magic
tech sky130A
magscale 1 2
timestamp 1623854003
<< checkpaint >>
rect -3932 -3932 21959 24103
<< locali >>
rect 3893 5763 3927 5865
rect 9321 5015 9355 5321
rect 6101 2295 6135 2465
rect 8953 2295 8987 2397
<< viali >>
rect 4537 17833 4571 17867
rect 6929 17765 6963 17799
rect 16405 17765 16439 17799
rect 1409 17697 1443 17731
rect 2329 17697 2363 17731
rect 3893 17697 3927 17731
rect 5549 17697 5583 17731
rect 7113 17697 7147 17731
rect 8953 17697 8987 17731
rect 10149 17697 10183 17731
rect 11989 17697 12023 17731
rect 14013 17697 14047 17731
rect 15393 17697 15427 17731
rect 16129 17697 16163 17731
rect 4169 17629 4203 17663
rect 10425 17629 10459 17663
rect 4537 17561 4571 17595
rect 16221 17561 16255 17595
rect 1593 17493 1627 17527
rect 2513 17493 2547 17527
rect 4077 17493 4111 17527
rect 5733 17493 5767 17527
rect 8769 17493 8803 17527
rect 12173 17493 12207 17527
rect 13829 17493 13863 17527
rect 15209 17493 15243 17527
rect 15945 17493 15979 17527
rect 4445 17289 4479 17323
rect 5089 17289 5123 17323
rect 6561 17289 6595 17323
rect 10977 17221 11011 17255
rect 11069 17221 11103 17255
rect 11713 17221 11747 17255
rect 12633 17221 12667 17255
rect 3801 17153 3835 17187
rect 3985 17153 4019 17187
rect 12173 17153 12207 17187
rect 12357 17153 12391 17187
rect 13185 17153 13219 17187
rect 1409 17085 1443 17119
rect 4537 17085 4571 17119
rect 5089 17085 5123 17119
rect 5641 17085 5675 17119
rect 5825 17085 5859 17119
rect 6653 17085 6687 17119
rect 6975 17085 7009 17119
rect 7078 17085 7112 17119
rect 7665 17085 7699 17119
rect 8401 17085 8435 17119
rect 9689 17085 9723 17119
rect 9965 17085 9999 17119
rect 10517 17085 10551 17119
rect 10609 17085 10643 17119
rect 11253 17085 11287 17119
rect 8585 17017 8619 17051
rect 9873 17017 9907 17051
rect 10057 17017 10091 17051
rect 12909 17017 12943 17051
rect 13093 17017 13127 17051
rect 1593 16949 1627 16983
rect 4077 16949 4111 16983
rect 10977 16949 11011 16983
rect 12081 16949 12115 16983
rect 4905 16745 4939 16779
rect 6009 16745 6043 16779
rect 10793 16745 10827 16779
rect 4629 16677 4663 16711
rect 7665 16677 7699 16711
rect 5089 16609 5123 16643
rect 5917 16609 5951 16643
rect 6193 16609 6227 16643
rect 6487 16609 6521 16643
rect 7205 16609 7239 16643
rect 7757 16609 7791 16643
rect 7941 16609 7975 16643
rect 8125 16609 8159 16643
rect 12449 16609 12483 16643
rect 13093 16609 13127 16643
rect 13369 16609 13403 16643
rect 13461 16609 13495 16643
rect 13921 16609 13955 16643
rect 14013 16541 14047 16575
rect 4721 16405 4755 16439
rect 10701 16405 10735 16439
rect 5641 16201 5675 16235
rect 8217 16201 8251 16235
rect 13829 16201 13863 16235
rect 4813 16133 4847 16167
rect 8677 16133 8711 16167
rect 8769 16133 8803 16167
rect 10517 16133 10551 16167
rect 2237 16065 2271 16099
rect 2421 16065 2455 16099
rect 4445 16065 4479 16099
rect 8309 16065 8343 16099
rect 2145 15997 2179 16031
rect 3801 15997 3835 16031
rect 4353 15997 4387 16031
rect 5825 15997 5859 16031
rect 7665 15997 7699 16031
rect 8217 15997 8251 16031
rect 8953 15997 8987 16031
rect 9505 15997 9539 16031
rect 10057 15997 10091 16031
rect 10149 15997 10183 16031
rect 13093 15997 13127 16031
rect 13645 15997 13679 16031
rect 4261 15929 4295 15963
rect 9965 15929 9999 15963
rect 13553 15929 13587 15963
rect 1777 15861 1811 15895
rect 4813 15861 4847 15895
rect 8677 15861 8711 15895
rect 10517 15861 10551 15895
rect 13737 15861 13771 15895
rect 2789 15657 2823 15691
rect 8677 15657 8711 15691
rect 14197 15657 14231 15691
rect 16313 15657 16347 15691
rect 2237 15589 2271 15623
rect 3249 15589 3283 15623
rect 11713 15589 11747 15623
rect 13277 15589 13311 15623
rect 1409 15521 1443 15555
rect 1777 15521 1811 15555
rect 2329 15521 2363 15555
rect 3065 15521 3099 15555
rect 3617 15521 3651 15555
rect 8585 15521 8619 15555
rect 13369 15521 13403 15555
rect 13829 15521 13863 15555
rect 14565 15521 14599 15555
rect 15761 15521 15795 15555
rect 16497 15521 16531 15555
rect 2421 15453 2455 15487
rect 13093 15453 13127 15487
rect 2789 15385 2823 15419
rect 3433 15385 3467 15419
rect 11897 15385 11931 15419
rect 13737 15385 13771 15419
rect 14197 15385 14231 15419
rect 14381 15385 14415 15419
rect 1593 15317 1627 15351
rect 15853 15317 15887 15351
rect 3985 15113 4019 15147
rect 7205 15113 7239 15147
rect 14105 15113 14139 15147
rect 15669 15113 15703 15147
rect 11713 15045 11747 15079
rect 16129 15045 16163 15079
rect 16221 15045 16255 15079
rect 4445 14977 4479 15011
rect 4629 14977 4663 15011
rect 6561 14977 6595 15011
rect 12173 14977 12207 15011
rect 12357 14977 12391 15011
rect 15761 14977 15795 15011
rect 1501 14909 1535 14943
rect 2237 14909 2271 14943
rect 2513 14909 2547 14943
rect 6745 14909 6779 14943
rect 15117 14909 15151 14943
rect 15669 14909 15703 14943
rect 16405 14909 16439 14943
rect 2421 14841 2455 14875
rect 4353 14841 4387 14875
rect 5457 14841 5491 14875
rect 5641 14841 5675 14875
rect 5825 14841 5859 14875
rect 5917 14841 5951 14875
rect 6101 14841 6135 14875
rect 6285 14841 6319 14875
rect 6837 14841 6871 14875
rect 11529 14841 11563 14875
rect 14013 14841 14047 14875
rect 2605 14773 2639 14807
rect 11437 14773 11471 14807
rect 12081 14773 12115 14807
rect 16129 14773 16163 14807
rect 4353 14569 4387 14603
rect 6377 14569 6411 14603
rect 8493 14569 8527 14603
rect 12265 14569 12299 14603
rect 7941 14501 7975 14535
rect 2605 14433 2639 14467
rect 4261 14433 4295 14467
rect 5733 14433 5767 14467
rect 5917 14433 5951 14467
rect 6193 14433 6227 14467
rect 6561 14433 6595 14467
rect 6745 14433 6779 14467
rect 6837 14433 6871 14467
rect 7481 14433 7515 14467
rect 8033 14433 8067 14467
rect 8585 14433 8619 14467
rect 9229 14433 9263 14467
rect 9781 14433 9815 14467
rect 10057 14433 10091 14467
rect 10425 14433 10459 14467
rect 10701 14433 10735 14467
rect 11253 14433 11287 14467
rect 11805 14433 11839 14467
rect 11897 14433 11931 14467
rect 12541 14433 12575 14467
rect 16497 14433 16531 14467
rect 1869 14365 1903 14399
rect 2513 14365 2547 14399
rect 4537 14365 4571 14399
rect 6653 14365 6687 14399
rect 8125 14365 8159 14399
rect 11437 14365 11471 14399
rect 6009 14297 6043 14331
rect 6101 14297 6135 14331
rect 8493 14297 8527 14331
rect 8677 14297 8711 14331
rect 12265 14297 12299 14331
rect 12357 14297 12391 14331
rect 3893 14229 3927 14263
rect 9229 14229 9263 14263
rect 10425 14229 10459 14263
rect 10609 14229 10643 14263
rect 16313 14229 16347 14263
rect 6193 14025 6227 14059
rect 13645 14025 13679 14059
rect 14105 14025 14139 14059
rect 16129 14025 16163 14059
rect 7849 13957 7883 13991
rect 8309 13957 8343 13991
rect 8401 13957 8435 13991
rect 15945 13957 15979 13991
rect 7941 13889 7975 13923
rect 15117 13889 15151 13923
rect 6101 13821 6135 13855
rect 7297 13821 7331 13855
rect 7849 13821 7883 13855
rect 8585 13821 8619 13855
rect 11805 13821 11839 13855
rect 11897 13821 11931 13855
rect 13093 13821 13127 13855
rect 13645 13821 13679 13855
rect 13737 13821 13771 13855
rect 14105 13821 14139 13855
rect 14933 13821 14967 13855
rect 15485 13821 15519 13855
rect 15577 13821 15611 13855
rect 16221 13821 16255 13855
rect 4721 13685 4755 13719
rect 4813 13685 4847 13719
rect 8309 13685 8343 13719
rect 12081 13685 12115 13719
rect 15945 13685 15979 13719
rect 2881 13481 2915 13515
rect 3249 13481 3283 13515
rect 4859 13481 4893 13515
rect 5825 13481 5859 13515
rect 8677 13481 8711 13515
rect 11805 13481 11839 13515
rect 12173 13481 12207 13515
rect 14105 13481 14139 13515
rect 2329 13413 2363 13447
rect 3985 13413 4019 13447
rect 10315 13413 10349 13447
rect 10793 13413 10827 13447
rect 12265 13413 12299 13447
rect 1869 13345 1903 13379
rect 2421 13345 2455 13379
rect 3157 13345 3191 13379
rect 3893 13345 3927 13379
rect 4445 13345 4479 13379
rect 5181 13345 5215 13379
rect 5733 13345 5767 13379
rect 8585 13345 8619 13379
rect 9781 13345 9815 13379
rect 10609 13345 10643 13379
rect 14013 13345 14047 13379
rect 2513 13277 2547 13311
rect 4537 13277 4571 13311
rect 6009 13277 6043 13311
rect 8769 13277 8803 13311
rect 9505 13277 9539 13311
rect 9689 13277 9723 13311
rect 10885 13277 10919 13311
rect 12403 13277 12437 13311
rect 2881 13209 2915 13243
rect 2973 13209 3007 13243
rect 4905 13209 4939 13243
rect 4997 13209 5031 13243
rect 5365 13209 5399 13243
rect 3341 13141 3375 13175
rect 8217 13141 8251 13175
rect 10149 13141 10183 13175
rect 6469 12937 6503 12971
rect 7113 12937 7147 12971
rect 7297 12937 7331 12971
rect 7573 12937 7607 12971
rect 11253 12937 11287 12971
rect 11713 12937 11747 12971
rect 14013 12937 14047 12971
rect 15393 12937 15427 12971
rect 4813 12869 4847 12903
rect 14473 12869 14507 12903
rect 14565 12869 14599 12903
rect 2329 12801 2363 12835
rect 4445 12801 4479 12835
rect 6653 12801 6687 12835
rect 6837 12801 6871 12835
rect 8125 12801 8159 12835
rect 9965 12801 9999 12835
rect 12357 12801 12391 12835
rect 15945 12801 15979 12835
rect 3249 12733 3283 12767
rect 3617 12733 3651 12767
rect 3801 12733 3835 12767
rect 4353 12733 4387 12767
rect 6745 12733 6779 12767
rect 6929 12733 6963 12767
rect 10793 12733 10827 12767
rect 10885 12733 10919 12767
rect 13461 12733 13495 12767
rect 14013 12733 14047 12767
rect 14105 12733 14139 12767
rect 14749 12733 14783 12767
rect 15853 12733 15887 12767
rect 2973 12665 3007 12699
rect 3433 12665 3467 12699
rect 3893 12665 3927 12699
rect 7265 12665 7299 12699
rect 7481 12665 7515 12699
rect 7941 12665 7975 12699
rect 11069 12665 11103 12699
rect 12173 12665 12207 12699
rect 4813 12597 4847 12631
rect 8033 12597 8067 12631
rect 12081 12597 12115 12631
rect 14473 12597 14507 12631
rect 15761 12597 15795 12631
rect 7113 12393 7147 12427
rect 9873 12393 9907 12427
rect 10609 12393 10643 12427
rect 11345 12393 11379 12427
rect 11989 12393 12023 12427
rect 15485 12393 15519 12427
rect 1869 12325 1903 12359
rect 11713 12325 11747 12359
rect 13001 12325 13035 12359
rect 1409 12257 1443 12291
rect 2053 12257 2087 12291
rect 6377 12257 6411 12291
rect 6837 12257 6871 12291
rect 7021 12257 7055 12291
rect 7573 12257 7607 12291
rect 7849 12257 7883 12291
rect 8033 12257 8067 12291
rect 10057 12257 10091 12291
rect 10333 12257 10367 12291
rect 10517 12257 10551 12291
rect 10793 12257 10827 12291
rect 11114 12257 11148 12291
rect 11253 12257 11287 12291
rect 11529 12257 11563 12291
rect 11805 12257 11839 12291
rect 11989 12257 12023 12291
rect 12449 12257 12483 12291
rect 12817 12257 12851 12291
rect 15761 12257 15795 12291
rect 15945 12257 15979 12291
rect 6101 12189 6135 12223
rect 8309 12189 8343 12223
rect 10885 12189 10919 12223
rect 15669 12189 15703 12223
rect 15853 12189 15887 12223
rect 1593 12121 1627 12155
rect 6561 12121 6595 12155
rect 10149 12121 10183 12155
rect 10241 12121 10275 12155
rect 10977 12121 11011 12155
rect 1777 12053 1811 12087
rect 6193 12053 6227 12087
rect 7757 12053 7791 12087
rect 7941 12053 7975 12087
rect 9689 11849 9723 11883
rect 10057 11849 10091 11883
rect 12633 11849 12667 11883
rect 13001 11849 13035 11883
rect 13737 11849 13771 11883
rect 15393 11849 15427 11883
rect 6653 11781 6687 11815
rect 7021 11781 7055 11815
rect 9229 11781 9263 11815
rect 13185 11781 13219 11815
rect 9137 11713 9171 11747
rect 9965 11713 9999 11747
rect 12173 11713 12207 11747
rect 14197 11713 14231 11747
rect 14381 11713 14415 11747
rect 15945 11713 15979 11747
rect 1593 11645 1627 11679
rect 2513 11645 2547 11679
rect 4997 11645 5031 11679
rect 6561 11645 6595 11679
rect 6745 11645 6779 11679
rect 6837 11645 6871 11679
rect 9045 11645 9079 11679
rect 9321 11645 9355 11679
rect 9505 11645 9539 11679
rect 10057 11645 10091 11679
rect 12081 11645 12115 11679
rect 12265 11645 12299 11679
rect 12357 11645 12391 11679
rect 12909 11645 12943 11679
rect 13093 11645 13127 11679
rect 13369 11645 13403 11679
rect 14841 11645 14875 11679
rect 15761 11645 15795 11679
rect 2237 11577 2271 11611
rect 14565 11577 14599 11611
rect 5089 11509 5123 11543
rect 8861 11509 8895 11543
rect 12541 11509 12575 11543
rect 14105 11509 14139 11543
rect 15853 11509 15887 11543
rect 5549 11305 5583 11339
rect 11253 11305 11287 11339
rect 16313 11305 16347 11339
rect 2973 11237 3007 11271
rect 4629 11237 4663 11271
rect 10333 11237 10367 11271
rect 14105 11237 14139 11271
rect 14473 11237 14507 11271
rect 15209 11237 15243 11271
rect 15393 11237 15427 11271
rect 1593 11169 1627 11203
rect 2329 11169 2363 11203
rect 4537 11169 4571 11203
rect 5089 11169 5123 11203
rect 5825 11169 5859 11203
rect 7757 11169 7791 11203
rect 7849 11169 7883 11203
rect 8493 11169 8527 11203
rect 8953 11169 8987 11203
rect 9965 11169 9999 11203
rect 10517 11169 10551 11203
rect 11161 11169 11195 11203
rect 11442 11169 11476 11203
rect 13185 11169 13219 11203
rect 14013 11169 14047 11203
rect 14381 11169 14415 11203
rect 14565 11169 14599 11203
rect 15485 11169 15519 11203
rect 16497 11169 16531 11203
rect 1961 11101 1995 11135
rect 2973 11101 3007 11135
rect 3065 11101 3099 11135
rect 5181 11101 5215 11135
rect 7941 11101 7975 11135
rect 10057 11101 10091 11135
rect 11529 11101 11563 11135
rect 2513 11033 2547 11067
rect 5549 11033 5583 11067
rect 5641 11033 5675 11067
rect 7389 11033 7423 11067
rect 8585 11033 8619 11067
rect 8769 11033 8803 11067
rect 10701 11033 10735 11067
rect 11805 11033 11839 11067
rect 14933 11033 14967 11067
rect 8217 10965 8251 10999
rect 8677 10965 8711 10999
rect 11621 10965 11655 10999
rect 13277 10965 13311 10999
rect 6469 10761 6503 10795
rect 6837 10761 6871 10795
rect 6929 10761 6963 10795
rect 7297 10761 7331 10795
rect 8125 10761 8159 10795
rect 8953 10761 8987 10795
rect 9413 10761 9447 10795
rect 10379 10761 10413 10795
rect 12817 10761 12851 10795
rect 3709 10693 3743 10727
rect 4353 10693 4387 10727
rect 6101 10693 6135 10727
rect 8493 10693 8527 10727
rect 9505 10693 9539 10727
rect 10241 10693 10275 10727
rect 11713 10693 11747 10727
rect 3157 10625 3191 10659
rect 4445 10625 4479 10659
rect 7941 10625 7975 10659
rect 8401 10625 8435 10659
rect 10149 10625 10183 10659
rect 12173 10625 12207 10659
rect 14473 10625 14507 10659
rect 1961 10557 1995 10591
rect 2789 10557 2823 10591
rect 3801 10557 3835 10591
rect 4353 10557 4387 10591
rect 4813 10557 4847 10591
rect 4905 10557 4939 10591
rect 5089 10557 5123 10591
rect 5917 10557 5951 10591
rect 6009 10557 6043 10591
rect 6193 10557 6227 10591
rect 6745 10557 6779 10591
rect 7021 10557 7055 10591
rect 7205 10557 7239 10591
rect 7665 10557 7699 10591
rect 8309 10557 8343 10591
rect 8585 10557 8619 10591
rect 8769 10557 8803 10591
rect 9229 10557 9263 10591
rect 9321 10557 9355 10591
rect 9689 10557 9723 10591
rect 10609 10557 10643 10591
rect 10793 10557 10827 10591
rect 11161 10557 11195 10591
rect 11437 10557 11471 10591
rect 11713 10557 11747 10591
rect 11897 10557 11931 10591
rect 12449 10557 12483 10591
rect 12633 10557 12667 10591
rect 12909 10557 12943 10591
rect 14197 10557 14231 10591
rect 14289 10557 14323 10591
rect 15669 10557 15703 10591
rect 2605 10489 2639 10523
rect 5733 10489 5767 10523
rect 9781 10489 9815 10523
rect 10517 10489 10551 10523
rect 3249 10421 3283 10455
rect 3341 10421 3375 10455
rect 4813 10421 4847 10455
rect 7757 10421 7791 10455
rect 11345 10421 11379 10455
rect 14473 10421 14507 10455
rect 15853 10421 15887 10455
rect 1593 10217 1627 10251
rect 12725 10149 12759 10183
rect 14933 10149 14967 10183
rect 1409 10081 1443 10115
rect 2145 10081 2179 10115
rect 3249 10081 3283 10115
rect 12449 10081 12483 10115
rect 13461 10081 13495 10115
rect 13737 10081 13771 10115
rect 13829 10081 13863 10115
rect 14381 10081 14415 10115
rect 2329 10013 2363 10047
rect 12725 10013 12759 10047
rect 14657 10013 14691 10047
rect 13553 9945 13587 9979
rect 14473 9945 14507 9979
rect 12541 9877 12575 9911
rect 14013 9877 14047 9911
rect 16405 9877 16439 9911
rect 12633 9673 12667 9707
rect 14473 9673 14507 9707
rect 4537 9605 4571 9639
rect 8217 9605 8251 9639
rect 10609 9605 10643 9639
rect 11253 9605 11287 9639
rect 13461 9605 13495 9639
rect 2513 9537 2547 9571
rect 5181 9537 5215 9571
rect 6469 9537 6503 9571
rect 11069 9537 11103 9571
rect 13369 9537 13403 9571
rect 2237 9469 2271 9503
rect 3525 9469 3559 9503
rect 3893 9469 3927 9503
rect 4537 9469 4571 9503
rect 5089 9469 5123 9503
rect 10057 9469 10091 9503
rect 10471 9469 10505 9503
rect 10885 9469 10919 9503
rect 11161 9469 11195 9503
rect 11345 9469 11379 9503
rect 11989 9469 12023 9503
rect 12173 9469 12207 9503
rect 12357 9469 12391 9503
rect 12817 9469 12851 9503
rect 13093 9469 13127 9503
rect 13277 9469 13311 9503
rect 13553 9469 13587 9503
rect 13829 9469 13863 9503
rect 13922 9469 13956 9503
rect 14105 9469 14139 9503
rect 14335 9469 14369 9503
rect 14565 9469 14599 9503
rect 15577 9469 15611 9503
rect 5365 9401 5399 9435
rect 6745 9401 6779 9435
rect 10241 9401 10275 9435
rect 10333 9401 10367 9435
rect 12265 9401 12299 9435
rect 13001 9401 13035 9435
rect 14197 9401 14231 9435
rect 14657 9401 14691 9435
rect 2053 9333 2087 9367
rect 3893 9333 3927 9367
rect 11529 9333 11563 9367
rect 12541 9333 12575 9367
rect 13737 9333 13771 9367
rect 15761 9333 15795 9367
rect 3617 9129 3651 9163
rect 4537 9129 4571 9163
rect 5825 9129 5859 9163
rect 6193 9129 6227 9163
rect 7021 9129 7055 9163
rect 9505 9129 9539 9163
rect 11621 9129 11655 9163
rect 16405 9129 16439 9163
rect 4353 9061 4387 9095
rect 5089 9061 5123 9095
rect 10701 9061 10735 9095
rect 11161 9061 11195 9095
rect 11529 9061 11563 9095
rect 12587 9061 12621 9095
rect 12725 9061 12759 9095
rect 12817 9061 12851 9095
rect 13093 9061 13127 9095
rect 14933 9061 14967 9095
rect 2053 8993 2087 9027
rect 3249 8993 3283 9027
rect 3893 8993 3927 9027
rect 4445 8993 4479 9027
rect 4721 8993 4755 9027
rect 5549 8993 5583 9027
rect 6837 8993 6871 9027
rect 9413 8993 9447 9027
rect 9919 8993 9953 9027
rect 10057 8993 10091 9027
rect 10149 8993 10183 9027
rect 10333 8993 10367 9027
rect 10609 8993 10643 9027
rect 10793 8993 10827 9027
rect 10911 8993 10945 9027
rect 11345 8993 11379 9027
rect 11621 8993 11655 9027
rect 11805 8993 11839 9027
rect 12909 8993 12943 9027
rect 13185 8993 13219 9027
rect 13369 8993 13403 9027
rect 2973 8925 3007 8959
rect 3157 8925 3191 8959
rect 4997 8925 5031 8959
rect 6285 8925 6319 8959
rect 6469 8925 6503 8959
rect 7113 8925 7147 8959
rect 7389 8925 7423 8959
rect 10425 8925 10459 8959
rect 11069 8925 11103 8959
rect 12449 8925 12483 8959
rect 13277 8925 13311 8959
rect 14657 8925 14691 8959
rect 8861 8857 8895 8891
rect 2421 8789 2455 8823
rect 9689 8789 9723 8823
rect 4905 8585 4939 8619
rect 6837 8585 6871 8619
rect 8493 8585 8527 8619
rect 9965 8585 9999 8619
rect 7389 8517 7423 8551
rect 7481 8449 7515 8483
rect 10425 8449 10459 8483
rect 10609 8449 10643 8483
rect 4813 8381 4847 8415
rect 6990 8381 7024 8415
rect 8677 8381 8711 8415
rect 13921 8381 13955 8415
rect 16497 8381 16531 8415
rect 7086 8313 7120 8347
rect 10333 8313 10367 8347
rect 14013 8245 14047 8279
rect 16313 8245 16347 8279
rect 1593 8041 1627 8075
rect 11621 8041 11655 8075
rect 14105 8041 14139 8075
rect 1409 7905 1443 7939
rect 2329 7905 2363 7939
rect 2973 7905 3007 7939
rect 3157 7905 3191 7939
rect 6653 7905 6687 7939
rect 9321 7905 9355 7939
rect 11805 7905 11839 7939
rect 11897 7905 11931 7939
rect 12173 7905 12207 7939
rect 13553 7905 13587 7939
rect 13829 7905 13863 7939
rect 13921 7905 13955 7939
rect 14381 7905 14415 7939
rect 14657 7905 14691 7939
rect 15669 7905 15703 7939
rect 2513 7701 2547 7735
rect 2789 7701 2823 7735
rect 6837 7701 6871 7735
rect 9137 7701 9171 7735
rect 12081 7701 12115 7735
rect 13645 7701 13679 7735
rect 14473 7701 14507 7735
rect 14749 7701 14783 7735
rect 15853 7701 15887 7735
rect 11897 7497 11931 7531
rect 12541 7497 12575 7531
rect 14473 7497 14507 7531
rect 16405 7497 16439 7531
rect 8217 7429 8251 7463
rect 14197 7429 14231 7463
rect 1685 7361 1719 7395
rect 3157 7361 3191 7395
rect 4537 7361 4571 7395
rect 5089 7361 5123 7395
rect 14289 7361 14323 7395
rect 14657 7361 14691 7395
rect 1409 7293 1443 7327
rect 3433 7293 3467 7327
rect 3617 7293 3651 7327
rect 3801 7293 3835 7327
rect 4077 7293 4111 7327
rect 4445 7293 4479 7327
rect 4905 7293 4939 7327
rect 5365 7293 5399 7327
rect 6469 7293 6503 7327
rect 10149 7293 10183 7327
rect 10793 7293 10827 7327
rect 10977 7293 11011 7327
rect 11253 7293 11287 7327
rect 11437 7293 11471 7327
rect 12081 7293 12115 7327
rect 12449 7293 12483 7327
rect 12541 7293 12575 7327
rect 12633 7293 12667 7327
rect 13553 7293 13587 7327
rect 13701 7293 13735 7327
rect 14018 7293 14052 7327
rect 14565 7293 14599 7327
rect 3525 7225 3559 7259
rect 4169 7225 4203 7259
rect 4261 7225 4295 7259
rect 4813 7225 4847 7259
rect 6745 7225 6779 7259
rect 9873 7225 9907 7259
rect 10333 7225 10367 7259
rect 12173 7225 12207 7259
rect 12265 7225 12299 7259
rect 13829 7225 13863 7259
rect 13921 7225 13955 7259
rect 14289 7225 14323 7259
rect 14933 7225 14967 7259
rect 3249 7157 3283 7191
rect 3893 7157 3927 7191
rect 4721 7157 4755 7191
rect 5181 7157 5215 7191
rect 8401 7157 8435 7191
rect 12909 7157 12943 7191
rect 3249 6953 3283 6987
rect 5733 6953 5767 6987
rect 6469 6885 6503 6919
rect 7941 6885 7975 6919
rect 8033 6885 8067 6919
rect 12633 6885 12667 6919
rect 6285 6817 6319 6851
rect 6561 6817 6595 6851
rect 7757 6817 7791 6851
rect 8149 6817 8183 6851
rect 10425 6817 10459 6851
rect 10517 6817 10551 6851
rect 11345 6817 11379 6851
rect 11713 6817 11747 6851
rect 12081 6817 12115 6851
rect 12357 6817 12391 6851
rect 12725 6817 12759 6851
rect 13737 6817 13771 6851
rect 13829 6817 13863 6851
rect 14105 6817 14139 6851
rect 1501 6749 1535 6783
rect 1777 6749 1811 6783
rect 3985 6749 4019 6783
rect 4261 6749 4295 6783
rect 11529 6749 11563 6783
rect 11989 6749 12023 6783
rect 12449 6749 12483 6783
rect 14013 6749 14047 6783
rect 6285 6681 6319 6715
rect 8309 6681 8343 6715
rect 11415 6681 11449 6715
rect 11805 6681 11839 6715
rect 11621 6613 11655 6647
rect 13553 6613 13587 6647
rect 2513 6409 2547 6443
rect 10701 6409 10735 6443
rect 12081 6409 12115 6443
rect 13369 6409 13403 6443
rect 15301 6409 15335 6443
rect 16313 6409 16347 6443
rect 11713 6341 11747 6375
rect 10241 6273 10275 6307
rect 11989 6273 12023 6307
rect 13829 6273 13863 6307
rect 2329 6205 2363 6239
rect 5181 6205 5215 6239
rect 6837 6205 6871 6239
rect 8217 6205 8251 6239
rect 8309 6205 8343 6239
rect 8585 6205 8619 6239
rect 8769 6205 8803 6239
rect 9965 6205 9999 6239
rect 10149 6205 10183 6239
rect 10333 6205 10367 6239
rect 10517 6205 10551 6239
rect 10793 6205 10827 6239
rect 10977 6205 11011 6239
rect 12081 6205 12115 6239
rect 13461 6205 13495 6239
rect 13553 6205 13587 6239
rect 15761 6205 15795 6239
rect 16497 6205 16531 6239
rect 8401 6137 8435 6171
rect 5273 6069 5307 6103
rect 6929 6069 6963 6103
rect 8033 6069 8067 6103
rect 8861 6069 8895 6103
rect 11069 6069 11103 6103
rect 15945 6069 15979 6103
rect 1593 5865 1627 5899
rect 3893 5865 3927 5899
rect 13737 5865 13771 5899
rect 14657 5865 14691 5899
rect 3433 5797 3467 5831
rect 10057 5797 10091 5831
rect 12265 5797 12299 5831
rect 16221 5797 16255 5831
rect 1409 5729 1443 5763
rect 3341 5729 3375 5763
rect 3525 5729 3559 5763
rect 3709 5729 3743 5763
rect 3893 5729 3927 5763
rect 3985 5729 4019 5763
rect 4169 5729 4203 5763
rect 7389 5729 7423 5763
rect 9321 5729 9355 5763
rect 9689 5729 9723 5763
rect 10149 5729 10183 5763
rect 14473 5729 14507 5763
rect 16497 5729 16531 5763
rect 7113 5661 7147 5695
rect 9413 5661 9447 5695
rect 9965 5661 9999 5695
rect 11989 5661 12023 5695
rect 3157 5525 3191 5559
rect 4169 5525 4203 5559
rect 5641 5525 5675 5559
rect 14749 5525 14783 5559
rect 6285 5321 6319 5355
rect 6469 5321 6503 5355
rect 9229 5321 9263 5355
rect 9321 5321 9355 5355
rect 13185 5321 13219 5355
rect 3893 5253 3927 5287
rect 4445 5253 4479 5287
rect 8125 5253 8159 5287
rect 1593 5185 1627 5219
rect 1869 5185 1903 5219
rect 3801 5185 3835 5219
rect 6929 5185 6963 5219
rect 7389 5185 7423 5219
rect 8309 5185 8343 5219
rect 8401 5185 8435 5219
rect 4320 5117 4354 5151
rect 4721 5117 4755 5151
rect 4997 5117 5031 5151
rect 6101 5117 6135 5151
rect 6653 5117 6687 5151
rect 6837 5117 6871 5151
rect 7021 5117 7055 5151
rect 7205 5117 7239 5151
rect 7297 5117 7331 5151
rect 7481 5117 7515 5151
rect 8861 5117 8895 5151
rect 9045 5117 9079 5151
rect 11253 5253 11287 5287
rect 9965 5185 9999 5219
rect 10425 5185 10459 5219
rect 9689 5117 9723 5151
rect 9873 5117 9907 5151
rect 10057 5117 10091 5151
rect 10241 5117 10275 5151
rect 10517 5117 10551 5151
rect 11529 5117 11563 5151
rect 11897 5117 11931 5151
rect 11989 5117 12023 5151
rect 12173 5117 12207 5151
rect 13001 5117 13035 5151
rect 9505 5049 9539 5083
rect 11253 5049 11287 5083
rect 11437 5049 11471 5083
rect 3341 4981 3375 5015
rect 4261 4981 4295 5015
rect 4537 4981 4571 5015
rect 4905 4981 4939 5015
rect 8769 4981 8803 5015
rect 9321 4981 9355 5015
rect 11805 4981 11839 5015
rect 12173 4981 12207 5015
rect 9689 4777 9723 4811
rect 16313 4777 16347 4811
rect 3985 4709 4019 4743
rect 9505 4709 9539 4743
rect 10057 4709 10091 4743
rect 11989 4709 12023 4743
rect 4077 4641 4111 4675
rect 4353 4641 4387 4675
rect 4445 4641 4479 4675
rect 5273 4641 5307 4675
rect 5452 4641 5486 4675
rect 5568 4641 5602 4675
rect 5687 4641 5721 4675
rect 6009 4641 6043 4675
rect 6193 4641 6227 4675
rect 9229 4641 9263 4675
rect 9413 4641 9447 4675
rect 9597 4641 9631 4675
rect 10149 4641 10183 4675
rect 10425 4641 10459 4675
rect 11069 4641 11103 4675
rect 11253 4641 11287 4675
rect 11805 4641 11839 4675
rect 12173 4641 12207 4675
rect 12569 4641 12603 4675
rect 12725 4641 12759 4675
rect 14013 4641 14047 4675
rect 15485 4641 15519 4675
rect 16497 4641 16531 4675
rect 6377 4573 6411 4607
rect 12357 4573 12391 4607
rect 12449 4573 12483 4607
rect 5917 4505 5951 4539
rect 4629 4437 4663 4471
rect 13829 4437 13863 4471
rect 15669 4437 15703 4471
rect 14828 4233 14862 4267
rect 5733 4165 5767 4199
rect 11345 4097 11379 4131
rect 12725 4097 12759 4131
rect 14565 4097 14599 4131
rect 5089 4029 5123 4063
rect 5181 4029 5215 4063
rect 5457 4029 5491 4063
rect 5641 4029 5675 4063
rect 6653 4029 6687 4063
rect 6745 4029 6779 4063
rect 7113 4029 7147 4063
rect 7389 4029 7423 4063
rect 11253 4029 11287 4063
rect 12081 4029 12115 4063
rect 12265 4029 12299 4063
rect 12449 4029 12483 4063
rect 6929 3961 6963 3995
rect 7024 3961 7058 3995
rect 7652 3961 7686 3995
rect 12357 3961 12391 3995
rect 13001 3961 13035 3995
rect 7297 3893 7331 3927
rect 9137 3893 9171 3927
rect 12633 3893 12667 3927
rect 14473 3893 14507 3927
rect 16313 3893 16347 3927
rect 1593 3689 1627 3723
rect 4445 3689 4479 3723
rect 4629 3689 4663 3723
rect 7205 3689 7239 3723
rect 8585 3689 8619 3723
rect 12081 3689 12115 3723
rect 1409 3553 1443 3587
rect 2329 3553 2363 3587
rect 3157 3553 3191 3587
rect 4570 3553 4604 3587
rect 5181 3553 5215 3587
rect 5365 3553 5399 3587
rect 6929 3553 6963 3587
rect 7113 3553 7147 3587
rect 7297 3553 7331 3587
rect 8401 3553 8435 3587
rect 10977 3553 11011 3587
rect 11345 3553 11379 3587
rect 11989 3553 12023 3587
rect 12541 3553 12575 3587
rect 12909 3553 12943 3587
rect 13001 3553 13035 3587
rect 15577 3553 15611 3587
rect 15761 3553 15795 3587
rect 16313 3553 16347 3587
rect 5089 3485 5123 3519
rect 5273 3485 5307 3519
rect 11805 3485 11839 3519
rect 16405 3485 16439 3519
rect 7481 3417 7515 3451
rect 11069 3417 11103 3451
rect 2513 3349 2547 3383
rect 3341 3349 3375 3383
rect 4997 3349 5031 3383
rect 15301 3349 15335 3383
rect 5365 3145 5399 3179
rect 6193 3145 6227 3179
rect 7573 3145 7607 3179
rect 10609 3145 10643 3179
rect 11345 3145 11379 3179
rect 13369 3145 13403 3179
rect 16497 3145 16531 3179
rect 5273 3077 5307 3111
rect 9965 3077 9999 3111
rect 13001 3077 13035 3111
rect 1409 3009 1443 3043
rect 3525 3009 3559 3043
rect 6837 3009 6871 3043
rect 7102 3009 7136 3043
rect 7297 3009 7331 3043
rect 11437 3009 11471 3043
rect 14749 3009 14783 3043
rect 15025 3009 15059 3043
rect 3433 2941 3467 2975
rect 5549 2941 5583 2975
rect 5641 2941 5675 2975
rect 5917 2941 5951 2975
rect 6285 2941 6319 2975
rect 7008 2941 7042 2975
rect 7205 2941 7239 2975
rect 7481 2941 7515 2975
rect 8401 2941 8435 2975
rect 8585 2941 8619 2975
rect 8677 2941 8711 2975
rect 8769 2941 8803 2975
rect 8953 2941 8987 2975
rect 9413 2941 9447 2975
rect 10057 2941 10091 2975
rect 10149 2941 10183 2975
rect 10425 2941 10459 2975
rect 10977 2941 11011 2975
rect 11069 2941 11103 2975
rect 11529 2941 11563 2975
rect 11713 2941 11747 2975
rect 11897 2941 11931 2975
rect 12081 2941 12115 2975
rect 12449 2941 12483 2975
rect 12817 2941 12851 2975
rect 13553 2941 13587 2975
rect 1685 2873 1719 2907
rect 3801 2873 3835 2907
rect 6009 2873 6043 2907
rect 9137 2873 9171 2907
rect 9229 2873 9263 2907
rect 11989 2873 12023 2907
rect 12633 2873 12667 2907
rect 12725 2873 12759 2907
rect 9597 2805 9631 2839
rect 10333 2805 10367 2839
rect 12265 2805 12299 2839
rect 1593 2601 1627 2635
rect 3893 2601 3927 2635
rect 5273 2601 5307 2635
rect 6377 2601 6411 2635
rect 7021 2601 7055 2635
rect 8309 2601 8343 2635
rect 11897 2601 11931 2635
rect 12081 2601 12115 2635
rect 12633 2601 12667 2635
rect 14565 2601 14599 2635
rect 15209 2601 15243 2635
rect 15761 2601 15795 2635
rect 16037 2601 16071 2635
rect 4169 2533 4203 2567
rect 4997 2533 5031 2567
rect 6745 2533 6779 2567
rect 7481 2533 7515 2567
rect 8769 2533 8803 2567
rect 9505 2533 9539 2567
rect 11253 2533 11287 2567
rect 1409 2465 1443 2499
rect 1869 2465 1903 2499
rect 3525 2465 3559 2499
rect 4077 2465 4111 2499
rect 4261 2465 4295 2499
rect 4445 2465 4479 2499
rect 4721 2465 4755 2499
rect 4813 2465 4847 2499
rect 5089 2465 5123 2499
rect 5733 2465 5767 2499
rect 6101 2465 6135 2499
rect 6193 2465 6227 2499
rect 7389 2465 7423 2499
rect 7757 2465 7791 2499
rect 8493 2465 8527 2499
rect 8677 2465 8711 2499
rect 11713 2465 11747 2499
rect 12022 2465 12056 2499
rect 12449 2465 12483 2499
rect 14381 2465 14415 2499
rect 14749 2465 14783 2499
rect 15393 2465 15427 2499
rect 15577 2465 15611 2499
rect 16221 2465 16255 2499
rect 16497 2465 16531 2499
rect 5825 2397 5859 2431
rect 4997 2329 5031 2363
rect 7297 2397 7331 2431
rect 7481 2397 7515 2431
rect 8953 2397 8987 2431
rect 9229 2397 9263 2431
rect 12541 2397 12575 2431
rect 14105 2397 14139 2431
rect 6929 2329 6963 2363
rect 16313 2329 16347 2363
rect 2053 2261 2087 2295
rect 3709 2261 3743 2295
rect 6101 2261 6135 2295
rect 7297 2261 7331 2295
rect 7665 2261 7699 2295
rect 8953 2261 8987 2295
rect 11529 2261 11563 2295
<< metal1 >>
rect 1104 17978 16836 18000
rect 1104 17926 6226 17978
rect 6278 17926 6290 17978
rect 6342 17926 6354 17978
rect 6406 17926 6418 17978
rect 6470 17926 11470 17978
rect 11522 17926 11534 17978
rect 11586 17926 11598 17978
rect 11650 17926 11662 17978
rect 11714 17926 16836 17978
rect 1104 17904 16836 17926
rect 4525 17867 4583 17873
rect 4525 17833 4537 17867
rect 4571 17864 4583 17867
rect 5074 17864 5080 17876
rect 4571 17836 5080 17864
rect 4571 17833 4583 17836
rect 4525 17827 4583 17833
rect 5074 17824 5080 17836
rect 5132 17824 5138 17876
rect 6914 17796 6920 17808
rect 6875 17768 6920 17796
rect 6914 17756 6920 17768
rect 6972 17756 6978 17808
rect 16393 17799 16451 17805
rect 16393 17765 16405 17799
rect 16439 17796 16451 17799
rect 17034 17796 17040 17808
rect 16439 17768 17040 17796
rect 16439 17765 16451 17768
rect 16393 17759 16451 17765
rect 17034 17756 17040 17768
rect 17092 17756 17098 17808
rect 474 17688 480 17740
rect 532 17728 538 17740
rect 1397 17731 1455 17737
rect 1397 17728 1409 17731
rect 532 17700 1409 17728
rect 532 17688 538 17700
rect 1397 17697 1409 17700
rect 1443 17697 1455 17731
rect 2314 17728 2320 17740
rect 2275 17700 2320 17728
rect 1397 17691 1455 17697
rect 2314 17688 2320 17700
rect 2372 17688 2378 17740
rect 3694 17688 3700 17740
rect 3752 17728 3758 17740
rect 3881 17731 3939 17737
rect 3881 17728 3893 17731
rect 3752 17700 3893 17728
rect 3752 17688 3758 17700
rect 3881 17697 3893 17700
rect 3927 17697 3939 17731
rect 5534 17728 5540 17740
rect 5495 17700 5540 17728
rect 3881 17691 3939 17697
rect 5534 17688 5540 17700
rect 5592 17688 5598 17740
rect 6546 17688 6552 17740
rect 6604 17728 6610 17740
rect 7101 17731 7159 17737
rect 7101 17728 7113 17731
rect 6604 17700 7113 17728
rect 6604 17688 6610 17700
rect 7101 17697 7113 17700
rect 7147 17697 7159 17731
rect 7101 17691 7159 17697
rect 8754 17688 8760 17740
rect 8812 17728 8818 17740
rect 8941 17731 8999 17737
rect 8941 17728 8953 17731
rect 8812 17700 8953 17728
rect 8812 17688 8818 17700
rect 8941 17697 8953 17700
rect 8987 17697 8999 17731
rect 10134 17728 10140 17740
rect 10095 17700 10140 17728
rect 8941 17691 8999 17697
rect 10134 17688 10140 17700
rect 10192 17688 10198 17740
rect 11974 17728 11980 17740
rect 11935 17700 11980 17728
rect 11974 17688 11980 17700
rect 12032 17688 12038 17740
rect 13814 17688 13820 17740
rect 13872 17728 13878 17740
rect 14001 17731 14059 17737
rect 14001 17728 14013 17731
rect 13872 17700 14013 17728
rect 13872 17688 13878 17700
rect 14001 17697 14013 17700
rect 14047 17697 14059 17731
rect 14001 17691 14059 17697
rect 15194 17688 15200 17740
rect 15252 17728 15258 17740
rect 15381 17731 15439 17737
rect 15381 17728 15393 17731
rect 15252 17700 15393 17728
rect 15252 17688 15258 17700
rect 15381 17697 15393 17700
rect 15427 17697 15439 17731
rect 16114 17728 16120 17740
rect 16075 17700 16120 17728
rect 15381 17691 15439 17697
rect 16114 17688 16120 17700
rect 16172 17688 16178 17740
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17660 4215 17663
rect 4430 17660 4436 17672
rect 4203 17632 4436 17660
rect 4203 17629 4215 17632
rect 4157 17623 4215 17629
rect 4430 17620 4436 17632
rect 4488 17620 4494 17672
rect 10413 17663 10471 17669
rect 10413 17629 10425 17663
rect 10459 17660 10471 17663
rect 12434 17660 12440 17672
rect 10459 17632 12440 17660
rect 10459 17629 10471 17632
rect 10413 17623 10471 17629
rect 12434 17620 12440 17632
rect 12492 17620 12498 17672
rect 4246 17552 4252 17604
rect 4304 17592 4310 17604
rect 4525 17595 4583 17601
rect 4304 17564 4476 17592
rect 4304 17552 4310 17564
rect 1578 17524 1584 17536
rect 1539 17496 1584 17524
rect 1578 17484 1584 17496
rect 1636 17484 1642 17536
rect 2501 17527 2559 17533
rect 2501 17493 2513 17527
rect 2547 17524 2559 17527
rect 3970 17524 3976 17536
rect 2547 17496 3976 17524
rect 2547 17493 2559 17496
rect 2501 17487 2559 17493
rect 3970 17484 3976 17496
rect 4028 17484 4034 17536
rect 4065 17527 4123 17533
rect 4065 17493 4077 17527
rect 4111 17524 4123 17527
rect 4338 17524 4344 17536
rect 4111 17496 4344 17524
rect 4111 17493 4123 17496
rect 4065 17487 4123 17493
rect 4338 17484 4344 17496
rect 4396 17484 4402 17536
rect 4448 17524 4476 17564
rect 4525 17561 4537 17595
rect 4571 17592 4583 17595
rect 4890 17592 4896 17604
rect 4571 17564 4896 17592
rect 4571 17561 4583 17564
rect 4525 17555 4583 17561
rect 4890 17552 4896 17564
rect 4948 17552 4954 17604
rect 16209 17595 16267 17601
rect 16209 17592 16221 17595
rect 5092 17564 16221 17592
rect 5092 17524 5120 17564
rect 16209 17561 16221 17564
rect 16255 17561 16267 17595
rect 16209 17555 16267 17561
rect 5718 17524 5724 17536
rect 4448 17496 5120 17524
rect 5679 17496 5724 17524
rect 5718 17484 5724 17496
rect 5776 17484 5782 17536
rect 8662 17484 8668 17536
rect 8720 17524 8726 17536
rect 8757 17527 8815 17533
rect 8757 17524 8769 17527
rect 8720 17496 8769 17524
rect 8720 17484 8726 17496
rect 8757 17493 8769 17496
rect 8803 17493 8815 17527
rect 12158 17524 12164 17536
rect 12119 17496 12164 17524
rect 8757 17487 8815 17493
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 13817 17527 13875 17533
rect 13817 17493 13829 17527
rect 13863 17524 13875 17527
rect 15010 17524 15016 17536
rect 13863 17496 15016 17524
rect 13863 17493 13875 17496
rect 13817 17487 13875 17493
rect 15010 17484 15016 17496
rect 15068 17484 15074 17536
rect 15194 17524 15200 17536
rect 15155 17496 15200 17524
rect 15194 17484 15200 17496
rect 15252 17484 15258 17536
rect 15930 17524 15936 17536
rect 15891 17496 15936 17524
rect 15930 17484 15936 17496
rect 15988 17484 15994 17536
rect 1104 17434 16836 17456
rect 1104 17382 3604 17434
rect 3656 17382 3668 17434
rect 3720 17382 3732 17434
rect 3784 17382 3796 17434
rect 3848 17382 8848 17434
rect 8900 17382 8912 17434
rect 8964 17382 8976 17434
rect 9028 17382 9040 17434
rect 9092 17382 14092 17434
rect 14144 17382 14156 17434
rect 14208 17382 14220 17434
rect 14272 17382 14284 17434
rect 14336 17382 16836 17434
rect 1104 17360 16836 17382
rect 4430 17320 4436 17332
rect 4391 17292 4436 17320
rect 4430 17280 4436 17292
rect 4488 17280 4494 17332
rect 5074 17320 5080 17332
rect 5035 17292 5080 17320
rect 5074 17280 5080 17292
rect 5132 17280 5138 17332
rect 6546 17320 6552 17332
rect 6507 17292 6552 17320
rect 6546 17280 6552 17292
rect 6604 17280 6610 17332
rect 15194 17320 15200 17332
rect 12176 17292 15200 17320
rect 2682 17212 2688 17264
rect 2740 17252 2746 17264
rect 4246 17252 4252 17264
rect 2740 17224 4252 17252
rect 2740 17212 2746 17224
rect 4246 17212 4252 17224
rect 4304 17212 4310 17264
rect 3789 17187 3847 17193
rect 3789 17153 3801 17187
rect 3835 17153 3847 17187
rect 3970 17184 3976 17196
rect 3931 17156 3976 17184
rect 3789 17147 3847 17153
rect 1394 17116 1400 17128
rect 1355 17088 1400 17116
rect 1394 17076 1400 17088
rect 1452 17076 1458 17128
rect 3804 17116 3832 17147
rect 3970 17144 3976 17156
rect 4028 17144 4034 17196
rect 4062 17116 4068 17128
rect 3804 17088 4068 17116
rect 4062 17076 4068 17088
rect 4120 17076 4126 17128
rect 4448 17116 4476 17280
rect 10965 17255 11023 17261
rect 10965 17221 10977 17255
rect 11011 17252 11023 17255
rect 11057 17255 11115 17261
rect 11057 17252 11069 17255
rect 11011 17224 11069 17252
rect 11011 17221 11023 17224
rect 10965 17215 11023 17221
rect 11057 17221 11069 17224
rect 11103 17221 11115 17255
rect 11057 17215 11115 17221
rect 11701 17255 11759 17261
rect 11701 17221 11713 17255
rect 11747 17221 11759 17255
rect 11701 17215 11759 17221
rect 10778 17184 10784 17196
rect 5828 17156 10784 17184
rect 4525 17119 4583 17125
rect 4525 17116 4537 17119
rect 4448 17088 4537 17116
rect 4525 17085 4537 17088
rect 4571 17085 4583 17119
rect 4525 17079 4583 17085
rect 5077 17119 5135 17125
rect 5077 17085 5089 17119
rect 5123 17116 5135 17119
rect 5166 17116 5172 17128
rect 5123 17088 5172 17116
rect 5123 17085 5135 17088
rect 5077 17079 5135 17085
rect 5166 17076 5172 17088
rect 5224 17116 5230 17128
rect 5828 17125 5856 17156
rect 10778 17144 10784 17156
rect 10836 17144 10842 17196
rect 11716 17184 11744 17215
rect 12176 17193 12204 17292
rect 15194 17280 15200 17292
rect 15252 17280 15258 17332
rect 12618 17252 12624 17264
rect 12579 17224 12624 17252
rect 12618 17212 12624 17224
rect 12676 17212 12682 17264
rect 10888 17156 11744 17184
rect 12161 17187 12219 17193
rect 5629 17119 5687 17125
rect 5629 17116 5641 17119
rect 5224 17088 5641 17116
rect 5224 17076 5230 17088
rect 5629 17085 5641 17088
rect 5675 17085 5687 17119
rect 5629 17079 5687 17085
rect 5813 17119 5871 17125
rect 5813 17085 5825 17119
rect 5859 17085 5871 17119
rect 5813 17079 5871 17085
rect 6641 17119 6699 17125
rect 6641 17085 6653 17119
rect 6687 17116 6699 17119
rect 6963 17119 7021 17125
rect 6963 17116 6975 17119
rect 6687 17088 6975 17116
rect 6687 17085 6699 17088
rect 6641 17079 6699 17085
rect 6963 17085 6975 17088
rect 7009 17085 7021 17119
rect 6963 17079 7021 17085
rect 7066 17119 7124 17125
rect 7066 17085 7078 17119
rect 7112 17116 7124 17119
rect 7112 17085 7144 17116
rect 7066 17079 7144 17085
rect 5994 17048 6000 17060
rect 1596 17020 6000 17048
rect 1596 16989 1624 17020
rect 5994 17008 6000 17020
rect 6052 17008 6058 17060
rect 7116 17048 7144 17079
rect 7190 17076 7196 17128
rect 7248 17116 7254 17128
rect 7653 17119 7711 17125
rect 7653 17116 7665 17119
rect 7248 17088 7665 17116
rect 7248 17076 7254 17088
rect 7653 17085 7665 17088
rect 7699 17085 7711 17119
rect 8386 17116 8392 17128
rect 8299 17088 8392 17116
rect 7653 17079 7711 17085
rect 8386 17076 8392 17088
rect 8444 17116 8450 17128
rect 9677 17119 9735 17125
rect 9677 17116 9689 17119
rect 8444 17088 9689 17116
rect 8444 17076 8450 17088
rect 9677 17085 9689 17088
rect 9723 17085 9735 17119
rect 9677 17079 9735 17085
rect 9953 17119 10011 17125
rect 9953 17085 9965 17119
rect 9999 17085 10011 17119
rect 9953 17079 10011 17085
rect 10505 17119 10563 17125
rect 10505 17085 10517 17119
rect 10551 17116 10563 17119
rect 10597 17119 10655 17125
rect 10597 17116 10609 17119
rect 10551 17088 10609 17116
rect 10551 17085 10563 17088
rect 10505 17079 10563 17085
rect 10597 17085 10609 17088
rect 10643 17116 10655 17119
rect 10888 17116 10916 17156
rect 12161 17153 12173 17187
rect 12207 17153 12219 17187
rect 12161 17147 12219 17153
rect 12345 17187 12403 17193
rect 12345 17153 12357 17187
rect 12391 17184 12403 17187
rect 12434 17184 12440 17196
rect 12391 17156 12440 17184
rect 12391 17153 12403 17156
rect 12345 17147 12403 17153
rect 12434 17144 12440 17156
rect 12492 17184 12498 17196
rect 13170 17184 13176 17196
rect 12492 17156 13176 17184
rect 12492 17144 12498 17156
rect 13170 17144 13176 17156
rect 13228 17144 13234 17196
rect 10643 17088 10916 17116
rect 10643 17085 10655 17088
rect 10597 17079 10655 17085
rect 8404 17048 8432 17076
rect 8570 17048 8576 17060
rect 7116 17020 8432 17048
rect 8531 17020 8576 17048
rect 8570 17008 8576 17020
rect 8628 17008 8634 17060
rect 9858 17048 9864 17060
rect 9771 17020 9864 17048
rect 9858 17008 9864 17020
rect 9916 17048 9922 17060
rect 9968 17048 9996 17079
rect 10962 17076 10968 17128
rect 11020 17116 11026 17128
rect 11241 17119 11299 17125
rect 11241 17116 11253 17119
rect 11020 17088 11253 17116
rect 11020 17076 11026 17088
rect 11241 17085 11253 17088
rect 11287 17085 11299 17119
rect 15930 17116 15936 17128
rect 11241 17079 11299 17085
rect 13096 17088 15936 17116
rect 9916 17020 9996 17048
rect 9916 17008 9922 17020
rect 1581 16983 1639 16989
rect 1581 16949 1593 16983
rect 1627 16949 1639 16983
rect 1581 16943 1639 16949
rect 4065 16983 4123 16989
rect 4065 16949 4077 16983
rect 4111 16980 4123 16983
rect 5626 16980 5632 16992
rect 4111 16952 5632 16980
rect 4111 16949 4123 16952
rect 4065 16943 4123 16949
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 9968 16980 9996 17020
rect 10045 17051 10103 17057
rect 10045 17017 10057 17051
rect 10091 17048 10103 17051
rect 10778 17048 10784 17060
rect 10091 17020 10784 17048
rect 10091 17017 10103 17020
rect 10045 17011 10103 17017
rect 10778 17008 10784 17020
rect 10836 17048 10842 17060
rect 10836 17020 11008 17048
rect 10836 17008 10842 17020
rect 10870 16980 10876 16992
rect 9968 16952 10876 16980
rect 10870 16940 10876 16952
rect 10928 16940 10934 16992
rect 10980 16989 11008 17020
rect 11054 17008 11060 17060
rect 11112 17048 11118 17060
rect 12526 17048 12532 17060
rect 11112 17020 12532 17048
rect 11112 17008 11118 17020
rect 12526 17008 12532 17020
rect 12584 17008 12590 17060
rect 12894 17048 12900 17060
rect 12855 17020 12900 17048
rect 12894 17008 12900 17020
rect 12952 17008 12958 17060
rect 13096 17057 13124 17088
rect 15930 17076 15936 17088
rect 15988 17076 15994 17128
rect 13081 17051 13139 17057
rect 13081 17017 13093 17051
rect 13127 17017 13139 17051
rect 13081 17011 13139 17017
rect 10965 16983 11023 16989
rect 10965 16949 10977 16983
rect 11011 16949 11023 16983
rect 12066 16980 12072 16992
rect 12027 16952 12072 16980
rect 10965 16943 11023 16949
rect 12066 16940 12072 16952
rect 12124 16940 12130 16992
rect 1104 16890 16836 16912
rect 1104 16838 6226 16890
rect 6278 16838 6290 16890
rect 6342 16838 6354 16890
rect 6406 16838 6418 16890
rect 6470 16838 11470 16890
rect 11522 16838 11534 16890
rect 11586 16838 11598 16890
rect 11650 16838 11662 16890
rect 11714 16838 16836 16890
rect 1104 16816 16836 16838
rect 4890 16776 4896 16788
rect 4851 16748 4896 16776
rect 4890 16736 4896 16748
rect 4948 16736 4954 16788
rect 5074 16736 5080 16788
rect 5132 16736 5138 16788
rect 5994 16776 6000 16788
rect 5955 16748 6000 16776
rect 5994 16736 6000 16748
rect 6052 16736 6058 16788
rect 10778 16776 10784 16788
rect 10739 16748 10784 16776
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 4617 16711 4675 16717
rect 4617 16677 4629 16711
rect 4663 16708 4675 16711
rect 5092 16708 5120 16736
rect 4663 16680 5120 16708
rect 7653 16711 7711 16717
rect 4663 16677 4675 16680
rect 4617 16671 4675 16677
rect 7653 16677 7665 16711
rect 7699 16708 7711 16711
rect 8386 16708 8392 16720
rect 7699 16680 8392 16708
rect 7699 16677 7711 16680
rect 7653 16671 7711 16677
rect 8386 16668 8392 16680
rect 8444 16668 8450 16720
rect 12618 16708 12624 16720
rect 12452 16680 12624 16708
rect 5074 16640 5080 16652
rect 5035 16612 5080 16640
rect 5074 16600 5080 16612
rect 5132 16600 5138 16652
rect 5902 16640 5908 16652
rect 5863 16612 5908 16640
rect 5902 16600 5908 16612
rect 5960 16600 5966 16652
rect 6086 16600 6092 16652
rect 6144 16640 6150 16652
rect 6181 16643 6239 16649
rect 6181 16640 6193 16643
rect 6144 16612 6193 16640
rect 6144 16600 6150 16612
rect 6181 16609 6193 16612
rect 6227 16609 6239 16643
rect 6181 16603 6239 16609
rect 6475 16643 6533 16649
rect 6475 16609 6487 16643
rect 6521 16640 6533 16643
rect 7190 16640 7196 16652
rect 6521 16612 7196 16640
rect 6521 16609 6533 16612
rect 6475 16603 6533 16609
rect 7190 16600 7196 16612
rect 7248 16600 7254 16652
rect 7745 16643 7803 16649
rect 7745 16609 7757 16643
rect 7791 16640 7803 16643
rect 7929 16643 7987 16649
rect 7929 16640 7941 16643
rect 7791 16612 7941 16640
rect 7791 16609 7803 16612
rect 7745 16603 7803 16609
rect 7929 16609 7941 16612
rect 7975 16609 7987 16643
rect 8110 16640 8116 16652
rect 8071 16612 8116 16640
rect 7929 16603 7987 16609
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 12452 16649 12480 16680
rect 12618 16668 12624 16680
rect 12676 16708 12682 16720
rect 12676 16680 13492 16708
rect 12676 16668 12682 16680
rect 12437 16643 12495 16649
rect 12437 16609 12449 16643
rect 12483 16609 12495 16643
rect 12437 16603 12495 16609
rect 12526 16600 12532 16652
rect 12584 16640 12590 16652
rect 13081 16643 13139 16649
rect 13081 16640 13093 16643
rect 12584 16612 13093 16640
rect 12584 16600 12590 16612
rect 13081 16609 13093 16612
rect 13127 16609 13139 16643
rect 13354 16640 13360 16652
rect 13315 16612 13360 16640
rect 13081 16603 13139 16609
rect 13096 16572 13124 16603
rect 13354 16600 13360 16612
rect 13412 16600 13418 16652
rect 13464 16649 13492 16680
rect 13449 16643 13507 16649
rect 13449 16609 13461 16643
rect 13495 16609 13507 16643
rect 13909 16643 13967 16649
rect 13909 16640 13921 16643
rect 13449 16603 13507 16609
rect 13556 16612 13921 16640
rect 13556 16572 13584 16612
rect 13909 16609 13921 16612
rect 13955 16609 13967 16643
rect 13909 16603 13967 16609
rect 13096 16544 13584 16572
rect 13814 16532 13820 16584
rect 13872 16572 13878 16584
rect 14001 16575 14059 16581
rect 14001 16572 14013 16575
rect 13872 16544 14013 16572
rect 13872 16532 13878 16544
rect 14001 16541 14013 16544
rect 14047 16541 14059 16575
rect 14001 16535 14059 16541
rect 4706 16436 4712 16448
rect 4667 16408 4712 16436
rect 4706 16396 4712 16408
rect 4764 16396 4770 16448
rect 10686 16436 10692 16448
rect 10647 16408 10692 16436
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 1104 16346 16836 16368
rect 1104 16294 3604 16346
rect 3656 16294 3668 16346
rect 3720 16294 3732 16346
rect 3784 16294 3796 16346
rect 3848 16294 8848 16346
rect 8900 16294 8912 16346
rect 8964 16294 8976 16346
rect 9028 16294 9040 16346
rect 9092 16294 14092 16346
rect 14144 16294 14156 16346
rect 14208 16294 14220 16346
rect 14272 16294 14284 16346
rect 14336 16294 16836 16346
rect 1104 16272 16836 16294
rect 4062 16232 4068 16244
rect 2746 16204 4068 16232
rect 1578 16056 1584 16108
rect 1636 16096 1642 16108
rect 2225 16099 2283 16105
rect 2225 16096 2237 16099
rect 1636 16068 2237 16096
rect 1636 16056 1642 16068
rect 2225 16065 2237 16068
rect 2271 16065 2283 16099
rect 2225 16059 2283 16065
rect 2409 16099 2467 16105
rect 2409 16065 2421 16099
rect 2455 16096 2467 16099
rect 2746 16096 2774 16204
rect 4062 16192 4068 16204
rect 4120 16192 4126 16244
rect 5626 16232 5632 16244
rect 5587 16204 5632 16232
rect 5626 16192 5632 16204
rect 5684 16192 5690 16244
rect 8110 16192 8116 16244
rect 8168 16232 8174 16244
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 8168 16204 8217 16232
rect 8168 16192 8174 16204
rect 8205 16201 8217 16204
rect 8251 16201 8263 16235
rect 13814 16232 13820 16244
rect 8205 16195 8263 16201
rect 8312 16204 12434 16232
rect 13775 16204 13820 16232
rect 2455 16068 2774 16096
rect 3712 16136 4660 16164
rect 2455 16065 2467 16068
rect 2409 16059 2467 16065
rect 2133 16031 2191 16037
rect 2133 15997 2145 16031
rect 2179 16028 2191 16031
rect 3712 16028 3740 16136
rect 4433 16099 4491 16105
rect 4433 16096 4445 16099
rect 3988 16068 4445 16096
rect 3988 16040 4016 16068
rect 4433 16065 4445 16068
rect 4479 16065 4491 16099
rect 4632 16096 4660 16136
rect 4706 16124 4712 16176
rect 4764 16164 4770 16176
rect 4801 16167 4859 16173
rect 4801 16164 4813 16167
rect 4764 16136 4813 16164
rect 4764 16124 4770 16136
rect 4801 16133 4813 16136
rect 4847 16133 4859 16167
rect 4801 16127 4859 16133
rect 6822 16096 6828 16108
rect 4632 16068 6828 16096
rect 4433 16059 4491 16065
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 8312 16105 8340 16204
rect 8665 16167 8723 16173
rect 8665 16133 8677 16167
rect 8711 16164 8723 16167
rect 8757 16167 8815 16173
rect 8757 16164 8769 16167
rect 8711 16136 8769 16164
rect 8711 16133 8723 16136
rect 8665 16127 8723 16133
rect 8757 16133 8769 16136
rect 8803 16133 8815 16167
rect 8757 16127 8815 16133
rect 9490 16124 9496 16176
rect 9548 16164 9554 16176
rect 10505 16167 10563 16173
rect 9548 16136 10180 16164
rect 9548 16124 9554 16136
rect 8297 16099 8355 16105
rect 8297 16096 8309 16099
rect 7668 16068 8309 16096
rect 2179 16000 3740 16028
rect 3789 16031 3847 16037
rect 2179 15997 2191 16000
rect 2133 15991 2191 15997
rect 3789 15997 3801 16031
rect 3835 16028 3847 16031
rect 3970 16028 3976 16040
rect 3835 16000 3976 16028
rect 3835 15997 3847 16000
rect 3789 15991 3847 15997
rect 3970 15988 3976 16000
rect 4028 15988 4034 16040
rect 4341 16031 4399 16037
rect 4341 15997 4353 16031
rect 4387 16028 4399 16031
rect 5074 16028 5080 16040
rect 4387 16000 5080 16028
rect 4387 15997 4399 16000
rect 4341 15991 4399 15997
rect 5074 15988 5080 16000
rect 5132 15988 5138 16040
rect 5626 15988 5632 16040
rect 5684 16028 5690 16040
rect 7668 16037 7696 16068
rect 8297 16065 8309 16068
rect 8343 16065 8355 16099
rect 8297 16059 8355 16065
rect 5813 16031 5871 16037
rect 5813 16028 5825 16031
rect 5684 16000 5825 16028
rect 5684 15988 5690 16000
rect 5813 15997 5825 16000
rect 5859 15997 5871 16031
rect 5813 15991 5871 15997
rect 7653 16031 7711 16037
rect 7653 15997 7665 16031
rect 7699 15997 7711 16031
rect 7653 15991 7711 15997
rect 8205 16031 8263 16037
rect 8205 15997 8217 16031
rect 8251 16028 8263 16031
rect 8570 16028 8576 16040
rect 8251 16000 8576 16028
rect 8251 15997 8263 16000
rect 8205 15991 8263 15997
rect 8570 15988 8576 16000
rect 8628 16028 8634 16040
rect 8941 16031 8999 16037
rect 8941 16028 8953 16031
rect 8628 16000 8953 16028
rect 8628 15988 8634 16000
rect 8941 15997 8953 16000
rect 8987 15997 8999 16031
rect 9490 16028 9496 16040
rect 9451 16000 9496 16028
rect 8941 15991 8999 15997
rect 9490 15988 9496 16000
rect 9548 15988 9554 16040
rect 9858 15988 9864 16040
rect 9916 16028 9922 16040
rect 10152 16037 10180 16136
rect 10505 16133 10517 16167
rect 10551 16164 10563 16167
rect 10686 16164 10692 16176
rect 10551 16136 10692 16164
rect 10551 16133 10563 16136
rect 10505 16127 10563 16133
rect 10686 16124 10692 16136
rect 10744 16124 10750 16176
rect 12406 16164 12434 16204
rect 13814 16192 13820 16204
rect 13872 16192 13878 16244
rect 14918 16164 14924 16176
rect 12406 16136 14924 16164
rect 14918 16124 14924 16136
rect 14976 16124 14982 16176
rect 13354 16056 13360 16108
rect 13412 16096 13418 16108
rect 13412 16068 13676 16096
rect 13412 16056 13418 16068
rect 10045 16031 10103 16037
rect 10045 16028 10057 16031
rect 9916 16000 10057 16028
rect 9916 15988 9922 16000
rect 10045 15997 10057 16000
rect 10091 15997 10103 16031
rect 10045 15991 10103 15997
rect 10137 16031 10195 16037
rect 10137 15997 10149 16031
rect 10183 15997 10195 16031
rect 10137 15991 10195 15997
rect 13081 16031 13139 16037
rect 13081 15997 13093 16031
rect 13127 16028 13139 16031
rect 13446 16028 13452 16040
rect 13127 16000 13452 16028
rect 13127 15997 13139 16000
rect 13081 15991 13139 15997
rect 13446 15988 13452 16000
rect 13504 15988 13510 16040
rect 13648 16037 13676 16068
rect 13633 16031 13691 16037
rect 13633 15997 13645 16031
rect 13679 16028 13691 16031
rect 13906 16028 13912 16040
rect 13679 16000 13912 16028
rect 13679 15997 13691 16000
rect 13633 15991 13691 15997
rect 13906 15988 13912 16000
rect 13964 15988 13970 16040
rect 4249 15963 4307 15969
rect 4249 15929 4261 15963
rect 4295 15929 4307 15963
rect 4249 15923 4307 15929
rect 9953 15963 10011 15969
rect 9953 15929 9965 15963
rect 9999 15929 10011 15963
rect 9953 15923 10011 15929
rect 13541 15963 13599 15969
rect 13541 15929 13553 15963
rect 13587 15929 13599 15963
rect 13541 15923 13599 15929
rect 1762 15892 1768 15904
rect 1723 15864 1768 15892
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 3234 15852 3240 15904
rect 3292 15892 3298 15904
rect 4264 15892 4292 15923
rect 4801 15895 4859 15901
rect 4801 15892 4813 15895
rect 3292 15864 4813 15892
rect 3292 15852 3298 15864
rect 4801 15861 4813 15864
rect 4847 15861 4859 15895
rect 4801 15855 4859 15861
rect 8110 15852 8116 15904
rect 8168 15892 8174 15904
rect 8665 15895 8723 15901
rect 8665 15892 8677 15895
rect 8168 15864 8677 15892
rect 8168 15852 8174 15864
rect 8665 15861 8677 15864
rect 8711 15861 8723 15895
rect 9968 15892 9996 15923
rect 10502 15892 10508 15904
rect 9968 15864 10508 15892
rect 8665 15855 8723 15861
rect 10502 15852 10508 15864
rect 10560 15852 10566 15904
rect 13556 15892 13584 15923
rect 13722 15892 13728 15904
rect 13556 15864 13728 15892
rect 13722 15852 13728 15864
rect 13780 15852 13786 15904
rect 1104 15802 16836 15824
rect 1104 15750 6226 15802
rect 6278 15750 6290 15802
rect 6342 15750 6354 15802
rect 6406 15750 6418 15802
rect 6470 15750 11470 15802
rect 11522 15750 11534 15802
rect 11586 15750 11598 15802
rect 11650 15750 11662 15802
rect 11714 15750 16836 15802
rect 1104 15728 16836 15750
rect 2498 15688 2504 15700
rect 2240 15660 2504 15688
rect 2240 15629 2268 15660
rect 2498 15648 2504 15660
rect 2556 15688 2562 15700
rect 2777 15691 2835 15697
rect 2777 15688 2789 15691
rect 2556 15660 2789 15688
rect 2556 15648 2562 15660
rect 2777 15657 2789 15660
rect 2823 15657 2835 15691
rect 2777 15651 2835 15657
rect 8570 15648 8576 15700
rect 8628 15688 8634 15700
rect 8665 15691 8723 15697
rect 8665 15688 8677 15691
rect 8628 15660 8677 15688
rect 8628 15648 8634 15660
rect 8665 15657 8677 15660
rect 8711 15657 8723 15691
rect 8665 15651 8723 15657
rect 13722 15648 13728 15700
rect 13780 15688 13786 15700
rect 14185 15691 14243 15697
rect 14185 15688 14197 15691
rect 13780 15660 14197 15688
rect 13780 15648 13786 15660
rect 14185 15657 14197 15660
rect 14231 15657 14243 15691
rect 14185 15651 14243 15657
rect 16301 15691 16359 15697
rect 16301 15657 16313 15691
rect 16347 15657 16359 15691
rect 16301 15651 16359 15657
rect 2225 15623 2283 15629
rect 2225 15589 2237 15623
rect 2271 15589 2283 15623
rect 3234 15620 3240 15632
rect 3195 15592 3240 15620
rect 2225 15583 2283 15589
rect 3234 15580 3240 15592
rect 3292 15580 3298 15632
rect 10502 15580 10508 15632
rect 10560 15620 10566 15632
rect 11701 15623 11759 15629
rect 11701 15620 11713 15623
rect 10560 15592 11713 15620
rect 10560 15580 10566 15592
rect 11701 15589 11713 15592
rect 11747 15589 11759 15623
rect 11701 15583 11759 15589
rect 13265 15623 13323 15629
rect 13265 15589 13277 15623
rect 13311 15620 13323 15623
rect 16316 15620 16344 15651
rect 13311 15592 16344 15620
rect 13311 15589 13323 15592
rect 13265 15583 13323 15589
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 1762 15552 1768 15564
rect 1723 15524 1768 15552
rect 1762 15512 1768 15524
rect 1820 15512 1826 15564
rect 2314 15552 2320 15564
rect 2227 15524 2320 15552
rect 2314 15512 2320 15524
rect 2372 15552 2378 15564
rect 3053 15555 3111 15561
rect 3053 15552 3065 15555
rect 2372 15524 3065 15552
rect 2372 15512 2378 15524
rect 3053 15521 3065 15524
rect 3099 15552 3111 15555
rect 3605 15555 3663 15561
rect 3605 15552 3617 15555
rect 3099 15524 3617 15552
rect 3099 15521 3111 15524
rect 3053 15515 3111 15521
rect 3605 15521 3617 15524
rect 3651 15521 3663 15555
rect 8570 15552 8576 15564
rect 8531 15524 8576 15552
rect 3605 15515 3663 15521
rect 8570 15512 8576 15524
rect 8628 15512 8634 15564
rect 13354 15552 13360 15564
rect 13315 15524 13360 15552
rect 13354 15512 13360 15524
rect 13412 15512 13418 15564
rect 13446 15512 13452 15564
rect 13504 15552 13510 15564
rect 13817 15555 13875 15561
rect 13817 15552 13829 15555
rect 13504 15524 13829 15552
rect 13504 15512 13510 15524
rect 1780 15484 1808 15512
rect 2409 15487 2467 15493
rect 2409 15484 2421 15487
rect 1780 15456 2421 15484
rect 2409 15453 2421 15456
rect 2455 15453 2467 15487
rect 2409 15447 2467 15453
rect 12434 15444 12440 15496
rect 12492 15484 12498 15496
rect 13081 15487 13139 15493
rect 13081 15484 13093 15487
rect 12492 15456 13093 15484
rect 12492 15444 12498 15456
rect 13081 15453 13093 15456
rect 13127 15484 13139 15487
rect 13170 15484 13176 15496
rect 13127 15456 13176 15484
rect 13127 15453 13139 15456
rect 13081 15447 13139 15453
rect 13170 15444 13176 15456
rect 13228 15444 13234 15496
rect 2777 15419 2835 15425
rect 2777 15385 2789 15419
rect 2823 15416 2835 15419
rect 3421 15419 3479 15425
rect 3421 15416 3433 15419
rect 2823 15388 3433 15416
rect 2823 15385 2835 15388
rect 2777 15379 2835 15385
rect 3421 15385 3433 15388
rect 3467 15385 3479 15419
rect 3421 15379 3479 15385
rect 11885 15419 11943 15425
rect 11885 15385 11897 15419
rect 11931 15416 11943 15419
rect 13630 15416 13636 15428
rect 11931 15388 13636 15416
rect 11931 15385 11943 15388
rect 11885 15379 11943 15385
rect 13630 15376 13636 15388
rect 13688 15376 13694 15428
rect 13740 15425 13768 15524
rect 13817 15521 13829 15524
rect 13863 15521 13875 15555
rect 13817 15515 13875 15521
rect 13906 15512 13912 15564
rect 13964 15552 13970 15564
rect 14553 15555 14611 15561
rect 14553 15552 14565 15555
rect 13964 15524 14565 15552
rect 13964 15512 13970 15524
rect 14553 15521 14565 15524
rect 14599 15521 14611 15555
rect 15746 15552 15752 15564
rect 15707 15524 15752 15552
rect 14553 15515 14611 15521
rect 15746 15512 15752 15524
rect 15804 15512 15810 15564
rect 16482 15552 16488 15564
rect 16443 15524 16488 15552
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 13725 15419 13783 15425
rect 13725 15385 13737 15419
rect 13771 15385 13783 15419
rect 13725 15379 13783 15385
rect 14185 15419 14243 15425
rect 14185 15385 14197 15419
rect 14231 15416 14243 15419
rect 14369 15419 14427 15425
rect 14369 15416 14381 15419
rect 14231 15388 14381 15416
rect 14231 15385 14243 15388
rect 14185 15379 14243 15385
rect 14369 15385 14381 15388
rect 14415 15385 14427 15419
rect 14369 15379 14427 15385
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15348 1639 15351
rect 4430 15348 4436 15360
rect 1627 15320 4436 15348
rect 1627 15317 1639 15320
rect 1581 15311 1639 15317
rect 4430 15308 4436 15320
rect 4488 15308 4494 15360
rect 15838 15348 15844 15360
rect 15799 15320 15844 15348
rect 15838 15308 15844 15320
rect 15896 15308 15902 15360
rect 1104 15258 16836 15280
rect 1104 15206 3604 15258
rect 3656 15206 3668 15258
rect 3720 15206 3732 15258
rect 3784 15206 3796 15258
rect 3848 15206 8848 15258
rect 8900 15206 8912 15258
rect 8964 15206 8976 15258
rect 9028 15206 9040 15258
rect 9092 15206 14092 15258
rect 14144 15206 14156 15258
rect 14208 15206 14220 15258
rect 14272 15206 14284 15258
rect 14336 15206 16836 15258
rect 1104 15184 16836 15206
rect 3970 15144 3976 15156
rect 3931 15116 3976 15144
rect 3970 15104 3976 15116
rect 4028 15104 4034 15156
rect 7193 15147 7251 15153
rect 7193 15113 7205 15147
rect 7239 15144 7251 15147
rect 9490 15144 9496 15156
rect 7239 15116 9496 15144
rect 7239 15113 7251 15116
rect 7193 15107 7251 15113
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 13906 15104 13912 15156
rect 13964 15144 13970 15156
rect 14093 15147 14151 15153
rect 14093 15144 14105 15147
rect 13964 15116 14105 15144
rect 13964 15104 13970 15116
rect 14093 15113 14105 15116
rect 14139 15113 14151 15147
rect 14093 15107 14151 15113
rect 15657 15147 15715 15153
rect 15657 15113 15669 15147
rect 15703 15144 15715 15147
rect 15746 15144 15752 15156
rect 15703 15116 15752 15144
rect 15703 15113 15715 15116
rect 15657 15107 15715 15113
rect 15746 15104 15752 15116
rect 15804 15104 15810 15156
rect 4062 15036 4068 15088
rect 4120 15076 4126 15088
rect 5902 15076 5908 15088
rect 4120 15048 5908 15076
rect 4120 15036 4126 15048
rect 2406 15008 2412 15020
rect 2240 14980 2412 15008
rect 1486 14940 1492 14952
rect 1447 14912 1492 14940
rect 1486 14900 1492 14912
rect 1544 14900 1550 14952
rect 2240 14949 2268 14980
rect 2406 14968 2412 14980
rect 2464 14968 2470 15020
rect 4430 15008 4436 15020
rect 4391 14980 4436 15008
rect 4430 14968 4436 14980
rect 4488 14968 4494 15020
rect 4522 14968 4528 15020
rect 4580 15008 4586 15020
rect 4632 15017 4660 15048
rect 5902 15036 5908 15048
rect 5960 15076 5966 15088
rect 5960 15048 6592 15076
rect 5960 15036 5966 15048
rect 6564 15020 6592 15048
rect 10042 15036 10048 15088
rect 10100 15076 10106 15088
rect 11701 15079 11759 15085
rect 11701 15076 11713 15079
rect 10100 15048 11713 15076
rect 10100 15036 10106 15048
rect 11701 15045 11713 15048
rect 11747 15045 11759 15079
rect 11701 15039 11759 15045
rect 16117 15079 16175 15085
rect 16117 15045 16129 15079
rect 16163 15076 16175 15079
rect 16209 15079 16267 15085
rect 16209 15076 16221 15079
rect 16163 15048 16221 15076
rect 16163 15045 16175 15048
rect 16117 15039 16175 15045
rect 16209 15045 16221 15048
rect 16255 15045 16267 15079
rect 16209 15039 16267 15045
rect 4617 15011 4675 15017
rect 4617 15008 4629 15011
rect 4580 14980 4629 15008
rect 4580 14968 4586 14980
rect 4617 14977 4629 14980
rect 4663 14977 4675 15011
rect 4617 14971 4675 14977
rect 5810 14968 5816 15020
rect 5868 14968 5874 15020
rect 6546 15008 6552 15020
rect 6507 14980 6552 15008
rect 6546 14968 6552 14980
rect 6604 14968 6610 15020
rect 12158 15008 12164 15020
rect 12119 14980 12164 15008
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 12345 15011 12403 15017
rect 12345 14977 12357 15011
rect 12391 15008 12403 15011
rect 12434 15008 12440 15020
rect 12391 14980 12440 15008
rect 12391 14977 12403 14980
rect 12345 14971 12403 14977
rect 12434 14968 12440 14980
rect 12492 14968 12498 15020
rect 15749 15011 15807 15017
rect 15749 15008 15761 15011
rect 15212 14980 15761 15008
rect 2225 14943 2283 14949
rect 2225 14909 2237 14943
rect 2271 14909 2283 14943
rect 2498 14940 2504 14952
rect 2459 14912 2504 14940
rect 2225 14903 2283 14909
rect 2498 14900 2504 14912
rect 2556 14900 2562 14952
rect 5828 14940 5856 14968
rect 15212 14952 15240 14980
rect 15749 14977 15761 14980
rect 15795 14977 15807 15011
rect 15749 14971 15807 14977
rect 6733 14943 6791 14949
rect 6733 14940 6745 14943
rect 5828 14912 6745 14940
rect 6733 14909 6745 14912
rect 6779 14909 6791 14943
rect 6733 14903 6791 14909
rect 6914 14900 6920 14952
rect 6972 14940 6978 14952
rect 6972 14912 12112 14940
rect 6972 14900 6978 14912
rect 2314 14832 2320 14884
rect 2372 14872 2378 14884
rect 2409 14875 2467 14881
rect 2409 14872 2421 14875
rect 2372 14844 2421 14872
rect 2372 14832 2378 14844
rect 2409 14841 2421 14844
rect 2455 14841 2467 14875
rect 2409 14835 2467 14841
rect 4341 14875 4399 14881
rect 4341 14841 4353 14875
rect 4387 14872 4399 14875
rect 5445 14875 5503 14881
rect 5445 14872 5457 14875
rect 4387 14844 5457 14872
rect 4387 14841 4399 14844
rect 4341 14835 4399 14841
rect 5445 14841 5457 14844
rect 5491 14841 5503 14875
rect 5445 14835 5503 14841
rect 5534 14832 5540 14884
rect 5592 14872 5598 14884
rect 5629 14875 5687 14881
rect 5629 14872 5641 14875
rect 5592 14844 5641 14872
rect 5592 14832 5598 14844
rect 5629 14841 5641 14844
rect 5675 14841 5687 14875
rect 5629 14835 5687 14841
rect 5813 14875 5871 14881
rect 5813 14841 5825 14875
rect 5859 14872 5871 14875
rect 5905 14875 5963 14881
rect 5905 14872 5917 14875
rect 5859 14844 5917 14872
rect 5859 14841 5871 14844
rect 5813 14835 5871 14841
rect 5905 14841 5917 14844
rect 5951 14841 5963 14875
rect 5905 14835 5963 14841
rect 2590 14764 2596 14816
rect 2648 14804 2654 14816
rect 2648 14776 2693 14804
rect 2648 14764 2654 14776
rect 5350 14764 5356 14816
rect 5408 14804 5414 14816
rect 5920 14804 5948 14835
rect 5994 14832 6000 14884
rect 6052 14872 6058 14884
rect 6089 14875 6147 14881
rect 6089 14872 6101 14875
rect 6052 14844 6101 14872
rect 6052 14832 6058 14844
rect 6089 14841 6101 14844
rect 6135 14841 6147 14875
rect 6089 14835 6147 14841
rect 6273 14875 6331 14881
rect 6273 14841 6285 14875
rect 6319 14872 6331 14875
rect 6825 14875 6883 14881
rect 6825 14872 6837 14875
rect 6319 14844 6837 14872
rect 6319 14841 6331 14844
rect 6273 14835 6331 14841
rect 6825 14841 6837 14844
rect 6871 14841 6883 14875
rect 6825 14835 6883 14841
rect 11330 14832 11336 14884
rect 11388 14872 11394 14884
rect 11517 14875 11575 14881
rect 11517 14872 11529 14875
rect 11388 14844 11529 14872
rect 11388 14832 11394 14844
rect 11517 14841 11529 14844
rect 11563 14841 11575 14875
rect 11517 14835 11575 14841
rect 6914 14804 6920 14816
rect 5408 14776 6920 14804
rect 5408 14764 5414 14776
rect 6914 14764 6920 14776
rect 6972 14764 6978 14816
rect 10410 14764 10416 14816
rect 10468 14804 10474 14816
rect 12084 14813 12112 14912
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 15105 14943 15163 14949
rect 13688 14912 15056 14940
rect 13688 14900 13694 14912
rect 13906 14832 13912 14884
rect 13964 14872 13970 14884
rect 14001 14875 14059 14881
rect 14001 14872 14013 14875
rect 13964 14844 14013 14872
rect 13964 14832 13970 14844
rect 14001 14841 14013 14844
rect 14047 14841 14059 14875
rect 15028 14872 15056 14912
rect 15105 14909 15117 14943
rect 15151 14940 15163 14943
rect 15194 14940 15200 14952
rect 15151 14912 15200 14940
rect 15151 14909 15163 14912
rect 15105 14903 15163 14909
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 15657 14943 15715 14949
rect 15657 14909 15669 14943
rect 15703 14940 15715 14943
rect 16393 14943 16451 14949
rect 16393 14940 16405 14943
rect 15703 14912 16405 14940
rect 15703 14909 15715 14912
rect 15657 14903 15715 14909
rect 16393 14909 16405 14912
rect 16439 14909 16451 14943
rect 16393 14903 16451 14909
rect 15672 14872 15700 14903
rect 15028 14844 15700 14872
rect 14001 14835 14059 14841
rect 11425 14807 11483 14813
rect 11425 14804 11437 14807
rect 10468 14776 11437 14804
rect 10468 14764 10474 14776
rect 11425 14773 11437 14776
rect 11471 14773 11483 14807
rect 11425 14767 11483 14773
rect 12069 14807 12127 14813
rect 12069 14773 12081 14807
rect 12115 14804 12127 14807
rect 12342 14804 12348 14816
rect 12115 14776 12348 14804
rect 12115 14773 12127 14776
rect 12069 14767 12127 14773
rect 12342 14764 12348 14776
rect 12400 14764 12406 14816
rect 15746 14764 15752 14816
rect 15804 14804 15810 14816
rect 16117 14807 16175 14813
rect 16117 14804 16129 14807
rect 15804 14776 16129 14804
rect 15804 14764 15810 14776
rect 16117 14773 16129 14776
rect 16163 14773 16175 14807
rect 16117 14767 16175 14773
rect 1104 14714 16836 14736
rect 1104 14662 6226 14714
rect 6278 14662 6290 14714
rect 6342 14662 6354 14714
rect 6406 14662 6418 14714
rect 6470 14662 11470 14714
rect 11522 14662 11534 14714
rect 11586 14662 11598 14714
rect 11650 14662 11662 14714
rect 11714 14662 16836 14714
rect 1104 14640 16836 14662
rect 4338 14600 4344 14612
rect 4299 14572 4344 14600
rect 4338 14560 4344 14572
rect 4396 14560 4402 14612
rect 6086 14560 6092 14612
rect 6144 14600 6150 14612
rect 6365 14603 6423 14609
rect 6365 14600 6377 14603
rect 6144 14572 6377 14600
rect 6144 14560 6150 14572
rect 6365 14569 6377 14572
rect 6411 14569 6423 14603
rect 6365 14563 6423 14569
rect 8481 14603 8539 14609
rect 8481 14569 8493 14603
rect 8527 14600 8539 14603
rect 8570 14600 8576 14612
rect 8527 14572 8576 14600
rect 8527 14569 8539 14572
rect 8481 14563 8539 14569
rect 5534 14492 5540 14544
rect 5592 14532 5598 14544
rect 7929 14535 7987 14541
rect 5592 14504 6776 14532
rect 5592 14492 5598 14504
rect 2590 14464 2596 14476
rect 2551 14436 2596 14464
rect 2590 14424 2596 14436
rect 2648 14424 2654 14476
rect 4249 14467 4307 14473
rect 4249 14433 4261 14467
rect 4295 14464 4307 14467
rect 5721 14467 5779 14473
rect 5721 14464 5733 14467
rect 4295 14436 5733 14464
rect 4295 14433 4307 14436
rect 4249 14427 4307 14433
rect 5721 14433 5733 14436
rect 5767 14433 5779 14467
rect 5721 14427 5779 14433
rect 5905 14467 5963 14473
rect 5905 14433 5917 14467
rect 5951 14433 5963 14467
rect 5905 14427 5963 14433
rect 1486 14356 1492 14408
rect 1544 14396 1550 14408
rect 1857 14399 1915 14405
rect 1857 14396 1869 14399
rect 1544 14368 1869 14396
rect 1544 14356 1550 14368
rect 1857 14365 1869 14368
rect 1903 14396 1915 14399
rect 2314 14396 2320 14408
rect 1903 14368 2320 14396
rect 1903 14365 1915 14368
rect 1857 14359 1915 14365
rect 2314 14356 2320 14368
rect 2372 14356 2378 14408
rect 2406 14356 2412 14408
rect 2464 14396 2470 14408
rect 2501 14399 2559 14405
rect 2501 14396 2513 14399
rect 2464 14368 2513 14396
rect 2464 14356 2470 14368
rect 2501 14365 2513 14368
rect 2547 14365 2559 14399
rect 4522 14396 4528 14408
rect 4483 14368 4528 14396
rect 2501 14359 2559 14365
rect 4522 14356 4528 14368
rect 4580 14356 4586 14408
rect 5626 14356 5632 14408
rect 5684 14396 5690 14408
rect 5920 14396 5948 14427
rect 6178 14424 6184 14476
rect 6236 14464 6242 14476
rect 6748 14473 6776 14504
rect 7929 14501 7941 14535
rect 7975 14532 7987 14535
rect 8496 14532 8524 14563
rect 8570 14560 8576 14572
rect 8628 14560 8634 14612
rect 12253 14603 12311 14609
rect 9232 14572 11284 14600
rect 7975 14504 8524 14532
rect 7975 14501 7987 14504
rect 7929 14495 7987 14501
rect 9232 14476 9260 14572
rect 6549 14467 6607 14473
rect 6236 14436 6281 14464
rect 6236 14424 6242 14436
rect 6549 14433 6561 14467
rect 6595 14433 6607 14467
rect 6549 14427 6607 14433
rect 6733 14467 6791 14473
rect 6733 14433 6745 14467
rect 6779 14433 6791 14467
rect 6733 14427 6791 14433
rect 6825 14467 6883 14473
rect 6825 14433 6837 14467
rect 6871 14464 6883 14467
rect 6914 14464 6920 14476
rect 6871 14436 6920 14464
rect 6871 14433 6883 14436
rect 6825 14427 6883 14433
rect 6564 14396 6592 14427
rect 6914 14424 6920 14436
rect 6972 14424 6978 14476
rect 7469 14467 7527 14473
rect 7469 14433 7481 14467
rect 7515 14464 7527 14467
rect 7558 14464 7564 14476
rect 7515 14436 7564 14464
rect 7515 14433 7527 14436
rect 7469 14427 7527 14433
rect 7558 14424 7564 14436
rect 7616 14424 7622 14476
rect 8018 14464 8024 14476
rect 7979 14436 8024 14464
rect 8018 14424 8024 14436
rect 8076 14424 8082 14476
rect 8294 14424 8300 14476
rect 8352 14464 8358 14476
rect 8573 14467 8631 14473
rect 8573 14464 8585 14467
rect 8352 14436 8585 14464
rect 8352 14424 8358 14436
rect 8573 14433 8585 14436
rect 8619 14433 8631 14467
rect 9214 14464 9220 14476
rect 9175 14436 9220 14464
rect 8573 14427 8631 14433
rect 9214 14424 9220 14436
rect 9272 14424 9278 14476
rect 9769 14467 9827 14473
rect 9769 14433 9781 14467
rect 9815 14464 9827 14467
rect 10042 14464 10048 14476
rect 9815 14436 10048 14464
rect 9815 14433 9827 14436
rect 9769 14427 9827 14433
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 10410 14464 10416 14476
rect 10371 14436 10416 14464
rect 10410 14424 10416 14436
rect 10468 14424 10474 14476
rect 11256 14473 11284 14572
rect 12253 14569 12265 14603
rect 12299 14569 12311 14603
rect 12253 14563 12311 14569
rect 10689 14467 10747 14473
rect 10689 14433 10701 14467
rect 10735 14433 10747 14467
rect 10689 14427 10747 14433
rect 11241 14467 11299 14473
rect 11241 14433 11253 14467
rect 11287 14433 11299 14467
rect 11241 14427 11299 14433
rect 11793 14467 11851 14473
rect 11793 14433 11805 14467
rect 11839 14464 11851 14467
rect 11882 14464 11888 14476
rect 11839 14436 11888 14464
rect 11839 14433 11851 14436
rect 11793 14427 11851 14433
rect 5684 14368 6592 14396
rect 5684 14356 5690 14368
rect 5994 14328 6000 14340
rect 5955 14300 6000 14328
rect 5994 14288 6000 14300
rect 6052 14288 6058 14340
rect 6089 14331 6147 14337
rect 6089 14297 6101 14331
rect 6135 14297 6147 14331
rect 6564 14328 6592 14368
rect 6638 14356 6644 14408
rect 6696 14396 6702 14408
rect 7576 14396 7604 14424
rect 8113 14399 8171 14405
rect 8113 14396 8125 14399
rect 6696 14368 6741 14396
rect 7576 14368 8125 14396
rect 6696 14356 6702 14368
rect 8113 14365 8125 14368
rect 8159 14365 8171 14399
rect 10704 14396 10732 14427
rect 8113 14359 8171 14365
rect 10428 14368 10732 14396
rect 6914 14328 6920 14340
rect 6564 14300 6920 14328
rect 6089 14291 6147 14297
rect 3142 14220 3148 14272
rect 3200 14260 3206 14272
rect 3881 14263 3939 14269
rect 3881 14260 3893 14263
rect 3200 14232 3893 14260
rect 3200 14220 3206 14232
rect 3881 14229 3893 14232
rect 3927 14229 3939 14263
rect 3881 14223 3939 14229
rect 5902 14220 5908 14272
rect 5960 14260 5966 14272
rect 6104 14260 6132 14291
rect 6914 14288 6920 14300
rect 6972 14288 6978 14340
rect 8481 14331 8539 14337
rect 8481 14297 8493 14331
rect 8527 14328 8539 14331
rect 8665 14331 8723 14337
rect 8665 14328 8677 14331
rect 8527 14300 8677 14328
rect 8527 14297 8539 14300
rect 8481 14291 8539 14297
rect 8665 14297 8677 14300
rect 8711 14297 8723 14331
rect 8665 14291 8723 14297
rect 10428 14269 10456 14368
rect 5960 14232 6132 14260
rect 9217 14263 9275 14269
rect 5960 14220 5966 14232
rect 9217 14229 9229 14263
rect 9263 14260 9275 14263
rect 10413 14263 10471 14269
rect 10413 14260 10425 14263
rect 9263 14232 10425 14260
rect 9263 14229 9275 14232
rect 9217 14223 9275 14229
rect 10413 14229 10425 14232
rect 10459 14229 10471 14263
rect 10594 14260 10600 14272
rect 10555 14232 10600 14260
rect 10413 14223 10471 14229
rect 10594 14220 10600 14232
rect 10652 14220 10658 14272
rect 11256 14260 11284 14427
rect 11882 14424 11888 14436
rect 11940 14424 11946 14476
rect 11330 14356 11336 14408
rect 11388 14396 11394 14408
rect 11425 14399 11483 14405
rect 11425 14396 11437 14399
rect 11388 14368 11437 14396
rect 11388 14356 11394 14368
rect 11425 14365 11437 14368
rect 11471 14396 11483 14399
rect 12268 14396 12296 14563
rect 12529 14467 12587 14473
rect 12529 14433 12541 14467
rect 12575 14433 12587 14467
rect 16482 14464 16488 14476
rect 16443 14436 16488 14464
rect 12529 14427 12587 14433
rect 11471 14368 12296 14396
rect 11471 14365 11483 14368
rect 11425 14359 11483 14365
rect 12253 14331 12311 14337
rect 12253 14297 12265 14331
rect 12299 14328 12311 14331
rect 12345 14331 12403 14337
rect 12345 14328 12357 14331
rect 12299 14300 12357 14328
rect 12299 14297 12311 14300
rect 12253 14291 12311 14297
rect 12345 14297 12357 14300
rect 12391 14297 12403 14331
rect 12345 14291 12403 14297
rect 12544 14260 12572 14427
rect 16482 14424 16488 14436
rect 16540 14424 16546 14476
rect 16298 14260 16304 14272
rect 11256 14232 12572 14260
rect 16259 14232 16304 14260
rect 16298 14220 16304 14232
rect 16356 14220 16362 14272
rect 1104 14170 16836 14192
rect 1104 14118 3604 14170
rect 3656 14118 3668 14170
rect 3720 14118 3732 14170
rect 3784 14118 3796 14170
rect 3848 14118 8848 14170
rect 8900 14118 8912 14170
rect 8964 14118 8976 14170
rect 9028 14118 9040 14170
rect 9092 14118 14092 14170
rect 14144 14118 14156 14170
rect 14208 14118 14220 14170
rect 14272 14118 14284 14170
rect 14336 14118 16836 14170
rect 1104 14096 16836 14118
rect 6181 14059 6239 14065
rect 6181 14025 6193 14059
rect 6227 14056 6239 14059
rect 9214 14056 9220 14068
rect 6227 14028 9220 14056
rect 6227 14025 6239 14028
rect 6181 14019 6239 14025
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 13633 14059 13691 14065
rect 13633 14025 13645 14059
rect 13679 14056 13691 14059
rect 13906 14056 13912 14068
rect 13679 14028 13912 14056
rect 13679 14025 13691 14028
rect 13633 14019 13691 14025
rect 13906 14016 13912 14028
rect 13964 14056 13970 14068
rect 14093 14059 14151 14065
rect 14093 14056 14105 14059
rect 13964 14028 14105 14056
rect 13964 14016 13970 14028
rect 14093 14025 14105 14028
rect 14139 14025 14151 14059
rect 14093 14019 14151 14025
rect 14826 14016 14832 14068
rect 14884 14056 14890 14068
rect 16117 14059 16175 14065
rect 16117 14056 16129 14059
rect 14884 14028 16129 14056
rect 14884 14016 14890 14028
rect 16117 14025 16129 14028
rect 16163 14025 16175 14059
rect 16117 14019 16175 14025
rect 7837 13991 7895 13997
rect 7837 13957 7849 13991
rect 7883 13988 7895 13991
rect 8202 13988 8208 14000
rect 7883 13960 8208 13988
rect 7883 13957 7895 13960
rect 7837 13951 7895 13957
rect 8202 13948 8208 13960
rect 8260 13948 8266 14000
rect 8297 13991 8355 13997
rect 8297 13957 8309 13991
rect 8343 13988 8355 13991
rect 8389 13991 8447 13997
rect 8389 13988 8401 13991
rect 8343 13960 8401 13988
rect 8343 13957 8355 13960
rect 8297 13951 8355 13957
rect 8389 13957 8401 13960
rect 8435 13957 8447 13991
rect 8389 13951 8447 13957
rect 13722 13948 13728 14000
rect 13780 13988 13786 14000
rect 13780 13960 14964 13988
rect 13780 13948 13786 13960
rect 7929 13923 7987 13929
rect 7929 13920 7941 13923
rect 7300 13892 7941 13920
rect 7300 13864 7328 13892
rect 7929 13889 7941 13892
rect 7975 13889 7987 13923
rect 7929 13883 7987 13889
rect 13096 13892 13768 13920
rect 5626 13812 5632 13864
rect 5684 13852 5690 13864
rect 6089 13855 6147 13861
rect 6089 13852 6101 13855
rect 5684 13824 6101 13852
rect 5684 13812 5690 13824
rect 6089 13821 6101 13824
rect 6135 13821 6147 13855
rect 7282 13852 7288 13864
rect 7243 13824 7288 13852
rect 6089 13815 6147 13821
rect 7282 13812 7288 13824
rect 7340 13812 7346 13864
rect 7837 13855 7895 13861
rect 7837 13821 7849 13855
rect 7883 13852 7895 13855
rect 8018 13852 8024 13864
rect 7883 13824 8024 13852
rect 7883 13821 7895 13824
rect 7837 13815 7895 13821
rect 8018 13812 8024 13824
rect 8076 13852 8082 13864
rect 8573 13855 8631 13861
rect 8573 13852 8585 13855
rect 8076 13824 8585 13852
rect 8076 13812 8082 13824
rect 8573 13821 8585 13824
rect 8619 13852 8631 13855
rect 10594 13852 10600 13864
rect 8619 13824 10600 13852
rect 8619 13821 8631 13824
rect 8573 13815 8631 13821
rect 10594 13812 10600 13824
rect 10652 13812 10658 13864
rect 11790 13852 11796 13864
rect 11751 13824 11796 13852
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 11885 13855 11943 13861
rect 11885 13821 11897 13855
rect 11931 13852 11943 13855
rect 12066 13852 12072 13864
rect 11931 13824 12072 13852
rect 11931 13821 11943 13824
rect 11885 13815 11943 13821
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 13096 13861 13124 13892
rect 13740 13864 13768 13892
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 13633 13855 13691 13861
rect 13633 13821 13645 13855
rect 13679 13821 13691 13855
rect 13633 13815 13691 13821
rect 13648 13784 13676 13815
rect 13722 13812 13728 13864
rect 13780 13852 13786 13864
rect 14090 13852 14096 13864
rect 13780 13824 13825 13852
rect 14051 13824 14096 13852
rect 13780 13812 13786 13824
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 14936 13861 14964 13960
rect 15838 13948 15844 14000
rect 15896 13988 15902 14000
rect 15933 13991 15991 13997
rect 15933 13988 15945 13991
rect 15896 13960 15945 13988
rect 15896 13948 15902 13960
rect 15933 13957 15945 13960
rect 15979 13957 15991 13991
rect 15933 13951 15991 13957
rect 15105 13923 15163 13929
rect 15105 13889 15117 13923
rect 15151 13920 15163 13923
rect 15151 13892 16252 13920
rect 15151 13889 15163 13892
rect 15105 13883 15163 13889
rect 14921 13855 14979 13861
rect 14921 13821 14933 13855
rect 14967 13821 14979 13855
rect 14921 13815 14979 13821
rect 15378 13812 15384 13864
rect 15436 13852 15442 13864
rect 15473 13855 15531 13861
rect 15473 13852 15485 13855
rect 15436 13824 15485 13852
rect 15436 13812 15442 13824
rect 15473 13821 15485 13824
rect 15519 13852 15531 13855
rect 15565 13855 15623 13861
rect 15565 13852 15577 13855
rect 15519 13824 15577 13852
rect 15519 13821 15531 13824
rect 15473 13815 15531 13821
rect 15565 13821 15577 13824
rect 15611 13821 15623 13855
rect 15565 13815 15623 13821
rect 14826 13784 14832 13796
rect 13648 13756 14832 13784
rect 14826 13744 14832 13756
rect 14884 13744 14890 13796
rect 4246 13676 4252 13728
rect 4304 13716 4310 13728
rect 4709 13719 4767 13725
rect 4709 13716 4721 13719
rect 4304 13688 4721 13716
rect 4304 13676 4310 13688
rect 4709 13685 4721 13688
rect 4755 13685 4767 13719
rect 4709 13679 4767 13685
rect 4798 13676 4804 13728
rect 4856 13716 4862 13728
rect 8294 13716 8300 13728
rect 4856 13688 4901 13716
rect 8255 13688 8300 13716
rect 4856 13676 4862 13688
rect 8294 13676 8300 13688
rect 8352 13676 8358 13728
rect 12066 13716 12072 13728
rect 12027 13688 12072 13716
rect 12066 13676 12072 13688
rect 12124 13676 12130 13728
rect 15948 13725 15976 13892
rect 16224 13861 16252 13892
rect 16209 13855 16267 13861
rect 16209 13821 16221 13855
rect 16255 13821 16267 13855
rect 16209 13815 16267 13821
rect 15933 13719 15991 13725
rect 15933 13685 15945 13719
rect 15979 13685 15991 13719
rect 15933 13679 15991 13685
rect 1104 13626 16836 13648
rect 1104 13574 6226 13626
rect 6278 13574 6290 13626
rect 6342 13574 6354 13626
rect 6406 13574 6418 13626
rect 6470 13574 11470 13626
rect 11522 13574 11534 13626
rect 11586 13574 11598 13626
rect 11650 13574 11662 13626
rect 11714 13574 16836 13626
rect 1104 13552 16836 13574
rect 2869 13515 2927 13521
rect 2869 13512 2881 13515
rect 2746 13484 2881 13512
rect 2317 13447 2375 13453
rect 2317 13413 2329 13447
rect 2363 13444 2375 13447
rect 2746 13444 2774 13484
rect 2869 13481 2881 13484
rect 2915 13512 2927 13515
rect 3237 13515 3295 13521
rect 3237 13512 3249 13515
rect 2915 13484 3249 13512
rect 2915 13481 2927 13484
rect 2869 13475 2927 13481
rect 3237 13481 3249 13484
rect 3283 13481 3295 13515
rect 4847 13515 4905 13521
rect 4847 13512 4859 13515
rect 3237 13475 3295 13481
rect 4264 13484 4859 13512
rect 4264 13456 4292 13484
rect 4847 13481 4859 13484
rect 4893 13481 4905 13515
rect 4847 13475 4905 13481
rect 5718 13472 5724 13524
rect 5776 13512 5782 13524
rect 5813 13515 5871 13521
rect 5813 13512 5825 13515
rect 5776 13484 5825 13512
rect 5776 13472 5782 13484
rect 5813 13481 5825 13484
rect 5859 13481 5871 13515
rect 8662 13512 8668 13524
rect 8623 13484 8668 13512
rect 5813 13475 5871 13481
rect 8662 13472 8668 13484
rect 8720 13472 8726 13524
rect 11793 13515 11851 13521
rect 11793 13481 11805 13515
rect 11839 13512 11851 13515
rect 11882 13512 11888 13524
rect 11839 13484 11888 13512
rect 11839 13481 11851 13484
rect 11793 13475 11851 13481
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 12066 13472 12072 13524
rect 12124 13512 12130 13524
rect 12161 13515 12219 13521
rect 12161 13512 12173 13515
rect 12124 13484 12173 13512
rect 12124 13472 12130 13484
rect 12161 13481 12173 13484
rect 12207 13481 12219 13515
rect 14090 13512 14096 13524
rect 14051 13484 14096 13512
rect 12161 13475 12219 13481
rect 14090 13472 14096 13484
rect 14148 13472 14154 13524
rect 2363 13416 2774 13444
rect 3973 13447 4031 13453
rect 2363 13413 2375 13416
rect 2317 13407 2375 13413
rect 3973 13413 3985 13447
rect 4019 13444 4031 13447
rect 4246 13444 4252 13456
rect 4019 13416 4252 13444
rect 4019 13413 4031 13416
rect 3973 13407 4031 13413
rect 4246 13404 4252 13416
rect 4304 13404 4310 13456
rect 10303 13447 10361 13453
rect 10303 13444 10315 13447
rect 4356 13416 4844 13444
rect 1857 13379 1915 13385
rect 1857 13345 1869 13379
rect 1903 13345 1915 13379
rect 2406 13376 2412 13388
rect 2367 13348 2412 13376
rect 1857 13339 1915 13345
rect 1872 13308 1900 13339
rect 2406 13336 2412 13348
rect 2464 13376 2470 13388
rect 3145 13379 3203 13385
rect 3145 13376 3157 13379
rect 2464 13348 3157 13376
rect 2464 13336 2470 13348
rect 3145 13345 3157 13348
rect 3191 13345 3203 13379
rect 3878 13376 3884 13388
rect 3839 13348 3884 13376
rect 3145 13339 3203 13345
rect 3878 13336 3884 13348
rect 3936 13336 3942 13388
rect 2501 13311 2559 13317
rect 2501 13308 2513 13311
rect 1872 13280 2513 13308
rect 2501 13277 2513 13280
rect 2547 13308 2559 13311
rect 4356 13308 4384 13416
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13345 4491 13379
rect 4816 13376 4844 13416
rect 5000 13416 10315 13444
rect 5000 13376 5028 13416
rect 10303 13413 10315 13416
rect 10349 13413 10361 13447
rect 10303 13407 10361 13413
rect 10502 13404 10508 13456
rect 10560 13444 10566 13456
rect 10781 13447 10839 13453
rect 10781 13444 10793 13447
rect 10560 13416 10793 13444
rect 10560 13404 10566 13416
rect 10781 13413 10793 13416
rect 10827 13413 10839 13447
rect 10781 13407 10839 13413
rect 12253 13447 12311 13453
rect 12253 13413 12265 13447
rect 12299 13444 12311 13447
rect 16206 13444 16212 13456
rect 12299 13416 16212 13444
rect 12299 13413 12311 13416
rect 12253 13407 12311 13413
rect 16206 13404 16212 13416
rect 16264 13404 16270 13456
rect 5166 13376 5172 13388
rect 4816 13348 5028 13376
rect 5127 13348 5172 13376
rect 4433 13339 4491 13345
rect 2547 13280 4384 13308
rect 4448 13308 4476 13339
rect 5166 13336 5172 13348
rect 5224 13336 5230 13388
rect 5721 13379 5779 13385
rect 5721 13345 5733 13379
rect 5767 13376 5779 13379
rect 6454 13376 6460 13388
rect 5767 13348 6460 13376
rect 5767 13345 5779 13348
rect 5721 13339 5779 13345
rect 6454 13336 6460 13348
rect 6512 13336 6518 13388
rect 8570 13376 8576 13388
rect 8531 13348 8576 13376
rect 8570 13336 8576 13348
rect 8628 13336 8634 13388
rect 9769 13379 9827 13385
rect 9769 13345 9781 13379
rect 9815 13376 9827 13379
rect 9858 13376 9864 13388
rect 9815 13348 9864 13376
rect 9815 13345 9827 13348
rect 9769 13339 9827 13345
rect 9858 13336 9864 13348
rect 9916 13336 9922 13388
rect 10594 13376 10600 13388
rect 10555 13348 10600 13376
rect 10594 13336 10600 13348
rect 10652 13336 10658 13388
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 14001 13379 14059 13385
rect 14001 13376 14013 13379
rect 13964 13348 14013 13376
rect 13964 13336 13970 13348
rect 14001 13345 14013 13348
rect 14047 13345 14059 13379
rect 14001 13339 14059 13345
rect 4525 13311 4583 13317
rect 4525 13308 4537 13311
rect 4448 13280 4537 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 4525 13277 4537 13280
rect 4571 13308 4583 13311
rect 5994 13308 6000 13320
rect 4571 13280 5396 13308
rect 5907 13280 6000 13308
rect 4571 13277 4583 13280
rect 4525 13271 4583 13277
rect 5368 13249 5396 13280
rect 5994 13268 6000 13280
rect 6052 13308 6058 13320
rect 6546 13308 6552 13320
rect 6052 13280 6552 13308
rect 6052 13268 6058 13280
rect 6546 13268 6552 13280
rect 6604 13308 6610 13320
rect 8662 13308 8668 13320
rect 6604 13280 8668 13308
rect 6604 13268 6610 13280
rect 8662 13268 8668 13280
rect 8720 13308 8726 13320
rect 8757 13311 8815 13317
rect 8757 13308 8769 13311
rect 8720 13280 8769 13308
rect 8720 13268 8726 13280
rect 8757 13277 8769 13280
rect 8803 13277 8815 13311
rect 8757 13271 8815 13277
rect 9493 13311 9551 13317
rect 9493 13277 9505 13311
rect 9539 13277 9551 13311
rect 9493 13271 9551 13277
rect 2869 13243 2927 13249
rect 2869 13209 2881 13243
rect 2915 13240 2927 13243
rect 2961 13243 3019 13249
rect 2961 13240 2973 13243
rect 2915 13212 2973 13240
rect 2915 13209 2927 13212
rect 2869 13203 2927 13209
rect 2961 13209 2973 13212
rect 3007 13209 3019 13243
rect 2961 13203 3019 13209
rect 4893 13243 4951 13249
rect 4893 13209 4905 13243
rect 4939 13240 4951 13243
rect 4985 13243 5043 13249
rect 4985 13240 4997 13243
rect 4939 13212 4997 13240
rect 4939 13209 4951 13212
rect 4893 13203 4951 13209
rect 4985 13209 4997 13212
rect 5031 13209 5043 13243
rect 4985 13203 5043 13209
rect 5353 13243 5411 13249
rect 5353 13209 5365 13243
rect 5399 13209 5411 13243
rect 9508 13240 9536 13271
rect 9674 13268 9680 13320
rect 9732 13308 9738 13320
rect 12434 13317 12440 13320
rect 10873 13311 10931 13317
rect 9732 13280 9777 13308
rect 9732 13268 9738 13280
rect 10873 13277 10885 13311
rect 10919 13277 10931 13311
rect 12391 13311 12440 13317
rect 12391 13308 12403 13311
rect 12347 13280 12403 13308
rect 10873 13271 10931 13277
rect 12391 13277 12403 13280
rect 12437 13277 12440 13311
rect 12391 13271 12440 13277
rect 10778 13240 10784 13252
rect 9508 13212 10784 13240
rect 5353 13203 5411 13209
rect 10778 13200 10784 13212
rect 10836 13240 10842 13252
rect 10888 13240 10916 13271
rect 12406 13268 12440 13271
rect 12492 13308 12498 13320
rect 15102 13308 15108 13320
rect 12492 13280 15108 13308
rect 12492 13268 12498 13280
rect 15102 13268 15108 13280
rect 15160 13268 15166 13320
rect 12406 13240 12434 13268
rect 10836 13212 12434 13240
rect 10836 13200 10842 13212
rect 3234 13132 3240 13184
rect 3292 13172 3298 13184
rect 3329 13175 3387 13181
rect 3329 13172 3341 13175
rect 3292 13144 3341 13172
rect 3292 13132 3298 13144
rect 3329 13141 3341 13144
rect 3375 13141 3387 13175
rect 3329 13135 3387 13141
rect 4430 13132 4436 13184
rect 4488 13172 4494 13184
rect 8205 13175 8263 13181
rect 8205 13172 8217 13175
rect 4488 13144 8217 13172
rect 4488 13132 4494 13144
rect 8205 13141 8217 13144
rect 8251 13141 8263 13175
rect 10134 13172 10140 13184
rect 10095 13144 10140 13172
rect 8205 13135 8263 13141
rect 10134 13132 10140 13144
rect 10192 13132 10198 13184
rect 1104 13082 16836 13104
rect 1104 13030 3604 13082
rect 3656 13030 3668 13082
rect 3720 13030 3732 13082
rect 3784 13030 3796 13082
rect 3848 13030 8848 13082
rect 8900 13030 8912 13082
rect 8964 13030 8976 13082
rect 9028 13030 9040 13082
rect 9092 13030 14092 13082
rect 14144 13030 14156 13082
rect 14208 13030 14220 13082
rect 14272 13030 14284 13082
rect 14336 13030 16836 13082
rect 1104 13008 16836 13030
rect 6454 12968 6460 12980
rect 6415 12940 6460 12968
rect 6454 12928 6460 12940
rect 6512 12928 6518 12980
rect 6546 12928 6552 12980
rect 6604 12968 6610 12980
rect 6822 12968 6828 12980
rect 6604 12940 6828 12968
rect 6604 12928 6610 12940
rect 6822 12928 6828 12940
rect 6880 12968 6886 12980
rect 7101 12971 7159 12977
rect 7101 12968 7113 12971
rect 6880 12940 7113 12968
rect 6880 12928 6886 12940
rect 7101 12937 7113 12940
rect 7147 12937 7159 12971
rect 7101 12931 7159 12937
rect 7190 12928 7196 12980
rect 7248 12968 7254 12980
rect 7285 12971 7343 12977
rect 7285 12968 7297 12971
rect 7248 12940 7297 12968
rect 7248 12928 7254 12940
rect 7285 12937 7297 12940
rect 7331 12937 7343 12971
rect 7558 12968 7564 12980
rect 7519 12940 7564 12968
rect 7285 12931 7343 12937
rect 4798 12900 4804 12912
rect 4759 12872 4804 12900
rect 4798 12860 4804 12872
rect 4856 12860 4862 12912
rect 7300 12900 7328 12931
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 8570 12928 8576 12980
rect 8628 12968 8634 12980
rect 11241 12971 11299 12977
rect 11241 12968 11253 12971
rect 8628 12940 11253 12968
rect 8628 12928 8634 12940
rect 11241 12937 11253 12940
rect 11287 12937 11299 12971
rect 11241 12931 11299 12937
rect 11701 12971 11759 12977
rect 11701 12937 11713 12971
rect 11747 12968 11759 12971
rect 11790 12968 11796 12980
rect 11747 12940 11796 12968
rect 11747 12937 11759 12940
rect 11701 12931 11759 12937
rect 8478 12900 8484 12912
rect 7300 12872 8484 12900
rect 8478 12860 8484 12872
rect 8536 12860 8542 12912
rect 11256 12900 11284 12931
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 13906 12928 13912 12980
rect 13964 12968 13970 12980
rect 14001 12971 14059 12977
rect 14001 12968 14013 12971
rect 13964 12940 14013 12968
rect 13964 12928 13970 12940
rect 14001 12937 14013 12940
rect 14047 12937 14059 12971
rect 15378 12968 15384 12980
rect 15339 12940 15384 12968
rect 14001 12931 14059 12937
rect 12158 12900 12164 12912
rect 11256 12872 12164 12900
rect 12158 12860 12164 12872
rect 12216 12860 12222 12912
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12832 2375 12835
rect 2774 12832 2780 12844
rect 2363 12804 2780 12832
rect 2363 12801 2375 12804
rect 2317 12795 2375 12801
rect 2774 12792 2780 12804
rect 2832 12832 2838 12844
rect 3142 12832 3148 12844
rect 2832 12804 3148 12832
rect 2832 12792 2838 12804
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 4430 12832 4436 12844
rect 4356 12804 4436 12832
rect 3234 12764 3240 12776
rect 3195 12736 3240 12764
rect 3234 12724 3240 12736
rect 3292 12724 3298 12776
rect 3605 12767 3663 12773
rect 3605 12733 3617 12767
rect 3651 12764 3663 12767
rect 3789 12767 3847 12773
rect 3789 12764 3801 12767
rect 3651 12736 3801 12764
rect 3651 12733 3663 12736
rect 3605 12727 3663 12733
rect 3789 12733 3801 12736
rect 3835 12764 3847 12767
rect 3970 12764 3976 12776
rect 3835 12736 3976 12764
rect 3835 12733 3847 12736
rect 3789 12727 3847 12733
rect 3970 12724 3976 12736
rect 4028 12724 4034 12776
rect 4356 12773 4384 12804
rect 4430 12792 4436 12804
rect 4488 12792 4494 12844
rect 5902 12792 5908 12844
rect 5960 12832 5966 12844
rect 6638 12832 6644 12844
rect 5960 12804 6644 12832
rect 5960 12792 5966 12804
rect 6638 12792 6644 12804
rect 6696 12792 6702 12844
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12832 6883 12835
rect 7098 12832 7104 12844
rect 6871 12804 7104 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 7098 12792 7104 12804
rect 7156 12792 7162 12844
rect 8113 12835 8171 12841
rect 8113 12801 8125 12835
rect 8159 12832 8171 12835
rect 8662 12832 8668 12844
rect 8159 12804 8668 12832
rect 8159 12801 8171 12804
rect 8113 12795 8171 12801
rect 8662 12792 8668 12804
rect 8720 12832 8726 12844
rect 9953 12835 10011 12841
rect 9953 12832 9965 12835
rect 8720 12804 9965 12832
rect 8720 12792 8726 12804
rect 9953 12801 9965 12804
rect 9999 12801 10011 12835
rect 9953 12795 10011 12801
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 10192 12804 11284 12832
rect 10192 12792 10198 12804
rect 4341 12767 4399 12773
rect 4341 12733 4353 12767
rect 4387 12733 4399 12767
rect 4341 12727 4399 12733
rect 6730 12724 6736 12776
rect 6788 12764 6794 12776
rect 6914 12764 6920 12776
rect 6788 12736 6833 12764
rect 6875 12736 6920 12764
rect 6788 12724 6794 12736
rect 6914 12724 6920 12736
rect 6972 12724 6978 12776
rect 7116 12764 7144 12792
rect 8202 12764 8208 12776
rect 7116 12736 8208 12764
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 10778 12764 10784 12776
rect 10739 12736 10784 12764
rect 10778 12724 10784 12736
rect 10836 12724 10842 12776
rect 10870 12724 10876 12776
rect 10928 12764 10934 12776
rect 11256 12764 11284 12804
rect 11330 12792 11336 12844
rect 11388 12832 11394 12844
rect 12345 12835 12403 12841
rect 12345 12832 12357 12835
rect 11388 12804 12357 12832
rect 11388 12792 11394 12804
rect 12345 12801 12357 12804
rect 12391 12832 12403 12835
rect 12802 12832 12808 12844
rect 12391 12804 12808 12832
rect 12391 12801 12403 12804
rect 12345 12795 12403 12801
rect 12802 12792 12808 12804
rect 12860 12792 12866 12844
rect 14016 12832 14044 12931
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 14461 12903 14519 12909
rect 14461 12869 14473 12903
rect 14507 12900 14519 12903
rect 14553 12903 14611 12909
rect 14553 12900 14565 12903
rect 14507 12872 14565 12900
rect 14507 12869 14519 12872
rect 14461 12863 14519 12869
rect 14553 12869 14565 12872
rect 14599 12869 14611 12903
rect 14553 12863 14611 12869
rect 14016 12804 14228 12832
rect 13449 12767 13507 12773
rect 13449 12764 13461 12767
rect 10928 12736 11192 12764
rect 11256 12736 13461 12764
rect 10928 12724 10934 12736
rect 2222 12656 2228 12708
rect 2280 12696 2286 12708
rect 2961 12699 3019 12705
rect 2961 12696 2973 12699
rect 2280 12668 2973 12696
rect 2280 12656 2286 12668
rect 2961 12665 2973 12668
rect 3007 12696 3019 12699
rect 3421 12699 3479 12705
rect 3421 12696 3433 12699
rect 3007 12668 3433 12696
rect 3007 12665 3019 12668
rect 2961 12659 3019 12665
rect 3421 12665 3433 12668
rect 3467 12665 3479 12699
rect 3421 12659 3479 12665
rect 3881 12699 3939 12705
rect 3881 12665 3893 12699
rect 3927 12696 3939 12699
rect 3927 12668 4844 12696
rect 3927 12665 3939 12668
rect 3881 12659 3939 12665
rect 4816 12637 4844 12668
rect 6086 12656 6092 12708
rect 6144 12696 6150 12708
rect 7253 12699 7311 12705
rect 7253 12696 7265 12699
rect 6144 12668 7265 12696
rect 6144 12656 6150 12668
rect 7253 12665 7265 12668
rect 7299 12696 7311 12699
rect 7374 12696 7380 12708
rect 7299 12668 7380 12696
rect 7299 12665 7311 12668
rect 7253 12659 7311 12665
rect 7374 12656 7380 12668
rect 7432 12656 7438 12708
rect 7469 12699 7527 12705
rect 7469 12665 7481 12699
rect 7515 12665 7527 12699
rect 7469 12659 7527 12665
rect 7929 12699 7987 12705
rect 7929 12665 7941 12699
rect 7975 12696 7987 12699
rect 8294 12696 8300 12708
rect 7975 12668 8300 12696
rect 7975 12665 7987 12668
rect 7929 12659 7987 12665
rect 4801 12631 4859 12637
rect 4801 12597 4813 12631
rect 4847 12628 4859 12631
rect 4982 12628 4988 12640
rect 4847 12600 4988 12628
rect 4847 12597 4859 12600
rect 4801 12591 4859 12597
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 6914 12588 6920 12640
rect 6972 12628 6978 12640
rect 7484 12628 7512 12659
rect 8294 12656 8300 12668
rect 8352 12656 8358 12708
rect 11057 12699 11115 12705
rect 11057 12665 11069 12699
rect 11103 12665 11115 12699
rect 11164 12696 11192 12736
rect 13449 12733 13461 12736
rect 13495 12733 13507 12767
rect 13998 12764 14004 12776
rect 13959 12736 14004 12764
rect 13449 12727 13507 12733
rect 11330 12696 11336 12708
rect 11164 12668 11336 12696
rect 11057 12659 11115 12665
rect 7834 12628 7840 12640
rect 6972 12600 7840 12628
rect 6972 12588 6978 12600
rect 7834 12588 7840 12600
rect 7892 12588 7898 12640
rect 8018 12588 8024 12640
rect 8076 12628 8082 12640
rect 8076 12600 8121 12628
rect 8076 12588 8082 12600
rect 10318 12588 10324 12640
rect 10376 12628 10382 12640
rect 11072 12628 11100 12659
rect 11330 12656 11336 12668
rect 11388 12696 11394 12708
rect 12161 12699 12219 12705
rect 12161 12696 12173 12699
rect 11388 12668 12173 12696
rect 11388 12656 11394 12668
rect 12161 12665 12173 12668
rect 12207 12665 12219 12699
rect 13464 12696 13492 12727
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 14093 12767 14151 12773
rect 14093 12733 14105 12767
rect 14139 12733 14151 12767
rect 14093 12727 14151 12733
rect 14108 12696 14136 12727
rect 13464 12668 14136 12696
rect 12161 12659 12219 12665
rect 11238 12628 11244 12640
rect 10376 12600 11244 12628
rect 10376 12588 10382 12600
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 12069 12631 12127 12637
rect 12069 12628 12081 12631
rect 11848 12600 12081 12628
rect 11848 12588 11854 12600
rect 12069 12597 12081 12600
rect 12115 12597 12127 12631
rect 14200 12628 14228 12804
rect 15102 12792 15108 12844
rect 15160 12832 15166 12844
rect 15933 12835 15991 12841
rect 15933 12832 15945 12835
rect 15160 12804 15945 12832
rect 15160 12792 15166 12804
rect 15933 12801 15945 12804
rect 15979 12801 15991 12835
rect 15933 12795 15991 12801
rect 14274 12724 14280 12776
rect 14332 12764 14338 12776
rect 14737 12767 14795 12773
rect 14737 12764 14749 12767
rect 14332 12736 14749 12764
rect 14332 12724 14338 12736
rect 14737 12733 14749 12736
rect 14783 12764 14795 12767
rect 14826 12764 14832 12776
rect 14783 12736 14832 12764
rect 14783 12733 14795 12736
rect 14737 12727 14795 12733
rect 14826 12724 14832 12736
rect 14884 12724 14890 12776
rect 15841 12767 15899 12773
rect 15841 12733 15853 12767
rect 15887 12764 15899 12767
rect 16298 12764 16304 12776
rect 15887 12736 16304 12764
rect 15887 12733 15899 12736
rect 15841 12727 15899 12733
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 14461 12631 14519 12637
rect 14461 12628 14473 12631
rect 14200 12600 14473 12628
rect 12069 12591 12127 12597
rect 14461 12597 14473 12600
rect 14507 12597 14519 12631
rect 15746 12628 15752 12640
rect 15707 12600 15752 12628
rect 14461 12591 14519 12597
rect 15746 12588 15752 12600
rect 15804 12588 15810 12640
rect 1104 12538 16836 12560
rect 1104 12486 6226 12538
rect 6278 12486 6290 12538
rect 6342 12486 6354 12538
rect 6406 12486 6418 12538
rect 6470 12486 11470 12538
rect 11522 12486 11534 12538
rect 11586 12486 11598 12538
rect 11650 12486 11662 12538
rect 11714 12486 16836 12538
rect 1104 12464 16836 12486
rect 7101 12427 7159 12433
rect 7101 12393 7113 12427
rect 7147 12424 7159 12427
rect 7190 12424 7196 12436
rect 7147 12396 7196 12424
rect 7147 12393 7159 12396
rect 7101 12387 7159 12393
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 9858 12384 9864 12436
rect 9916 12424 9922 12436
rect 10594 12424 10600 12436
rect 9916 12396 9961 12424
rect 10555 12396 10600 12424
rect 9916 12384 9922 12396
rect 10594 12384 10600 12396
rect 10652 12384 10658 12436
rect 11330 12424 11336 12436
rect 11256 12396 11336 12424
rect 1857 12359 1915 12365
rect 1857 12325 1869 12359
rect 1903 12356 1915 12359
rect 2130 12356 2136 12368
rect 1903 12328 2136 12356
rect 1903 12325 1915 12328
rect 1857 12319 1915 12325
rect 2130 12316 2136 12328
rect 2188 12316 2194 12368
rect 7852 12328 8156 12356
rect 7852 12300 7880 12328
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 2041 12291 2099 12297
rect 2041 12257 2053 12291
rect 2087 12288 2099 12291
rect 2774 12288 2780 12300
rect 2087 12260 2780 12288
rect 2087 12257 2099 12260
rect 2041 12251 2099 12257
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 5350 12248 5356 12300
rect 5408 12288 5414 12300
rect 6365 12291 6423 12297
rect 6365 12288 6377 12291
rect 5408 12260 6377 12288
rect 5408 12248 5414 12260
rect 6365 12257 6377 12260
rect 6411 12257 6423 12291
rect 6365 12251 6423 12257
rect 6730 12248 6736 12300
rect 6788 12288 6794 12300
rect 6825 12291 6883 12297
rect 6825 12288 6837 12291
rect 6788 12260 6837 12288
rect 6788 12248 6794 12260
rect 6825 12257 6837 12260
rect 6871 12257 6883 12291
rect 6825 12251 6883 12257
rect 7009 12291 7067 12297
rect 7009 12257 7021 12291
rect 7055 12288 7067 12291
rect 7098 12288 7104 12300
rect 7055 12260 7104 12288
rect 7055 12257 7067 12260
rect 7009 12251 7067 12257
rect 7098 12248 7104 12260
rect 7156 12248 7162 12300
rect 7561 12291 7619 12297
rect 7561 12257 7573 12291
rect 7607 12257 7619 12291
rect 7834 12288 7840 12300
rect 7795 12260 7840 12288
rect 7561 12251 7619 12257
rect 6089 12223 6147 12229
rect 6089 12189 6101 12223
rect 6135 12220 6147 12223
rect 6914 12220 6920 12232
rect 6135 12192 6920 12220
rect 6135 12189 6147 12192
rect 6089 12183 6147 12189
rect 6914 12180 6920 12192
rect 6972 12180 6978 12232
rect 7190 12180 7196 12232
rect 7248 12220 7254 12232
rect 7576 12220 7604 12251
rect 7834 12248 7840 12260
rect 7892 12248 7898 12300
rect 8021 12291 8079 12297
rect 8021 12257 8033 12291
rect 8067 12257 8079 12291
rect 8128 12288 8156 12328
rect 8478 12316 8484 12368
rect 8536 12356 8542 12368
rect 10226 12356 10232 12368
rect 8536 12328 10232 12356
rect 8536 12316 8542 12328
rect 10226 12316 10232 12328
rect 10284 12316 10290 12368
rect 10870 12356 10876 12368
rect 10520 12328 10876 12356
rect 8128 12260 9996 12288
rect 8021 12251 8079 12257
rect 7248 12192 7604 12220
rect 7248 12180 7254 12192
rect 1578 12152 1584 12164
rect 1539 12124 1584 12152
rect 1578 12112 1584 12124
rect 1636 12112 1642 12164
rect 6549 12155 6607 12161
rect 6549 12152 6561 12155
rect 6104 12124 6561 12152
rect 6104 12096 6132 12124
rect 6549 12121 6561 12124
rect 6595 12152 6607 12155
rect 8036 12152 8064 12251
rect 8294 12220 8300 12232
rect 8255 12192 8300 12220
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 8386 12180 8392 12232
rect 8444 12220 8450 12232
rect 9674 12220 9680 12232
rect 8444 12192 9680 12220
rect 8444 12180 8450 12192
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 9968 12220 9996 12260
rect 10042 12248 10048 12300
rect 10100 12288 10106 12300
rect 10318 12288 10324 12300
rect 10100 12260 10145 12288
rect 10279 12260 10324 12288
rect 10100 12248 10106 12260
rect 10318 12248 10324 12260
rect 10376 12248 10382 12300
rect 10520 12297 10548 12328
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 10505 12291 10563 12297
rect 10505 12257 10517 12291
rect 10551 12257 10563 12291
rect 10778 12288 10784 12300
rect 10739 12260 10784 12288
rect 10505 12251 10563 12257
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 11146 12297 11152 12300
rect 11102 12291 11152 12297
rect 11102 12257 11114 12291
rect 11148 12257 11152 12291
rect 11102 12251 11152 12257
rect 11146 12248 11152 12251
rect 11204 12248 11210 12300
rect 11256 12297 11284 12396
rect 11330 12384 11336 12396
rect 11388 12384 11394 12436
rect 11974 12424 11980 12436
rect 11935 12396 11980 12424
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 12066 12384 12072 12436
rect 12124 12424 12130 12436
rect 12342 12424 12348 12436
rect 12124 12396 12348 12424
rect 12124 12384 12130 12396
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 15473 12427 15531 12433
rect 15473 12393 15485 12427
rect 15519 12424 15531 12427
rect 15746 12424 15752 12436
rect 15519 12396 15752 12424
rect 15519 12393 15531 12396
rect 15473 12387 15531 12393
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 11701 12359 11759 12365
rect 11701 12356 11713 12359
rect 11348 12328 11713 12356
rect 11241 12291 11299 12297
rect 11241 12257 11253 12291
rect 11287 12257 11299 12291
rect 11241 12251 11299 12257
rect 10336 12220 10364 12248
rect 10870 12220 10876 12232
rect 9968 12192 10364 12220
rect 10831 12192 10876 12220
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 11348 12220 11376 12328
rect 11701 12325 11713 12328
rect 11747 12356 11759 12359
rect 12989 12359 13047 12365
rect 12989 12356 13001 12359
rect 11747 12328 13001 12356
rect 11747 12325 11759 12328
rect 11701 12319 11759 12325
rect 12989 12325 13001 12328
rect 13035 12356 13047 12359
rect 13170 12356 13176 12368
rect 13035 12328 13176 12356
rect 13035 12325 13047 12328
rect 12989 12319 13047 12325
rect 13170 12316 13176 12328
rect 13228 12316 13234 12368
rect 14826 12316 14832 12368
rect 14884 12356 14890 12368
rect 14884 12328 15976 12356
rect 14884 12316 14890 12328
rect 11517 12291 11575 12297
rect 11517 12257 11529 12291
rect 11563 12257 11575 12291
rect 11790 12288 11796 12300
rect 11751 12260 11796 12288
rect 11517 12251 11575 12257
rect 10980 12192 11376 12220
rect 11532 12220 11560 12251
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 11974 12288 11980 12300
rect 11935 12260 11980 12288
rect 11974 12248 11980 12260
rect 12032 12248 12038 12300
rect 12066 12248 12072 12300
rect 12124 12288 12130 12300
rect 12437 12291 12495 12297
rect 12437 12288 12449 12291
rect 12124 12260 12449 12288
rect 12124 12248 12130 12260
rect 12437 12257 12449 12260
rect 12483 12257 12495 12291
rect 12802 12288 12808 12300
rect 12763 12260 12808 12288
rect 12437 12251 12495 12257
rect 12802 12248 12808 12260
rect 12860 12248 12866 12300
rect 15562 12248 15568 12300
rect 15620 12288 15626 12300
rect 15948 12297 15976 12328
rect 15749 12291 15807 12297
rect 15749 12288 15761 12291
rect 15620 12260 15761 12288
rect 15620 12248 15626 12260
rect 15749 12257 15761 12260
rect 15795 12257 15807 12291
rect 15749 12251 15807 12257
rect 15933 12291 15991 12297
rect 15933 12257 15945 12291
rect 15979 12257 15991 12291
rect 15933 12251 15991 12257
rect 13262 12220 13268 12232
rect 11532 12192 13268 12220
rect 9398 12152 9404 12164
rect 6595 12124 9404 12152
rect 6595 12121 6607 12124
rect 6549 12115 6607 12121
rect 9398 12112 9404 12124
rect 9456 12112 9462 12164
rect 9490 12112 9496 12164
rect 9548 12152 9554 12164
rect 10137 12155 10195 12161
rect 10137 12152 10149 12155
rect 9548 12124 10149 12152
rect 9548 12112 9554 12124
rect 10137 12121 10149 12124
rect 10183 12121 10195 12155
rect 10137 12115 10195 12121
rect 10226 12112 10232 12164
rect 10284 12152 10290 12164
rect 10980 12161 11008 12192
rect 10965 12155 11023 12161
rect 10965 12152 10977 12155
rect 10284 12124 10977 12152
rect 10284 12112 10290 12124
rect 10965 12121 10977 12124
rect 11011 12121 11023 12155
rect 10965 12115 11023 12121
rect 11146 12112 11152 12164
rect 11204 12152 11210 12164
rect 11532 12152 11560 12192
rect 13262 12180 13268 12192
rect 13320 12220 13326 12232
rect 15657 12223 15715 12229
rect 15657 12220 15669 12223
rect 13320 12192 15669 12220
rect 13320 12180 13326 12192
rect 15657 12189 15669 12192
rect 15703 12189 15715 12223
rect 15841 12223 15899 12229
rect 15841 12220 15853 12223
rect 15657 12183 15715 12189
rect 15764 12192 15853 12220
rect 11204 12124 11560 12152
rect 11204 12112 11210 12124
rect 11974 12112 11980 12164
rect 12032 12152 12038 12164
rect 14550 12152 14556 12164
rect 12032 12124 14556 12152
rect 12032 12112 12038 12124
rect 14550 12112 14556 12124
rect 14608 12112 14614 12164
rect 1762 12084 1768 12096
rect 1723 12056 1768 12084
rect 1762 12044 1768 12056
rect 1820 12044 1826 12096
rect 6086 12044 6092 12096
rect 6144 12044 6150 12096
rect 6178 12044 6184 12096
rect 6236 12084 6242 12096
rect 6236 12056 6281 12084
rect 6236 12044 6242 12056
rect 7650 12044 7656 12096
rect 7708 12084 7714 12096
rect 7745 12087 7803 12093
rect 7745 12084 7757 12087
rect 7708 12056 7757 12084
rect 7708 12044 7714 12056
rect 7745 12053 7757 12056
rect 7791 12053 7803 12087
rect 7926 12084 7932 12096
rect 7887 12056 7932 12084
rect 7745 12047 7803 12053
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 12342 12084 12348 12096
rect 8260 12056 12348 12084
rect 8260 12044 8266 12056
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 13814 12044 13820 12096
rect 13872 12084 13878 12096
rect 15764 12084 15792 12192
rect 15841 12189 15853 12192
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 13872 12056 15792 12084
rect 13872 12044 13878 12056
rect 1104 11994 16836 12016
rect 1104 11942 3604 11994
rect 3656 11942 3668 11994
rect 3720 11942 3732 11994
rect 3784 11942 3796 11994
rect 3848 11942 8848 11994
rect 8900 11942 8912 11994
rect 8964 11942 8976 11994
rect 9028 11942 9040 11994
rect 9092 11942 14092 11994
rect 14144 11942 14156 11994
rect 14208 11942 14220 11994
rect 14272 11942 14284 11994
rect 14336 11942 16836 11994
rect 1104 11920 16836 11942
rect 7926 11880 7932 11892
rect 6656 11852 7932 11880
rect 6656 11824 6684 11852
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 9677 11883 9735 11889
rect 8956 11852 9260 11880
rect 8956 11824 8984 11852
rect 6638 11812 6644 11824
rect 6599 11784 6644 11812
rect 6638 11772 6644 11784
rect 6696 11772 6702 11824
rect 7009 11815 7067 11821
rect 7009 11781 7021 11815
rect 7055 11812 7067 11815
rect 8846 11812 8852 11824
rect 7055 11784 8852 11812
rect 7055 11781 7067 11784
rect 7009 11775 7067 11781
rect 8846 11772 8852 11784
rect 8904 11772 8910 11824
rect 8938 11772 8944 11824
rect 8996 11772 9002 11824
rect 9232 11821 9260 11852
rect 9677 11849 9689 11883
rect 9723 11880 9735 11883
rect 9766 11880 9772 11892
rect 9723 11852 9772 11880
rect 9723 11849 9735 11852
rect 9677 11843 9735 11849
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 10045 11883 10103 11889
rect 10045 11849 10057 11883
rect 10091 11880 10103 11883
rect 10134 11880 10140 11892
rect 10091 11852 10140 11880
rect 10091 11849 10103 11852
rect 10045 11843 10103 11849
rect 10134 11840 10140 11852
rect 10192 11880 10198 11892
rect 12250 11880 12256 11892
rect 10192 11852 12256 11880
rect 10192 11840 10198 11852
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 12621 11883 12679 11889
rect 12621 11849 12633 11883
rect 12667 11880 12679 11883
rect 12894 11880 12900 11892
rect 12667 11852 12900 11880
rect 12667 11849 12679 11852
rect 12621 11843 12679 11849
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 12989 11883 13047 11889
rect 12989 11849 13001 11883
rect 13035 11880 13047 11883
rect 13262 11880 13268 11892
rect 13035 11852 13268 11880
rect 13035 11849 13047 11852
rect 12989 11843 13047 11849
rect 9217 11815 9275 11821
rect 9217 11781 9229 11815
rect 9263 11781 9275 11815
rect 9858 11812 9864 11824
rect 9217 11775 9275 11781
rect 9600 11784 9864 11812
rect 8570 11704 8576 11756
rect 8628 11744 8634 11756
rect 9125 11747 9183 11753
rect 9125 11744 9137 11747
rect 8628 11716 9137 11744
rect 8628 11704 8634 11716
rect 9125 11713 9137 11716
rect 9171 11713 9183 11747
rect 9125 11707 9183 11713
rect 1581 11679 1639 11685
rect 1581 11645 1593 11679
rect 1627 11676 1639 11679
rect 1762 11676 1768 11688
rect 1627 11648 1768 11676
rect 1627 11645 1639 11648
rect 1581 11639 1639 11645
rect 1762 11636 1768 11648
rect 1820 11636 1826 11688
rect 2406 11636 2412 11688
rect 2464 11676 2470 11688
rect 2501 11679 2559 11685
rect 2501 11676 2513 11679
rect 2464 11648 2513 11676
rect 2464 11636 2470 11648
rect 2501 11645 2513 11648
rect 2547 11645 2559 11679
rect 4982 11676 4988 11688
rect 4943 11648 4988 11676
rect 2501 11639 2559 11645
rect 4982 11636 4988 11648
rect 5040 11636 5046 11688
rect 6546 11676 6552 11688
rect 6507 11648 6552 11676
rect 6546 11636 6552 11648
rect 6604 11636 6610 11688
rect 6730 11676 6736 11688
rect 6691 11648 6736 11676
rect 6730 11636 6736 11648
rect 6788 11636 6794 11688
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 7190 11676 7196 11688
rect 6871 11648 7196 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 8478 11636 8484 11688
rect 8536 11676 8542 11688
rect 9033 11679 9091 11685
rect 9033 11676 9045 11679
rect 8536 11648 9045 11676
rect 8536 11636 8542 11648
rect 9033 11645 9045 11648
rect 9079 11645 9091 11679
rect 9033 11639 9091 11645
rect 9309 11679 9367 11685
rect 9309 11645 9321 11679
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 9493 11679 9551 11685
rect 9493 11645 9505 11679
rect 9539 11676 9551 11679
rect 9600 11676 9628 11784
rect 9858 11772 9864 11784
rect 9916 11772 9922 11824
rect 12434 11772 12440 11824
rect 12492 11812 12498 11824
rect 13004 11812 13032 11843
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 13722 11880 13728 11892
rect 13683 11852 13728 11880
rect 13722 11840 13728 11852
rect 13780 11840 13786 11892
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 15381 11883 15439 11889
rect 15381 11880 15393 11883
rect 15252 11852 15393 11880
rect 15252 11840 15258 11852
rect 15381 11849 15393 11852
rect 15427 11849 15439 11883
rect 15381 11843 15439 11849
rect 12492 11784 13032 11812
rect 12492 11772 12498 11784
rect 13078 11772 13084 11824
rect 13136 11812 13142 11824
rect 13173 11815 13231 11821
rect 13173 11812 13185 11815
rect 13136 11784 13185 11812
rect 13136 11772 13142 11784
rect 13173 11781 13185 11784
rect 13219 11781 13231 11815
rect 13173 11775 13231 11781
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11744 10011 11747
rect 11146 11744 11152 11756
rect 9999 11716 11152 11744
rect 9999 11713 10011 11716
rect 9953 11707 10011 11713
rect 11146 11704 11152 11716
rect 11204 11704 11210 11756
rect 11974 11744 11980 11756
rect 11256 11716 11980 11744
rect 9539 11648 9628 11676
rect 10045 11679 10103 11685
rect 9539 11645 9551 11648
rect 9493 11639 9551 11645
rect 10045 11645 10057 11679
rect 10091 11676 10103 11679
rect 10686 11676 10692 11688
rect 10091 11648 10692 11676
rect 10091 11645 10103 11648
rect 10045 11639 10103 11645
rect 2222 11608 2228 11620
rect 2183 11580 2228 11608
rect 2222 11568 2228 11580
rect 2280 11568 2286 11620
rect 6748 11608 6776 11636
rect 7650 11608 7656 11620
rect 6748 11580 7656 11608
rect 7650 11568 7656 11580
rect 7708 11568 7714 11620
rect 9324 11608 9352 11639
rect 10686 11636 10692 11648
rect 10744 11676 10750 11688
rect 11256 11676 11284 11716
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11744 12219 11747
rect 12802 11744 12808 11756
rect 12207 11716 12808 11744
rect 12207 11713 12219 11716
rect 12161 11707 12219 11713
rect 12802 11704 12808 11716
rect 12860 11744 12866 11756
rect 14185 11747 14243 11753
rect 12860 11716 13492 11744
rect 12860 11704 12866 11716
rect 12066 11676 12072 11688
rect 10744 11648 11284 11676
rect 12027 11648 12072 11676
rect 10744 11636 10750 11648
rect 12066 11636 12072 11648
rect 12124 11636 12130 11688
rect 12250 11676 12256 11688
rect 12211 11648 12256 11676
rect 12250 11636 12256 11648
rect 12308 11636 12314 11688
rect 12345 11679 12403 11685
rect 12345 11645 12357 11679
rect 12391 11676 12403 11679
rect 12434 11676 12440 11688
rect 12391 11648 12440 11676
rect 12391 11645 12403 11648
rect 12345 11639 12403 11645
rect 12434 11636 12440 11648
rect 12492 11636 12498 11688
rect 12710 11636 12716 11688
rect 12768 11676 12774 11688
rect 13096 11685 13124 11716
rect 12897 11679 12955 11685
rect 12897 11676 12909 11679
rect 12768 11648 12909 11676
rect 12768 11636 12774 11648
rect 12897 11645 12909 11648
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 13081 11679 13139 11685
rect 13081 11645 13093 11679
rect 13127 11645 13139 11679
rect 13081 11639 13139 11645
rect 13262 11636 13268 11688
rect 13320 11676 13326 11688
rect 13357 11679 13415 11685
rect 13357 11676 13369 11679
rect 13320 11648 13369 11676
rect 13320 11636 13326 11648
rect 13357 11645 13369 11648
rect 13403 11645 13415 11679
rect 13464 11676 13492 11716
rect 14185 11713 14197 11747
rect 14231 11744 14243 11747
rect 14274 11744 14280 11756
rect 14231 11716 14280 11744
rect 14231 11713 14243 11716
rect 14185 11707 14243 11713
rect 14274 11704 14280 11716
rect 14332 11704 14338 11756
rect 14369 11747 14427 11753
rect 14369 11713 14381 11747
rect 14415 11744 14427 11747
rect 15102 11744 15108 11756
rect 14415 11716 15108 11744
rect 14415 11713 14427 11716
rect 14369 11707 14427 11713
rect 15102 11704 15108 11716
rect 15160 11744 15166 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15160 11716 15945 11744
rect 15160 11704 15166 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 14826 11676 14832 11688
rect 13464 11648 14832 11676
rect 13357 11639 13415 11645
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 15746 11676 15752 11688
rect 15707 11648 15752 11676
rect 15746 11636 15752 11648
rect 15804 11636 15810 11688
rect 9674 11608 9680 11620
rect 9324 11580 9680 11608
rect 9674 11568 9680 11580
rect 9732 11568 9738 11620
rect 14550 11608 14556 11620
rect 14511 11580 14556 11608
rect 14550 11568 14556 11580
rect 14608 11568 14614 11620
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 5077 11543 5135 11549
rect 5077 11540 5089 11543
rect 4396 11512 5089 11540
rect 4396 11500 4402 11512
rect 5077 11509 5089 11512
rect 5123 11509 5135 11543
rect 5077 11503 5135 11509
rect 8849 11543 8907 11549
rect 8849 11509 8861 11543
rect 8895 11540 8907 11543
rect 9214 11540 9220 11552
rect 8895 11512 9220 11540
rect 8895 11509 8907 11512
rect 8849 11503 8907 11509
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 12529 11543 12587 11549
rect 12529 11509 12541 11543
rect 12575 11540 12587 11543
rect 13998 11540 14004 11552
rect 12575 11512 14004 11540
rect 12575 11509 12587 11512
rect 12529 11503 12587 11509
rect 13998 11500 14004 11512
rect 14056 11540 14062 11552
rect 14090 11540 14096 11552
rect 14056 11512 14096 11540
rect 14056 11500 14062 11512
rect 14090 11500 14096 11512
rect 14148 11500 14154 11552
rect 14274 11500 14280 11552
rect 14332 11540 14338 11552
rect 15746 11540 15752 11552
rect 14332 11512 15752 11540
rect 14332 11500 14338 11512
rect 15746 11500 15752 11512
rect 15804 11500 15810 11552
rect 15841 11543 15899 11549
rect 15841 11509 15853 11543
rect 15887 11540 15899 11543
rect 16022 11540 16028 11552
rect 15887 11512 16028 11540
rect 15887 11509 15899 11512
rect 15841 11503 15899 11509
rect 16022 11500 16028 11512
rect 16080 11500 16086 11552
rect 1104 11450 16836 11472
rect 1104 11398 6226 11450
rect 6278 11398 6290 11450
rect 6342 11398 6354 11450
rect 6406 11398 6418 11450
rect 6470 11398 11470 11450
rect 11522 11398 11534 11450
rect 11586 11398 11598 11450
rect 11650 11398 11662 11450
rect 11714 11398 16836 11450
rect 1104 11376 16836 11398
rect 5074 11336 5080 11348
rect 4632 11308 5080 11336
rect 2961 11271 3019 11277
rect 2961 11237 2973 11271
rect 3007 11268 3019 11271
rect 3326 11268 3332 11280
rect 3007 11240 3332 11268
rect 3007 11237 3019 11240
rect 2961 11231 3019 11237
rect 3326 11228 3332 11240
rect 3384 11228 3390 11280
rect 4632 11277 4660 11308
rect 5074 11296 5080 11308
rect 5132 11336 5138 11348
rect 5537 11339 5595 11345
rect 5537 11336 5549 11339
rect 5132 11308 5549 11336
rect 5132 11296 5138 11308
rect 5537 11305 5549 11308
rect 5583 11305 5595 11339
rect 5537 11299 5595 11305
rect 7834 11296 7840 11348
rect 7892 11336 7898 11348
rect 7892 11308 9168 11336
rect 7892 11296 7898 11308
rect 4617 11271 4675 11277
rect 4617 11237 4629 11271
rect 4663 11237 4675 11271
rect 9030 11268 9036 11280
rect 4617 11231 4675 11237
rect 5000 11240 5856 11268
rect 1578 11200 1584 11212
rect 1539 11172 1584 11200
rect 1578 11160 1584 11172
rect 1636 11160 1642 11212
rect 2317 11203 2375 11209
rect 2317 11169 2329 11203
rect 2363 11200 2375 11203
rect 2682 11200 2688 11212
rect 2363 11172 2688 11200
rect 2363 11169 2375 11172
rect 2317 11163 2375 11169
rect 2682 11160 2688 11172
rect 2740 11160 2746 11212
rect 4338 11160 4344 11212
rect 4396 11200 4402 11212
rect 4525 11203 4583 11209
rect 4525 11200 4537 11203
rect 4396 11172 4537 11200
rect 4396 11160 4402 11172
rect 4525 11169 4537 11172
rect 4571 11200 4583 11203
rect 5000 11200 5028 11240
rect 5828 11209 5856 11240
rect 8496 11240 9036 11268
rect 4571 11172 5028 11200
rect 5077 11203 5135 11209
rect 4571 11169 4583 11172
rect 4525 11163 4583 11169
rect 5077 11169 5089 11203
rect 5123 11169 5135 11203
rect 5077 11163 5135 11169
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11169 5871 11203
rect 7742 11200 7748 11212
rect 7703 11172 7748 11200
rect 5813 11163 5871 11169
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11101 2007 11135
rect 1949 11095 2007 11101
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 3142 11132 3148 11144
rect 3099 11104 3148 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 1964 11064 1992 11095
rect 2130 11064 2136 11076
rect 1964 11036 2136 11064
rect 2130 11024 2136 11036
rect 2188 11024 2194 11076
rect 2314 11024 2320 11076
rect 2372 11064 2378 11076
rect 2501 11067 2559 11073
rect 2501 11064 2513 11067
rect 2372 11036 2513 11064
rect 2372 11024 2378 11036
rect 2501 11033 2513 11036
rect 2547 11033 2559 11067
rect 2976 11064 3004 11095
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 5092 11132 5120 11163
rect 7742 11160 7748 11172
rect 7800 11160 7806 11212
rect 7837 11203 7895 11209
rect 7837 11169 7849 11203
rect 7883 11200 7895 11203
rect 8294 11200 8300 11212
rect 7883 11172 8300 11200
rect 7883 11169 7895 11172
rect 7837 11163 7895 11169
rect 8294 11160 8300 11172
rect 8352 11160 8358 11212
rect 8496 11209 8524 11240
rect 9030 11228 9036 11240
rect 9088 11228 9094 11280
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11169 8539 11203
rect 8481 11163 8539 11169
rect 8662 11160 8668 11212
rect 8720 11200 8726 11212
rect 8938 11200 8944 11212
rect 8720 11172 8944 11200
rect 8720 11160 8726 11172
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 9140 11200 9168 11308
rect 9214 11296 9220 11348
rect 9272 11336 9278 11348
rect 9272 11308 10456 11336
rect 9272 11296 9278 11308
rect 9582 11228 9588 11280
rect 9640 11268 9646 11280
rect 10321 11271 10379 11277
rect 10321 11268 10333 11271
rect 9640 11240 10333 11268
rect 9640 11228 9646 11240
rect 10321 11237 10333 11240
rect 10367 11237 10379 11271
rect 10428 11268 10456 11308
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 11241 11339 11299 11345
rect 11241 11336 11253 11339
rect 10928 11308 11253 11336
rect 10928 11296 10934 11308
rect 11241 11305 11253 11308
rect 11287 11305 11299 11339
rect 13354 11336 13360 11348
rect 11241 11299 11299 11305
rect 11348 11308 13360 11336
rect 11348 11268 11376 11308
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 16206 11296 16212 11348
rect 16264 11336 16270 11348
rect 16301 11339 16359 11345
rect 16301 11336 16313 11339
rect 16264 11308 16313 11336
rect 16264 11296 16270 11308
rect 16301 11305 16313 11308
rect 16347 11305 16359 11339
rect 16301 11299 16359 11305
rect 13262 11268 13268 11280
rect 10428 11240 11376 11268
rect 12268 11240 13268 11268
rect 10321 11231 10379 11237
rect 9674 11200 9680 11212
rect 9140 11172 9680 11200
rect 9674 11160 9680 11172
rect 9732 11200 9738 11212
rect 9950 11200 9956 11212
rect 9732 11172 9956 11200
rect 9732 11160 9738 11172
rect 9950 11160 9956 11172
rect 10008 11200 10014 11212
rect 10410 11200 10416 11212
rect 10008 11172 10416 11200
rect 10008 11160 10014 11172
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 10505 11203 10563 11209
rect 10505 11169 10517 11203
rect 10551 11169 10563 11203
rect 11146 11200 11152 11212
rect 11107 11172 11152 11200
rect 10505 11163 10563 11169
rect 5169 11135 5227 11141
rect 5169 11132 5181 11135
rect 5092 11104 5181 11132
rect 5169 11101 5181 11104
rect 5215 11132 5227 11135
rect 7926 11132 7932 11144
rect 5215 11104 7420 11132
rect 7887 11104 7932 11132
rect 5215 11101 5227 11104
rect 5169 11095 5227 11101
rect 7392 11073 7420 11104
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 8956 11132 8984 11160
rect 10045 11135 10103 11141
rect 10045 11132 10057 11135
rect 8956 11104 10057 11132
rect 10045 11101 10057 11104
rect 10091 11132 10103 11135
rect 10520 11132 10548 11163
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 11422 11160 11428 11212
rect 11480 11209 11486 11212
rect 11480 11200 11488 11209
rect 11480 11172 11525 11200
rect 11480 11163 11488 11172
rect 11480 11160 11486 11163
rect 11514 11132 11520 11144
rect 10091 11104 10548 11132
rect 11475 11104 11520 11132
rect 10091 11101 10103 11104
rect 10045 11095 10103 11101
rect 11514 11092 11520 11104
rect 11572 11132 11578 11144
rect 12268 11132 12296 11240
rect 13262 11228 13268 11240
rect 13320 11268 13326 11280
rect 14093 11271 14151 11277
rect 14093 11268 14105 11271
rect 13320 11240 14105 11268
rect 13320 11228 13326 11240
rect 14093 11237 14105 11240
rect 14139 11237 14151 11271
rect 14093 11231 14151 11237
rect 14461 11271 14519 11277
rect 14461 11237 14473 11271
rect 14507 11268 14519 11271
rect 15197 11271 15255 11277
rect 15197 11268 15209 11271
rect 14507 11240 15209 11268
rect 14507 11237 14519 11240
rect 14461 11231 14519 11237
rect 15197 11237 15209 11240
rect 15243 11237 15255 11271
rect 15197 11231 15255 11237
rect 15381 11271 15439 11277
rect 15381 11237 15393 11271
rect 15427 11268 15439 11271
rect 15838 11268 15844 11280
rect 15427 11240 15844 11268
rect 15427 11237 15439 11240
rect 15381 11231 15439 11237
rect 15838 11228 15844 11240
rect 15896 11228 15902 11280
rect 13170 11200 13176 11212
rect 13131 11172 13176 11200
rect 13170 11160 13176 11172
rect 13228 11160 13234 11212
rect 13814 11200 13820 11212
rect 13280 11172 13820 11200
rect 11572 11104 12296 11132
rect 11572 11092 11578 11104
rect 12342 11092 12348 11144
rect 12400 11132 12406 11144
rect 13280 11132 13308 11172
rect 13814 11160 13820 11172
rect 13872 11200 13878 11212
rect 14001 11203 14059 11209
rect 14001 11200 14013 11203
rect 13872 11172 14013 11200
rect 13872 11160 13878 11172
rect 14001 11169 14013 11172
rect 14047 11169 14059 11203
rect 14001 11163 14059 11169
rect 14369 11203 14427 11209
rect 14369 11169 14381 11203
rect 14415 11169 14427 11203
rect 14550 11200 14556 11212
rect 14511 11172 14556 11200
rect 14369 11163 14427 11169
rect 12400 11104 13308 11132
rect 12400 11092 12406 11104
rect 5537 11067 5595 11073
rect 2976 11036 5488 11064
rect 2501 11027 2559 11033
rect 5460 10996 5488 11036
rect 5537 11033 5549 11067
rect 5583 11064 5595 11067
rect 5629 11067 5687 11073
rect 5629 11064 5641 11067
rect 5583 11036 5641 11064
rect 5583 11033 5595 11036
rect 5537 11027 5595 11033
rect 5629 11033 5641 11036
rect 5675 11033 5687 11067
rect 5629 11027 5687 11033
rect 7377 11067 7435 11073
rect 7377 11033 7389 11067
rect 7423 11033 7435 11067
rect 7377 11027 7435 11033
rect 7466 11024 7472 11076
rect 7524 11064 7530 11076
rect 8386 11064 8392 11076
rect 7524 11036 8392 11064
rect 7524 11024 7530 11036
rect 8386 11024 8392 11036
rect 8444 11064 8450 11076
rect 8573 11067 8631 11073
rect 8573 11064 8585 11067
rect 8444 11036 8585 11064
rect 8444 11024 8450 11036
rect 8573 11033 8585 11036
rect 8619 11033 8631 11067
rect 8573 11027 8631 11033
rect 8757 11067 8815 11073
rect 8757 11033 8769 11067
rect 8803 11064 8815 11067
rect 9766 11064 9772 11076
rect 8803 11036 9772 11064
rect 8803 11033 8815 11036
rect 8757 11027 8815 11033
rect 9766 11024 9772 11036
rect 9824 11024 9830 11076
rect 10689 11067 10747 11073
rect 10689 11033 10701 11067
rect 10735 11064 10747 11067
rect 11422 11064 11428 11076
rect 10735 11036 11428 11064
rect 10735 11033 10747 11036
rect 10689 11027 10747 11033
rect 11422 11024 11428 11036
rect 11480 11024 11486 11076
rect 11790 11064 11796 11076
rect 11703 11036 11796 11064
rect 11790 11024 11796 11036
rect 11848 11064 11854 11076
rect 11974 11064 11980 11076
rect 11848 11036 11980 11064
rect 11848 11024 11854 11036
rect 11974 11024 11980 11036
rect 12032 11024 12038 11076
rect 14384 11064 14412 11163
rect 14550 11160 14556 11172
rect 14608 11160 14614 11212
rect 15102 11160 15108 11212
rect 15160 11200 15166 11212
rect 15473 11203 15531 11209
rect 15473 11200 15485 11203
rect 15160 11172 15485 11200
rect 15160 11160 15166 11172
rect 15473 11169 15485 11172
rect 15519 11169 15531 11203
rect 16482 11200 16488 11212
rect 16443 11172 16488 11200
rect 15473 11163 15531 11169
rect 16482 11160 16488 11172
rect 16540 11160 16546 11212
rect 14918 11064 14924 11076
rect 13280 11036 14412 11064
rect 14879 11036 14924 11064
rect 13280 11008 13308 11036
rect 14918 11024 14924 11036
rect 14976 11024 14982 11076
rect 6454 10996 6460 11008
rect 5460 10968 6460 10996
rect 6454 10956 6460 10968
rect 6512 10956 6518 11008
rect 8202 10996 8208 11008
rect 8163 10968 8208 10996
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 8478 10956 8484 11008
rect 8536 10996 8542 11008
rect 8665 10999 8723 11005
rect 8665 10996 8677 10999
rect 8536 10968 8677 10996
rect 8536 10956 8542 10968
rect 8665 10965 8677 10968
rect 8711 10965 8723 10999
rect 11606 10996 11612 11008
rect 11567 10968 11612 10996
rect 8665 10959 8723 10965
rect 11606 10956 11612 10968
rect 11664 10956 11670 11008
rect 13262 10996 13268 11008
rect 13223 10968 13268 10996
rect 13262 10956 13268 10968
rect 13320 10956 13326 11008
rect 1104 10906 16836 10928
rect 1104 10854 3604 10906
rect 3656 10854 3668 10906
rect 3720 10854 3732 10906
rect 3784 10854 3796 10906
rect 3848 10854 8848 10906
rect 8900 10854 8912 10906
rect 8964 10854 8976 10906
rect 9028 10854 9040 10906
rect 9092 10854 14092 10906
rect 14144 10854 14156 10906
rect 14208 10854 14220 10906
rect 14272 10854 14284 10906
rect 14336 10854 16836 10906
rect 1104 10832 16836 10854
rect 6454 10792 6460 10804
rect 6415 10764 6460 10792
rect 6454 10752 6460 10764
rect 6512 10752 6518 10804
rect 6638 10752 6644 10804
rect 6696 10792 6702 10804
rect 6825 10795 6883 10801
rect 6825 10792 6837 10795
rect 6696 10764 6837 10792
rect 6696 10752 6702 10764
rect 6825 10761 6837 10764
rect 6871 10761 6883 10795
rect 6825 10755 6883 10761
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7282 10792 7288 10804
rect 6972 10764 7017 10792
rect 7243 10764 7288 10792
rect 6972 10752 6978 10764
rect 7282 10752 7288 10764
rect 7340 10752 7346 10804
rect 7742 10752 7748 10804
rect 7800 10792 7806 10804
rect 8113 10795 8171 10801
rect 8113 10792 8125 10795
rect 7800 10764 8125 10792
rect 7800 10752 7806 10764
rect 8113 10761 8125 10764
rect 8159 10761 8171 10795
rect 8113 10755 8171 10761
rect 8941 10795 8999 10801
rect 8941 10761 8953 10795
rect 8987 10792 8999 10795
rect 9214 10792 9220 10804
rect 8987 10764 9220 10792
rect 8987 10761 8999 10764
rect 8941 10755 8999 10761
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 9401 10795 9459 10801
rect 9401 10761 9413 10795
rect 9447 10792 9459 10795
rect 10134 10792 10140 10804
rect 9447 10764 10140 10792
rect 9447 10761 9459 10764
rect 9401 10755 9459 10761
rect 3697 10727 3755 10733
rect 3697 10693 3709 10727
rect 3743 10693 3755 10727
rect 3697 10687 3755 10693
rect 4341 10727 4399 10733
rect 4341 10693 4353 10727
rect 4387 10724 4399 10727
rect 4798 10724 4804 10736
rect 4387 10696 4804 10724
rect 4387 10693 4399 10696
rect 4341 10687 4399 10693
rect 3142 10656 3148 10668
rect 3103 10628 3148 10656
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 3712 10656 3740 10687
rect 4798 10684 4804 10696
rect 4856 10684 4862 10736
rect 5994 10684 6000 10736
rect 6052 10684 6058 10736
rect 6089 10727 6147 10733
rect 6089 10693 6101 10727
rect 6135 10724 6147 10727
rect 6932 10724 6960 10752
rect 6135 10696 6960 10724
rect 8481 10727 8539 10733
rect 6135 10693 6147 10696
rect 6089 10687 6147 10693
rect 8481 10693 8493 10727
rect 8527 10724 8539 10727
rect 8662 10724 8668 10736
rect 8527 10696 8668 10724
rect 8527 10693 8539 10696
rect 8481 10687 8539 10693
rect 8662 10684 8668 10696
rect 8720 10684 8726 10736
rect 9416 10724 9444 10755
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 10367 10795 10425 10801
rect 10367 10761 10379 10795
rect 10413 10792 10425 10795
rect 11146 10792 11152 10804
rect 10413 10764 11152 10792
rect 10413 10761 10425 10764
rect 10367 10755 10425 10761
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 11606 10752 11612 10804
rect 11664 10792 11670 10804
rect 12342 10792 12348 10804
rect 11664 10764 12348 10792
rect 11664 10752 11670 10764
rect 12342 10752 12348 10764
rect 12400 10792 12406 10804
rect 12805 10795 12863 10801
rect 12805 10792 12817 10795
rect 12400 10764 12817 10792
rect 12400 10752 12406 10764
rect 8772 10696 9444 10724
rect 9493 10727 9551 10733
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 3712 10628 4445 10656
rect 1949 10591 2007 10597
rect 1949 10557 1961 10591
rect 1995 10588 2007 10591
rect 2130 10588 2136 10600
rect 1995 10560 2136 10588
rect 1995 10557 2007 10560
rect 1949 10551 2007 10557
rect 2130 10548 2136 10560
rect 2188 10548 2194 10600
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 3804 10597 3832 10628
rect 4433 10625 4445 10628
rect 4479 10625 4491 10659
rect 6012 10656 6040 10684
rect 6546 10656 6552 10668
rect 6012 10628 6552 10656
rect 4433 10619 4491 10625
rect 6546 10616 6552 10628
rect 6604 10656 6610 10668
rect 7926 10656 7932 10668
rect 6604 10628 7932 10656
rect 6604 10616 6610 10628
rect 7926 10616 7932 10628
rect 7984 10616 7990 10668
rect 8386 10656 8392 10668
rect 8299 10628 8392 10656
rect 8386 10616 8392 10628
rect 8444 10656 8450 10668
rect 8772 10656 8800 10696
rect 9493 10693 9505 10727
rect 9539 10724 9551 10727
rect 9582 10724 9588 10736
rect 9539 10696 9588 10724
rect 9539 10693 9551 10696
rect 9493 10687 9551 10693
rect 9582 10684 9588 10696
rect 9640 10684 9646 10736
rect 10226 10724 10232 10736
rect 10187 10696 10232 10724
rect 10226 10684 10232 10696
rect 10284 10684 10290 10736
rect 11514 10724 11520 10736
rect 10336 10696 11520 10724
rect 8444 10628 8800 10656
rect 8444 10616 8450 10628
rect 8846 10616 8852 10668
rect 8904 10656 8910 10668
rect 10137 10659 10195 10665
rect 10137 10656 10149 10659
rect 8904 10628 10149 10656
rect 8904 10616 8910 10628
rect 10137 10625 10149 10628
rect 10183 10656 10195 10659
rect 10336 10656 10364 10696
rect 11514 10684 11520 10696
rect 11572 10684 11578 10736
rect 11698 10724 11704 10736
rect 11659 10696 11704 10724
rect 11698 10684 11704 10696
rect 11756 10684 11762 10736
rect 10183 10628 10364 10656
rect 10183 10625 10195 10628
rect 10137 10619 10195 10625
rect 10410 10616 10416 10668
rect 10468 10656 10474 10668
rect 10468 10628 10824 10656
rect 10468 10616 10474 10628
rect 3789 10591 3847 10597
rect 2832 10560 2877 10588
rect 2832 10548 2838 10560
rect 3789 10557 3801 10591
rect 3835 10557 3847 10591
rect 4338 10588 4344 10600
rect 4299 10560 4344 10588
rect 3789 10551 3847 10557
rect 4338 10548 4344 10560
rect 4396 10548 4402 10600
rect 4801 10591 4859 10597
rect 4801 10557 4813 10591
rect 4847 10588 4859 10591
rect 4893 10591 4951 10597
rect 4893 10588 4905 10591
rect 4847 10560 4905 10588
rect 4847 10557 4859 10560
rect 4801 10551 4859 10557
rect 4893 10557 4905 10560
rect 4939 10557 4951 10591
rect 5074 10588 5080 10600
rect 5035 10560 5080 10588
rect 4893 10551 4951 10557
rect 5074 10548 5080 10560
rect 5132 10548 5138 10600
rect 5905 10591 5963 10597
rect 5905 10557 5917 10591
rect 5951 10557 5963 10591
rect 5905 10551 5963 10557
rect 2222 10480 2228 10532
rect 2280 10520 2286 10532
rect 2593 10523 2651 10529
rect 2593 10520 2605 10523
rect 2280 10492 2605 10520
rect 2280 10480 2286 10492
rect 2593 10489 2605 10492
rect 2639 10489 2651 10523
rect 5721 10523 5779 10529
rect 5721 10520 5733 10523
rect 2593 10483 2651 10489
rect 4448 10492 5733 10520
rect 3234 10452 3240 10464
rect 3195 10424 3240 10452
rect 3234 10412 3240 10424
rect 3292 10412 3298 10464
rect 3329 10455 3387 10461
rect 3329 10421 3341 10455
rect 3375 10452 3387 10455
rect 4448 10452 4476 10492
rect 5721 10489 5733 10492
rect 5767 10489 5779 10523
rect 5920 10520 5948 10551
rect 5994 10548 6000 10600
rect 6052 10588 6058 10600
rect 6178 10588 6184 10600
rect 6052 10560 6097 10588
rect 6139 10560 6184 10588
rect 6052 10548 6058 10560
rect 6178 10548 6184 10560
rect 6236 10588 6242 10600
rect 6733 10591 6791 10597
rect 6733 10588 6745 10591
rect 6236 10560 6745 10588
rect 6236 10548 6242 10560
rect 6733 10557 6745 10560
rect 6779 10557 6791 10591
rect 7006 10588 7012 10600
rect 6967 10560 7012 10588
rect 6733 10551 6791 10557
rect 7006 10548 7012 10560
rect 7064 10548 7070 10600
rect 7190 10588 7196 10600
rect 7151 10560 7196 10588
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 7653 10591 7711 10597
rect 7653 10557 7665 10591
rect 7699 10588 7711 10591
rect 8202 10588 8208 10600
rect 7699 10560 8208 10588
rect 7699 10557 7711 10560
rect 7653 10551 7711 10557
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 8297 10591 8355 10597
rect 8297 10557 8309 10591
rect 8343 10557 8355 10591
rect 8570 10588 8576 10600
rect 8531 10560 8576 10588
rect 8297 10551 8355 10557
rect 7208 10520 7236 10548
rect 5920 10492 7236 10520
rect 8312 10520 8340 10551
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 8757 10591 8815 10597
rect 8757 10557 8769 10591
rect 8803 10588 8815 10591
rect 9030 10588 9036 10600
rect 8803 10560 9036 10588
rect 8803 10557 8815 10560
rect 8757 10551 8815 10557
rect 9030 10548 9036 10560
rect 9088 10548 9094 10600
rect 9214 10588 9220 10600
rect 9175 10560 9220 10588
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 9309 10591 9367 10597
rect 9309 10557 9321 10591
rect 9355 10557 9367 10591
rect 9674 10588 9680 10600
rect 9635 10560 9680 10588
rect 9309 10551 9367 10557
rect 8478 10520 8484 10532
rect 8312 10492 8484 10520
rect 5721 10483 5779 10489
rect 8478 10480 8484 10492
rect 8536 10520 8542 10532
rect 9324 10520 9352 10551
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 9858 10548 9864 10600
rect 9916 10588 9922 10600
rect 10796 10597 10824 10628
rect 10870 10616 10876 10668
rect 10928 10656 10934 10668
rect 12161 10659 12219 10665
rect 10928 10628 11744 10656
rect 10928 10616 10934 10628
rect 10597 10591 10655 10597
rect 10597 10588 10609 10591
rect 9916 10560 10609 10588
rect 9916 10548 9922 10560
rect 10597 10557 10609 10560
rect 10643 10557 10655 10591
rect 10597 10551 10655 10557
rect 10781 10591 10839 10597
rect 10781 10557 10793 10591
rect 10827 10557 10839 10591
rect 11146 10588 11152 10600
rect 11107 10560 11152 10588
rect 10781 10551 10839 10557
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 11422 10588 11428 10600
rect 11383 10560 11428 10588
rect 11422 10548 11428 10560
rect 11480 10548 11486 10600
rect 11716 10597 11744 10628
rect 12161 10625 12173 10659
rect 12207 10656 12219 10659
rect 12250 10656 12256 10668
rect 12207 10628 12256 10656
rect 12207 10625 12219 10628
rect 12161 10619 12219 10625
rect 12250 10616 12256 10628
rect 12308 10616 12314 10668
rect 11701 10591 11759 10597
rect 11701 10557 11713 10591
rect 11747 10557 11759 10591
rect 11701 10551 11759 10557
rect 11885 10591 11943 10597
rect 11885 10557 11897 10591
rect 11931 10557 11943 10591
rect 12434 10588 12440 10600
rect 12395 10560 12440 10588
rect 11885 10551 11943 10557
rect 8536 10492 9352 10520
rect 8536 10480 8542 10492
rect 4798 10452 4804 10464
rect 3375 10424 4476 10452
rect 4759 10424 4804 10452
rect 3375 10421 3387 10424
rect 3329 10415 3387 10421
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 6638 10452 6644 10464
rect 5592 10424 6644 10452
rect 5592 10412 5598 10424
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 7742 10452 7748 10464
rect 7703 10424 7748 10452
rect 7742 10412 7748 10424
rect 7800 10412 7806 10464
rect 9324 10452 9352 10492
rect 9490 10480 9496 10532
rect 9548 10520 9554 10532
rect 9769 10523 9827 10529
rect 9769 10520 9781 10523
rect 9548 10492 9781 10520
rect 9548 10480 9554 10492
rect 9769 10489 9781 10492
rect 9815 10489 9827 10523
rect 9769 10483 9827 10489
rect 10505 10523 10563 10529
rect 10505 10489 10517 10523
rect 10551 10520 10563 10523
rect 10686 10520 10692 10532
rect 10551 10492 10692 10520
rect 10551 10489 10563 10492
rect 10505 10483 10563 10489
rect 10520 10452 10548 10483
rect 10686 10480 10692 10492
rect 10744 10480 10750 10532
rect 11900 10520 11928 10551
rect 12434 10548 12440 10560
rect 12492 10548 12498 10600
rect 12636 10597 12664 10764
rect 12805 10761 12817 10764
rect 12851 10761 12863 10795
rect 12805 10755 12863 10761
rect 14458 10656 14464 10668
rect 14419 10628 14464 10656
rect 14458 10616 14464 10628
rect 14516 10616 14522 10668
rect 12621 10591 12679 10597
rect 12621 10557 12633 10591
rect 12667 10557 12679 10591
rect 12621 10551 12679 10557
rect 12710 10548 12716 10600
rect 12768 10588 12774 10600
rect 12897 10591 12955 10597
rect 12897 10588 12909 10591
rect 12768 10560 12909 10588
rect 12768 10548 12774 10560
rect 12897 10557 12909 10560
rect 12943 10588 12955 10591
rect 13078 10588 13084 10600
rect 12943 10560 13084 10588
rect 12943 10557 12955 10560
rect 12897 10551 12955 10557
rect 13078 10548 13084 10560
rect 13136 10548 13142 10600
rect 13354 10548 13360 10600
rect 13412 10588 13418 10600
rect 14185 10591 14243 10597
rect 14185 10588 14197 10591
rect 13412 10560 14197 10588
rect 13412 10548 13418 10560
rect 14185 10557 14197 10560
rect 14231 10557 14243 10591
rect 14185 10551 14243 10557
rect 14277 10591 14335 10597
rect 14277 10557 14289 10591
rect 14323 10588 14335 10591
rect 14642 10588 14648 10600
rect 14323 10560 14648 10588
rect 14323 10557 14335 10560
rect 14277 10551 14335 10557
rect 14642 10548 14648 10560
rect 14700 10548 14706 10600
rect 15654 10588 15660 10600
rect 15615 10560 15660 10588
rect 15654 10548 15660 10560
rect 15712 10548 15718 10600
rect 11348 10492 11928 10520
rect 11348 10464 11376 10492
rect 11146 10452 11152 10464
rect 9324 10424 11152 10452
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 11330 10452 11336 10464
rect 11291 10424 11336 10452
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 14461 10455 14519 10461
rect 14461 10421 14473 10455
rect 14507 10452 14519 10455
rect 14918 10452 14924 10464
rect 14507 10424 14924 10452
rect 14507 10421 14519 10424
rect 14461 10415 14519 10421
rect 14918 10412 14924 10424
rect 14976 10412 14982 10464
rect 15841 10455 15899 10461
rect 15841 10421 15853 10455
rect 15887 10452 15899 10455
rect 15930 10452 15936 10464
rect 15887 10424 15936 10452
rect 15887 10421 15899 10424
rect 15841 10415 15899 10421
rect 15930 10412 15936 10424
rect 15988 10412 15994 10464
rect 1104 10362 16836 10384
rect 1104 10310 6226 10362
rect 6278 10310 6290 10362
rect 6342 10310 6354 10362
rect 6406 10310 6418 10362
rect 6470 10310 11470 10362
rect 11522 10310 11534 10362
rect 11586 10310 11598 10362
rect 11650 10310 11662 10362
rect 11714 10310 16836 10362
rect 1104 10288 16836 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 3234 10248 3240 10260
rect 1627 10220 3240 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 3234 10208 3240 10220
rect 3292 10208 3298 10260
rect 5994 10208 6000 10260
rect 6052 10248 6058 10260
rect 6730 10248 6736 10260
rect 6052 10220 6736 10248
rect 6052 10208 6058 10220
rect 6730 10208 6736 10220
rect 6788 10248 6794 10260
rect 7006 10248 7012 10260
rect 6788 10220 7012 10248
rect 6788 10208 6794 10220
rect 7006 10208 7012 10220
rect 7064 10248 7070 10260
rect 10226 10248 10232 10260
rect 7064 10220 10232 10248
rect 7064 10208 7070 10220
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 6638 10140 6644 10192
rect 6696 10180 6702 10192
rect 10778 10180 10784 10192
rect 6696 10152 10784 10180
rect 6696 10140 6702 10152
rect 10778 10140 10784 10152
rect 10836 10180 10842 10192
rect 11330 10180 11336 10192
rect 10836 10152 11336 10180
rect 10836 10140 10842 10152
rect 11330 10140 11336 10152
rect 11388 10140 11394 10192
rect 12713 10183 12771 10189
rect 12713 10149 12725 10183
rect 12759 10180 12771 10183
rect 14918 10180 14924 10192
rect 12759 10152 14412 10180
rect 14879 10152 14924 10180
rect 12759 10149 12771 10152
rect 12713 10143 12771 10149
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 2130 10112 2136 10124
rect 2091 10084 2136 10112
rect 2130 10072 2136 10084
rect 2188 10072 2194 10124
rect 3142 10072 3148 10124
rect 3200 10112 3206 10124
rect 3237 10115 3295 10121
rect 3237 10112 3249 10115
rect 3200 10084 3249 10112
rect 3200 10072 3206 10084
rect 3237 10081 3249 10084
rect 3283 10112 3295 10115
rect 6546 10112 6552 10124
rect 3283 10084 6552 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 12342 10072 12348 10124
rect 12400 10112 12406 10124
rect 12437 10115 12495 10121
rect 12437 10112 12449 10115
rect 12400 10084 12449 10112
rect 12400 10072 12406 10084
rect 12437 10081 12449 10084
rect 12483 10081 12495 10115
rect 12437 10075 12495 10081
rect 13354 10072 13360 10124
rect 13412 10112 13418 10124
rect 13449 10115 13507 10121
rect 13449 10112 13461 10115
rect 13412 10084 13461 10112
rect 13412 10072 13418 10084
rect 13449 10081 13461 10084
rect 13495 10081 13507 10115
rect 13449 10075 13507 10081
rect 13725 10115 13783 10121
rect 13725 10081 13737 10115
rect 13771 10081 13783 10115
rect 13725 10075 13783 10081
rect 2314 10044 2320 10056
rect 2275 10016 2320 10044
rect 2314 10004 2320 10016
rect 2372 10004 2378 10056
rect 12710 10044 12716 10056
rect 12671 10016 12716 10044
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 13078 10004 13084 10056
rect 13136 10044 13142 10056
rect 13740 10044 13768 10075
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 14384 10121 14412 10152
rect 14918 10140 14924 10152
rect 14976 10140 14982 10192
rect 15930 10140 15936 10192
rect 15988 10140 15994 10192
rect 14369 10115 14427 10121
rect 13872 10084 13917 10112
rect 13872 10072 13878 10084
rect 14369 10081 14381 10115
rect 14415 10112 14427 10115
rect 14550 10112 14556 10124
rect 14415 10084 14556 10112
rect 14415 10081 14427 10084
rect 14369 10075 14427 10081
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 13136 10016 13768 10044
rect 13832 10044 13860 10072
rect 14645 10047 14703 10053
rect 13832 10016 14596 10044
rect 13136 10004 13142 10016
rect 11054 9936 11060 9988
rect 11112 9976 11118 9988
rect 12250 9976 12256 9988
rect 11112 9948 12256 9976
rect 11112 9936 11118 9948
rect 12250 9936 12256 9948
rect 12308 9976 12314 9988
rect 13541 9979 13599 9985
rect 13541 9976 13553 9979
rect 12308 9948 13553 9976
rect 12308 9936 12314 9948
rect 13541 9945 13553 9948
rect 13587 9945 13599 9979
rect 13541 9939 13599 9945
rect 13906 9936 13912 9988
rect 13964 9976 13970 9988
rect 14461 9979 14519 9985
rect 14461 9976 14473 9979
rect 13964 9948 14473 9976
rect 13964 9936 13970 9948
rect 14461 9945 14473 9948
rect 14507 9945 14519 9979
rect 14461 9939 14519 9945
rect 12526 9908 12532 9920
rect 12487 9880 12532 9908
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 14001 9911 14059 9917
rect 14001 9908 14013 9911
rect 13872 9880 14013 9908
rect 13872 9868 13878 9880
rect 14001 9877 14013 9880
rect 14047 9877 14059 9911
rect 14568 9908 14596 10016
rect 14645 10013 14657 10047
rect 14691 10044 14703 10047
rect 14918 10044 14924 10056
rect 14691 10016 14924 10044
rect 14691 10013 14703 10016
rect 14645 10007 14703 10013
rect 14918 10004 14924 10016
rect 14976 10004 14982 10056
rect 16393 9911 16451 9917
rect 16393 9908 16405 9911
rect 14568 9880 16405 9908
rect 14001 9871 14059 9877
rect 16393 9877 16405 9880
rect 16439 9877 16451 9911
rect 16393 9871 16451 9877
rect 1104 9818 16836 9840
rect 1104 9766 3604 9818
rect 3656 9766 3668 9818
rect 3720 9766 3732 9818
rect 3784 9766 3796 9818
rect 3848 9766 8848 9818
rect 8900 9766 8912 9818
rect 8964 9766 8976 9818
rect 9028 9766 9040 9818
rect 9092 9766 14092 9818
rect 14144 9766 14156 9818
rect 14208 9766 14220 9818
rect 14272 9766 14284 9818
rect 14336 9766 16836 9818
rect 1104 9744 16836 9766
rect 12526 9704 12532 9716
rect 12084 9676 12532 9704
rect 4525 9639 4583 9645
rect 4525 9605 4537 9639
rect 4571 9636 4583 9639
rect 5626 9636 5632 9648
rect 4571 9608 5632 9636
rect 4571 9605 4583 9608
rect 4525 9599 4583 9605
rect 5626 9596 5632 9608
rect 5684 9596 5690 9648
rect 7834 9596 7840 9648
rect 7892 9636 7898 9648
rect 8205 9639 8263 9645
rect 8205 9636 8217 9639
rect 7892 9608 8217 9636
rect 7892 9596 7898 9608
rect 8205 9605 8217 9608
rect 8251 9605 8263 9639
rect 8205 9599 8263 9605
rect 10597 9639 10655 9645
rect 10597 9605 10609 9639
rect 10643 9636 10655 9639
rect 11238 9636 11244 9648
rect 10643 9608 11244 9636
rect 10643 9605 10655 9608
rect 10597 9599 10655 9605
rect 11238 9596 11244 9608
rect 11296 9596 11302 9648
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2774 9568 2780 9580
rect 2547 9540 2780 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2774 9528 2780 9540
rect 2832 9528 2838 9580
rect 4706 9568 4712 9580
rect 4540 9540 4712 9568
rect 2222 9500 2228 9512
rect 2183 9472 2228 9500
rect 2222 9460 2228 9472
rect 2280 9460 2286 9512
rect 3513 9503 3571 9509
rect 3513 9469 3525 9503
rect 3559 9500 3571 9503
rect 3602 9500 3608 9512
rect 3559 9472 3608 9500
rect 3559 9469 3571 9472
rect 3513 9463 3571 9469
rect 3602 9460 3608 9472
rect 3660 9460 3666 9512
rect 3878 9500 3884 9512
rect 3839 9472 3884 9500
rect 3878 9460 3884 9472
rect 3936 9460 3942 9512
rect 4540 9509 4568 9540
rect 4706 9528 4712 9540
rect 4764 9568 4770 9580
rect 5169 9571 5227 9577
rect 5169 9568 5181 9571
rect 4764 9540 5181 9568
rect 4764 9528 4770 9540
rect 5169 9537 5181 9540
rect 5215 9537 5227 9571
rect 5169 9531 5227 9537
rect 6457 9571 6515 9577
rect 6457 9537 6469 9571
rect 6503 9568 6515 9571
rect 7098 9568 7104 9580
rect 6503 9540 7104 9568
rect 6503 9537 6515 9540
rect 6457 9531 6515 9537
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 10060 9540 10916 9568
rect 10060 9512 10088 9540
rect 10888 9512 10916 9540
rect 10962 9528 10968 9580
rect 11020 9568 11026 9580
rect 11057 9571 11115 9577
rect 11057 9568 11069 9571
rect 11020 9540 11069 9568
rect 11020 9528 11026 9540
rect 11057 9537 11069 9540
rect 11103 9537 11115 9571
rect 11057 9531 11115 9537
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9469 4583 9503
rect 4525 9463 4583 9469
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9500 5135 9503
rect 5534 9500 5540 9512
rect 5123 9472 5540 9500
rect 5123 9469 5135 9472
rect 5077 9463 5135 9469
rect 5534 9460 5540 9472
rect 5592 9460 5598 9512
rect 10042 9500 10048 9512
rect 9955 9472 10048 9500
rect 10042 9460 10048 9472
rect 10100 9460 10106 9512
rect 10459 9503 10517 9509
rect 10459 9469 10471 9503
rect 10505 9500 10517 9503
rect 10870 9500 10876 9512
rect 10505 9472 10640 9500
rect 10831 9472 10876 9500
rect 10505 9469 10517 9472
rect 10459 9463 10517 9469
rect 4798 9392 4804 9444
rect 4856 9432 4862 9444
rect 5353 9435 5411 9441
rect 5353 9432 5365 9435
rect 4856 9404 5365 9432
rect 4856 9392 4862 9404
rect 5353 9401 5365 9404
rect 5399 9401 5411 9435
rect 5353 9395 5411 9401
rect 6733 9435 6791 9441
rect 6733 9401 6745 9435
rect 6779 9432 6791 9435
rect 6822 9432 6828 9444
rect 6779 9404 6828 9432
rect 6779 9401 6791 9404
rect 6733 9395 6791 9401
rect 6822 9392 6828 9404
rect 6880 9392 6886 9444
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 7064 9404 7222 9432
rect 7064 9392 7070 9404
rect 9582 9392 9588 9444
rect 9640 9432 9646 9444
rect 10229 9435 10287 9441
rect 10229 9432 10241 9435
rect 9640 9404 10241 9432
rect 9640 9392 9646 9404
rect 10229 9401 10241 9404
rect 10275 9401 10287 9435
rect 10229 9395 10287 9401
rect 10321 9435 10379 9441
rect 10321 9401 10333 9435
rect 10367 9401 10379 9435
rect 10321 9395 10379 9401
rect 10612 9432 10640 9472
rect 10870 9460 10876 9472
rect 10928 9460 10934 9512
rect 11149 9503 11207 9509
rect 11149 9469 11161 9503
rect 11195 9469 11207 9503
rect 11149 9463 11207 9469
rect 11333 9503 11391 9509
rect 11333 9469 11345 9503
rect 11379 9500 11391 9503
rect 11790 9500 11796 9512
rect 11379 9472 11796 9500
rect 11379 9469 11391 9472
rect 11333 9463 11391 9469
rect 11054 9432 11060 9444
rect 10612 9404 11060 9432
rect 2038 9364 2044 9376
rect 1999 9336 2044 9364
rect 2038 9324 2044 9336
rect 2096 9324 2102 9376
rect 3881 9367 3939 9373
rect 3881 9333 3893 9367
rect 3927 9364 3939 9367
rect 4338 9364 4344 9376
rect 3927 9336 4344 9364
rect 3927 9333 3939 9336
rect 3881 9327 3939 9333
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 9766 9324 9772 9376
rect 9824 9364 9830 9376
rect 10336 9364 10364 9395
rect 9824 9336 10364 9364
rect 9824 9324 9830 9336
rect 10410 9324 10416 9376
rect 10468 9364 10474 9376
rect 10612 9364 10640 9404
rect 11054 9392 11060 9404
rect 11112 9392 11118 9444
rect 11164 9432 11192 9463
rect 11790 9460 11796 9472
rect 11848 9460 11854 9512
rect 11882 9460 11888 9512
rect 11940 9500 11946 9512
rect 11977 9503 12035 9509
rect 11977 9500 11989 9503
rect 11940 9472 11989 9500
rect 11940 9460 11946 9472
rect 11977 9469 11989 9472
rect 12023 9500 12035 9503
rect 12084 9500 12112 9676
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 12621 9707 12679 9713
rect 12621 9673 12633 9707
rect 12667 9704 12679 9707
rect 12710 9704 12716 9716
rect 12667 9676 12716 9704
rect 12667 9673 12679 9676
rect 12621 9667 12679 9673
rect 12710 9664 12716 9676
rect 12768 9664 12774 9716
rect 14458 9704 14464 9716
rect 14419 9676 14464 9704
rect 14458 9664 14464 9676
rect 14516 9664 14522 9716
rect 12342 9636 12348 9648
rect 12176 9608 12348 9636
rect 12176 9509 12204 9608
rect 12342 9596 12348 9608
rect 12400 9596 12406 9648
rect 12544 9636 12572 9664
rect 13078 9636 13084 9648
rect 12544 9608 13084 9636
rect 13078 9596 13084 9608
rect 13136 9596 13142 9648
rect 13449 9639 13507 9645
rect 13449 9605 13461 9639
rect 13495 9636 13507 9639
rect 13814 9636 13820 9648
rect 13495 9608 13820 9636
rect 13495 9605 13507 9608
rect 13449 9599 13507 9605
rect 13814 9596 13820 9608
rect 13872 9636 13878 9648
rect 13872 9608 14136 9636
rect 13872 9596 13878 9608
rect 13170 9568 13176 9580
rect 12452 9540 13176 9568
rect 12023 9472 12112 9500
rect 12161 9503 12219 9509
rect 12023 9469 12035 9472
rect 11977 9463 12035 9469
rect 12161 9469 12173 9503
rect 12207 9469 12219 9503
rect 12342 9500 12348 9512
rect 12303 9472 12348 9500
rect 12161 9463 12219 9469
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 11164 9404 11376 9432
rect 11348 9376 11376 9404
rect 12066 9392 12072 9444
rect 12124 9432 12130 9444
rect 12253 9435 12311 9441
rect 12253 9432 12265 9435
rect 12124 9404 12265 9432
rect 12124 9392 12130 9404
rect 12253 9401 12265 9404
rect 12299 9401 12311 9435
rect 12253 9395 12311 9401
rect 10468 9336 10640 9364
rect 10468 9324 10474 9336
rect 11330 9324 11336 9376
rect 11388 9324 11394 9376
rect 11517 9367 11575 9373
rect 11517 9333 11529 9367
rect 11563 9364 11575 9367
rect 12452 9364 12480 9540
rect 12820 9509 12848 9540
rect 13170 9528 13176 9540
rect 13228 9568 13234 9580
rect 13357 9571 13415 9577
rect 13357 9568 13369 9571
rect 13228 9540 13369 9568
rect 13228 9528 13234 9540
rect 13357 9537 13369 9540
rect 13403 9537 13415 9571
rect 13357 9531 13415 9537
rect 14108 9568 14136 9608
rect 14108 9540 14596 9568
rect 12805 9503 12863 9509
rect 12805 9469 12817 9503
rect 12851 9469 12863 9503
rect 13078 9500 13084 9512
rect 13039 9472 13084 9500
rect 12805 9463 12863 9469
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 13262 9500 13268 9512
rect 13223 9472 13268 9500
rect 13262 9460 13268 9472
rect 13320 9460 13326 9512
rect 13541 9503 13599 9509
rect 13541 9469 13553 9503
rect 13587 9469 13599 9503
rect 13541 9463 13599 9469
rect 12989 9435 13047 9441
rect 12989 9401 13001 9435
rect 13035 9432 13047 9435
rect 13354 9432 13360 9444
rect 13035 9404 13360 9432
rect 13035 9401 13047 9404
rect 12989 9395 13047 9401
rect 11563 9336 12480 9364
rect 12529 9367 12587 9373
rect 11563 9333 11575 9336
rect 11517 9327 11575 9333
rect 12529 9333 12541 9367
rect 12575 9364 12587 9367
rect 13004 9364 13032 9395
rect 13354 9392 13360 9404
rect 13412 9432 13418 9444
rect 13556 9432 13584 9463
rect 13630 9460 13636 9512
rect 13688 9500 13694 9512
rect 13817 9503 13875 9509
rect 13817 9500 13829 9503
rect 13688 9472 13829 9500
rect 13688 9460 13694 9472
rect 13817 9469 13829 9472
rect 13863 9469 13875 9503
rect 13817 9463 13875 9469
rect 13906 9460 13912 9512
rect 13964 9500 13970 9512
rect 14108 9509 14136 9540
rect 14093 9503 14151 9509
rect 13964 9472 14009 9500
rect 13964 9460 13970 9472
rect 14093 9469 14105 9503
rect 14139 9469 14151 9503
rect 14093 9463 14151 9469
rect 14323 9503 14381 9509
rect 14323 9469 14335 9503
rect 14369 9500 14381 9503
rect 14458 9500 14464 9512
rect 14369 9472 14464 9500
rect 14369 9469 14381 9472
rect 14323 9463 14381 9469
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 14568 9509 14596 9540
rect 14553 9503 14611 9509
rect 14553 9469 14565 9503
rect 14599 9469 14611 9503
rect 15562 9500 15568 9512
rect 15523 9472 15568 9500
rect 14553 9463 14611 9469
rect 15562 9460 15568 9472
rect 15620 9460 15626 9512
rect 13412 9404 13584 9432
rect 14185 9435 14243 9441
rect 13412 9392 13418 9404
rect 14185 9401 14197 9435
rect 14231 9432 14243 9435
rect 14645 9435 14703 9441
rect 14645 9432 14657 9435
rect 14231 9404 14657 9432
rect 14231 9401 14243 9404
rect 14185 9395 14243 9401
rect 14645 9401 14657 9404
rect 14691 9401 14703 9435
rect 14645 9395 14703 9401
rect 12575 9336 13032 9364
rect 13725 9367 13783 9373
rect 12575 9333 12587 9336
rect 12529 9327 12587 9333
rect 13725 9333 13737 9367
rect 13771 9364 13783 9367
rect 14550 9364 14556 9376
rect 13771 9336 14556 9364
rect 13771 9333 13783 9336
rect 13725 9327 13783 9333
rect 14550 9324 14556 9336
rect 14608 9324 14614 9376
rect 15654 9324 15660 9376
rect 15712 9364 15718 9376
rect 15749 9367 15807 9373
rect 15749 9364 15761 9367
rect 15712 9336 15761 9364
rect 15712 9324 15718 9336
rect 15749 9333 15761 9336
rect 15795 9333 15807 9367
rect 15749 9327 15807 9333
rect 1104 9274 16836 9296
rect 1104 9222 6226 9274
rect 6278 9222 6290 9274
rect 6342 9222 6354 9274
rect 6406 9222 6418 9274
rect 6470 9222 11470 9274
rect 11522 9222 11534 9274
rect 11586 9222 11598 9274
rect 11650 9222 11662 9274
rect 11714 9222 16836 9274
rect 1104 9200 16836 9222
rect 3602 9160 3608 9172
rect 3563 9132 3608 9160
rect 3602 9120 3608 9132
rect 3660 9120 3666 9172
rect 3878 9120 3884 9172
rect 3936 9160 3942 9172
rect 4525 9163 4583 9169
rect 4525 9160 4537 9163
rect 3936 9132 4537 9160
rect 3936 9120 3942 9132
rect 4525 9129 4537 9132
rect 4571 9129 4583 9163
rect 4525 9123 4583 9129
rect 5534 9120 5540 9172
rect 5592 9160 5598 9172
rect 5813 9163 5871 9169
rect 5813 9160 5825 9163
rect 5592 9132 5825 9160
rect 5592 9120 5598 9132
rect 5813 9129 5825 9132
rect 5859 9129 5871 9163
rect 5813 9123 5871 9129
rect 6086 9120 6092 9172
rect 6144 9160 6150 9172
rect 6181 9163 6239 9169
rect 6181 9160 6193 9163
rect 6144 9132 6193 9160
rect 6144 9120 6150 9132
rect 6181 9129 6193 9132
rect 6227 9129 6239 9163
rect 7006 9160 7012 9172
rect 6967 9132 7012 9160
rect 6181 9123 6239 9129
rect 7006 9120 7012 9132
rect 7064 9120 7070 9172
rect 9214 9160 9220 9172
rect 7760 9132 9220 9160
rect 3142 9052 3148 9104
rect 3200 9052 3206 9104
rect 2038 9024 2044 9036
rect 1999 8996 2044 9024
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 3160 9024 3188 9052
rect 2976 8996 3188 9024
rect 3237 9027 3295 9033
rect 2976 8965 3004 8996
rect 3237 8993 3249 9027
rect 3283 8993 3295 9027
rect 3620 9024 3648 9120
rect 4338 9092 4344 9104
rect 4299 9064 4344 9092
rect 4338 9052 4344 9064
rect 4396 9052 4402 9104
rect 5077 9095 5135 9101
rect 5077 9061 5089 9095
rect 5123 9092 5135 9095
rect 5626 9092 5632 9104
rect 5123 9064 5632 9092
rect 5123 9061 5135 9064
rect 5077 9055 5135 9061
rect 5626 9052 5632 9064
rect 5684 9052 5690 9104
rect 7760 9092 7788 9132
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 9493 9163 9551 9169
rect 9493 9129 9505 9163
rect 9539 9160 9551 9163
rect 9582 9160 9588 9172
rect 9539 9132 9588 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 11609 9163 11667 9169
rect 11609 9160 11621 9163
rect 10612 9132 11621 9160
rect 6104 9064 7788 9092
rect 8864 9064 9536 9092
rect 3881 9027 3939 9033
rect 3881 9024 3893 9027
rect 3620 8996 3893 9024
rect 3237 8987 3295 8993
rect 3881 8993 3893 8996
rect 3927 8993 3939 9027
rect 3881 8987 3939 8993
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 4706 9024 4712 9036
rect 4479 8996 4712 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 2961 8959 3019 8965
rect 2961 8925 2973 8959
rect 3007 8925 3019 8959
rect 3142 8956 3148 8968
rect 3103 8928 3148 8956
rect 2961 8919 3019 8925
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 3252 8888 3280 8987
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 5534 9024 5540 9036
rect 5495 8996 5540 9024
rect 5534 8984 5540 8996
rect 5592 8984 5598 9036
rect 4890 8916 4896 8968
rect 4948 8956 4954 8968
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 4948 8928 4997 8956
rect 4948 8916 4954 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 6104 8888 6132 9064
rect 6730 8984 6736 9036
rect 6788 9024 6794 9036
rect 6825 9027 6883 9033
rect 6825 9024 6837 9027
rect 6788 8996 6837 9024
rect 6788 8984 6794 8996
rect 6825 8993 6837 8996
rect 6871 8993 6883 9027
rect 6825 8987 6883 8993
rect 8478 8984 8484 9036
rect 8536 8984 8542 9036
rect 6273 8959 6331 8965
rect 6273 8925 6285 8959
rect 6319 8925 6331 8959
rect 6273 8919 6331 8925
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8956 6515 8959
rect 6546 8956 6552 8968
rect 6503 8928 6552 8956
rect 6503 8925 6515 8928
rect 6457 8919 6515 8925
rect 3252 8860 6132 8888
rect 2409 8823 2467 8829
rect 2409 8789 2421 8823
rect 2455 8820 2467 8823
rect 2590 8820 2596 8832
rect 2455 8792 2596 8820
rect 2455 8789 2467 8792
rect 2409 8783 2467 8789
rect 2590 8780 2596 8792
rect 2648 8780 2654 8832
rect 6288 8820 6316 8919
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 7098 8956 7104 8968
rect 7059 8928 7104 8956
rect 7098 8916 7104 8928
rect 7156 8916 7162 8968
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8956 7435 8959
rect 8864 8956 8892 9064
rect 9401 9027 9459 9033
rect 9401 8993 9413 9027
rect 9447 8993 9459 9027
rect 9401 8987 9459 8993
rect 7423 8928 8892 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 8849 8891 8907 8897
rect 8849 8857 8861 8891
rect 8895 8888 8907 8891
rect 9416 8888 9444 8987
rect 9508 8956 9536 9064
rect 9600 9024 9628 9120
rect 10152 9064 10548 9092
rect 9907 9027 9965 9033
rect 9907 9024 9919 9027
rect 9600 8996 9919 9024
rect 9907 8993 9919 8996
rect 9953 8993 9965 9027
rect 10042 9024 10048 9036
rect 10003 8996 10048 9024
rect 9907 8987 9965 8993
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 10152 9033 10180 9064
rect 10137 9027 10195 9033
rect 10137 8993 10149 9027
rect 10183 8993 10195 9027
rect 10318 9024 10324 9036
rect 10279 8996 10324 9024
rect 10137 8987 10195 8993
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 10413 8959 10471 8965
rect 10413 8956 10425 8959
rect 9508 8928 10425 8956
rect 10413 8925 10425 8928
rect 10459 8925 10471 8959
rect 10520 8956 10548 9064
rect 10612 9033 10640 9132
rect 11609 9129 11621 9132
rect 11655 9129 11667 9163
rect 11609 9123 11667 9129
rect 11790 9120 11796 9172
rect 11848 9160 11854 9172
rect 14642 9160 14648 9172
rect 11848 9132 14648 9160
rect 11848 9120 11854 9132
rect 10689 9095 10747 9101
rect 10689 9061 10701 9095
rect 10735 9092 10747 9095
rect 11149 9095 11207 9101
rect 11149 9092 11161 9095
rect 10735 9064 11161 9092
rect 10735 9061 10747 9064
rect 10689 9055 10747 9061
rect 11149 9061 11161 9064
rect 11195 9061 11207 9095
rect 11149 9055 11207 9061
rect 11238 9052 11244 9104
rect 11296 9092 11302 9104
rect 11517 9095 11575 9101
rect 11517 9092 11529 9095
rect 11296 9064 11529 9092
rect 11296 9052 11302 9064
rect 11517 9061 11529 9064
rect 11563 9092 11575 9095
rect 11563 9064 11836 9092
rect 11563 9061 11575 9064
rect 11517 9055 11575 9061
rect 10597 9027 10655 9033
rect 10597 8993 10609 9027
rect 10643 8993 10655 9027
rect 10778 9024 10784 9036
rect 10739 8996 10784 9024
rect 10597 8987 10655 8993
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 10899 9027 10957 9033
rect 10899 9024 10911 9027
rect 10888 8993 10911 9024
rect 10945 8993 10957 9027
rect 11330 9024 11336 9036
rect 11291 8996 11336 9024
rect 10888 8987 10957 8993
rect 10796 8956 10824 8984
rect 10520 8928 10824 8956
rect 10413 8919 10471 8925
rect 9766 8888 9772 8900
rect 8895 8860 9772 8888
rect 8895 8857 8907 8860
rect 8849 8851 8907 8857
rect 9766 8848 9772 8860
rect 9824 8888 9830 8900
rect 10226 8888 10232 8900
rect 9824 8860 10232 8888
rect 9824 8848 9830 8860
rect 10226 8848 10232 8860
rect 10284 8888 10290 8900
rect 10888 8888 10916 8987
rect 11330 8984 11336 8996
rect 11388 9024 11394 9036
rect 11808 9033 11836 9064
rect 12066 9052 12072 9104
rect 12124 9092 12130 9104
rect 12618 9101 12624 9104
rect 12575 9095 12624 9101
rect 12575 9092 12587 9095
rect 12124 9064 12587 9092
rect 12124 9052 12130 9064
rect 12575 9061 12587 9064
rect 12621 9061 12624 9095
rect 12575 9055 12624 9061
rect 12618 9052 12624 9055
rect 12676 9052 12682 9104
rect 12728 9101 12756 9132
rect 14642 9120 14648 9132
rect 14700 9120 14706 9172
rect 16298 9120 16304 9172
rect 16356 9160 16362 9172
rect 16393 9163 16451 9169
rect 16393 9160 16405 9163
rect 16356 9132 16405 9160
rect 16356 9120 16362 9132
rect 16393 9129 16405 9132
rect 16439 9129 16451 9163
rect 16393 9123 16451 9129
rect 12713 9095 12771 9101
rect 12713 9061 12725 9095
rect 12759 9061 12771 9095
rect 12713 9055 12771 9061
rect 12802 9052 12808 9104
rect 12860 9092 12866 9104
rect 13081 9095 13139 9101
rect 12860 9064 12905 9092
rect 12860 9052 12866 9064
rect 13081 9061 13093 9095
rect 13127 9092 13139 9095
rect 14921 9095 14979 9101
rect 14921 9092 14933 9095
rect 13127 9064 14933 9092
rect 13127 9061 13139 9064
rect 13081 9055 13139 9061
rect 14921 9061 14933 9064
rect 14967 9061 14979 9095
rect 14921 9055 14979 9061
rect 15654 9052 15660 9104
rect 15712 9052 15718 9104
rect 11609 9027 11667 9033
rect 11609 9024 11621 9027
rect 11388 8996 11621 9024
rect 11388 8984 11394 8996
rect 11609 8993 11621 8996
rect 11655 8993 11667 9027
rect 11609 8987 11667 8993
rect 11793 9027 11851 9033
rect 11793 8993 11805 9027
rect 11839 8993 11851 9027
rect 11793 8987 11851 8993
rect 12897 9027 12955 9033
rect 12897 8993 12909 9027
rect 12943 8993 12955 9027
rect 13170 9024 13176 9036
rect 13131 8996 13176 9024
rect 12897 8987 12955 8993
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8956 11115 8959
rect 12437 8959 12495 8965
rect 12437 8956 12449 8959
rect 11103 8928 12449 8956
rect 11103 8925 11115 8928
rect 11057 8919 11115 8925
rect 12437 8925 12449 8928
rect 12483 8925 12495 8959
rect 12912 8956 12940 8987
rect 13170 8984 13176 8996
rect 13228 8984 13234 9036
rect 13354 9024 13360 9036
rect 13315 8996 13360 9024
rect 13354 8984 13360 8996
rect 13412 8984 13418 9036
rect 13265 8959 13323 8965
rect 13265 8956 13277 8959
rect 12912 8928 13277 8956
rect 12437 8919 12495 8925
rect 13265 8925 13277 8928
rect 13311 8925 13323 8959
rect 13265 8919 13323 8925
rect 14645 8959 14703 8965
rect 14645 8925 14657 8959
rect 14691 8956 14703 8959
rect 14918 8956 14924 8968
rect 14691 8928 14924 8956
rect 14691 8925 14703 8928
rect 14645 8919 14703 8925
rect 10284 8860 10916 8888
rect 12452 8888 12480 8919
rect 14918 8916 14924 8928
rect 14976 8916 14982 8968
rect 13630 8888 13636 8900
rect 12452 8860 13636 8888
rect 10284 8848 10290 8860
rect 13630 8848 13636 8860
rect 13688 8848 13694 8900
rect 8570 8820 8576 8832
rect 6288 8792 8576 8820
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 9674 8820 9680 8832
rect 9635 8792 9680 8820
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 1104 8730 16836 8752
rect 1104 8678 3604 8730
rect 3656 8678 3668 8730
rect 3720 8678 3732 8730
rect 3784 8678 3796 8730
rect 3848 8678 8848 8730
rect 8900 8678 8912 8730
rect 8964 8678 8976 8730
rect 9028 8678 9040 8730
rect 9092 8678 14092 8730
rect 14144 8678 14156 8730
rect 14208 8678 14220 8730
rect 14272 8678 14284 8730
rect 14336 8678 16836 8730
rect 1104 8656 16836 8678
rect 4890 8616 4896 8628
rect 4851 8588 4896 8616
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 6822 8616 6828 8628
rect 6783 8588 6828 8616
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 8478 8616 8484 8628
rect 8439 8588 8484 8616
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 9953 8619 10011 8625
rect 9953 8585 9965 8619
rect 9999 8616 10011 8619
rect 10318 8616 10324 8628
rect 9999 8588 10324 8616
rect 9999 8585 10011 8588
rect 9953 8579 10011 8585
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 7377 8551 7435 8557
rect 7377 8517 7389 8551
rect 7423 8548 7435 8551
rect 9674 8548 9680 8560
rect 7423 8520 9680 8548
rect 7423 8517 7435 8520
rect 7377 8511 7435 8517
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8480 7527 8483
rect 7834 8480 7840 8492
rect 7515 8452 7840 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 4338 8372 4344 8424
rect 4396 8412 4402 8424
rect 4801 8415 4859 8421
rect 4801 8412 4813 8415
rect 4396 8384 4813 8412
rect 4396 8372 4402 8384
rect 4801 8381 4813 8384
rect 4847 8381 4859 8415
rect 4801 8375 4859 8381
rect 6978 8415 7036 8421
rect 6978 8381 6990 8415
rect 7024 8412 7036 8415
rect 7484 8412 7512 8443
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 7024 8384 7512 8412
rect 7024 8381 7036 8384
rect 6978 8375 7036 8381
rect 7074 8347 7132 8353
rect 7074 8313 7086 8347
rect 7120 8344 7132 8347
rect 7944 8344 7972 8520
rect 9674 8508 9680 8520
rect 9732 8508 9738 8560
rect 8570 8440 8576 8492
rect 8628 8480 8634 8492
rect 10410 8480 10416 8492
rect 8628 8452 9352 8480
rect 10371 8452 10416 8480
rect 8628 8440 8634 8452
rect 8662 8412 8668 8424
rect 8623 8384 8668 8412
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 9324 8412 9352 8452
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8480 10655 8483
rect 11330 8480 11336 8492
rect 10643 8452 11336 8480
rect 10643 8449 10655 8452
rect 10597 8443 10655 8449
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 13170 8412 13176 8424
rect 9324 8384 13176 8412
rect 13170 8372 13176 8384
rect 13228 8372 13234 8424
rect 13906 8412 13912 8424
rect 13867 8384 13912 8412
rect 13906 8372 13912 8384
rect 13964 8372 13970 8424
rect 16482 8412 16488 8424
rect 16443 8384 16488 8412
rect 16482 8372 16488 8384
rect 16540 8372 16546 8424
rect 7120 8316 7972 8344
rect 7120 8313 7132 8316
rect 7074 8307 7132 8313
rect 10226 8304 10232 8356
rect 10284 8344 10290 8356
rect 10321 8347 10379 8353
rect 10321 8344 10333 8347
rect 10284 8316 10333 8344
rect 10284 8304 10290 8316
rect 10321 8313 10333 8316
rect 10367 8313 10379 8347
rect 10321 8307 10379 8313
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 14001 8279 14059 8285
rect 14001 8276 14013 8279
rect 13872 8248 14013 8276
rect 13872 8236 13878 8248
rect 14001 8245 14013 8248
rect 14047 8245 14059 8279
rect 16298 8276 16304 8288
rect 16259 8248 16304 8276
rect 14001 8239 14059 8245
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 1104 8186 16836 8208
rect 1104 8134 6226 8186
rect 6278 8134 6290 8186
rect 6342 8134 6354 8186
rect 6406 8134 6418 8186
rect 6470 8134 11470 8186
rect 11522 8134 11534 8186
rect 11586 8134 11598 8186
rect 11650 8134 11662 8186
rect 11714 8134 16836 8186
rect 1104 8112 16836 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 3142 8072 3148 8084
rect 1627 8044 3148 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 3142 8032 3148 8044
rect 3200 8032 3206 8084
rect 11330 8032 11336 8084
rect 11388 8072 11394 8084
rect 11609 8075 11667 8081
rect 11609 8072 11621 8075
rect 11388 8044 11621 8072
rect 11388 8032 11394 8044
rect 11609 8041 11621 8044
rect 11655 8041 11667 8075
rect 11609 8035 11667 8041
rect 12342 8032 12348 8084
rect 12400 8072 12406 8084
rect 13078 8072 13084 8084
rect 12400 8044 13084 8072
rect 12400 8032 12406 8044
rect 13078 8032 13084 8044
rect 13136 8072 13142 8084
rect 13722 8072 13728 8084
rect 13136 8044 13728 8072
rect 13136 8032 13142 8044
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 13906 8032 13912 8084
rect 13964 8072 13970 8084
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 13964 8044 14105 8072
rect 13964 8032 13970 8044
rect 14093 8041 14105 8044
rect 14139 8041 14151 8075
rect 14093 8035 14151 8041
rect 11238 7964 11244 8016
rect 11296 8004 11302 8016
rect 13446 8004 13452 8016
rect 11296 7976 13452 8004
rect 11296 7964 11302 7976
rect 13446 7964 13452 7976
rect 13504 8004 13510 8016
rect 13504 7976 13952 8004
rect 13504 7964 13510 7976
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 2314 7936 2320 7948
rect 2275 7908 2320 7936
rect 2314 7896 2320 7908
rect 2372 7896 2378 7948
rect 2958 7936 2964 7948
rect 2919 7908 2964 7936
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 3145 7939 3203 7945
rect 3145 7905 3157 7939
rect 3191 7936 3203 7939
rect 4154 7936 4160 7948
rect 3191 7908 4160 7936
rect 3191 7905 3203 7908
rect 3145 7899 3203 7905
rect 4154 7896 4160 7908
rect 4212 7896 4218 7948
rect 6086 7896 6092 7948
rect 6144 7936 6150 7948
rect 6641 7939 6699 7945
rect 6641 7936 6653 7939
rect 6144 7908 6653 7936
rect 6144 7896 6150 7908
rect 6641 7905 6653 7908
rect 6687 7936 6699 7939
rect 6730 7936 6736 7948
rect 6687 7908 6736 7936
rect 6687 7905 6699 7908
rect 6641 7899 6699 7905
rect 6730 7896 6736 7908
rect 6788 7936 6794 7948
rect 8662 7936 8668 7948
rect 6788 7908 8668 7936
rect 6788 7896 6794 7908
rect 8662 7896 8668 7908
rect 8720 7936 8726 7948
rect 9309 7939 9367 7945
rect 9309 7936 9321 7939
rect 8720 7908 9321 7936
rect 8720 7896 8726 7908
rect 9309 7905 9321 7908
rect 9355 7905 9367 7939
rect 9309 7899 9367 7905
rect 11793 7939 11851 7945
rect 11793 7905 11805 7939
rect 11839 7905 11851 7939
rect 11793 7899 11851 7905
rect 11808 7868 11836 7899
rect 11882 7896 11888 7948
rect 11940 7936 11946 7948
rect 12161 7939 12219 7945
rect 11940 7908 11985 7936
rect 11940 7896 11946 7908
rect 12161 7905 12173 7939
rect 12207 7936 12219 7939
rect 12618 7936 12624 7948
rect 12207 7908 12624 7936
rect 12207 7905 12219 7908
rect 12161 7899 12219 7905
rect 12618 7896 12624 7908
rect 12676 7896 12682 7948
rect 13541 7939 13599 7945
rect 13541 7905 13553 7939
rect 13587 7936 13599 7939
rect 13587 7908 13676 7936
rect 13587 7905 13599 7908
rect 13541 7899 13599 7905
rect 12526 7868 12532 7880
rect 11808 7840 12532 7868
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 12250 7760 12256 7812
rect 12308 7800 12314 7812
rect 13648 7800 13676 7908
rect 13722 7896 13728 7948
rect 13780 7936 13786 7948
rect 13924 7945 13952 7976
rect 13817 7939 13875 7945
rect 13817 7936 13829 7939
rect 13780 7908 13829 7936
rect 13780 7896 13786 7908
rect 13817 7905 13829 7908
rect 13863 7905 13875 7939
rect 13817 7899 13875 7905
rect 13909 7939 13967 7945
rect 13909 7905 13921 7939
rect 13955 7905 13967 7939
rect 13909 7899 13967 7905
rect 14369 7939 14427 7945
rect 14369 7905 14381 7939
rect 14415 7905 14427 7939
rect 14369 7899 14427 7905
rect 13832 7868 13860 7899
rect 14384 7868 14412 7899
rect 14550 7896 14556 7948
rect 14608 7936 14614 7948
rect 14645 7939 14703 7945
rect 14645 7936 14657 7939
rect 14608 7908 14657 7936
rect 14608 7896 14614 7908
rect 14645 7905 14657 7908
rect 14691 7936 14703 7939
rect 15010 7936 15016 7948
rect 14691 7908 15016 7936
rect 14691 7905 14703 7908
rect 14645 7899 14703 7905
rect 15010 7896 15016 7908
rect 15068 7896 15074 7948
rect 15654 7936 15660 7948
rect 15615 7908 15660 7936
rect 15654 7896 15660 7908
rect 15712 7896 15718 7948
rect 13832 7840 14412 7868
rect 14826 7828 14832 7880
rect 14884 7828 14890 7880
rect 14844 7800 14872 7828
rect 16390 7800 16396 7812
rect 12308 7772 12664 7800
rect 13648 7772 16396 7800
rect 12308 7760 12314 7772
rect 2406 7692 2412 7744
rect 2464 7732 2470 7744
rect 2501 7735 2559 7741
rect 2501 7732 2513 7735
rect 2464 7704 2513 7732
rect 2464 7692 2470 7704
rect 2501 7701 2513 7704
rect 2547 7701 2559 7735
rect 2501 7695 2559 7701
rect 2682 7692 2688 7744
rect 2740 7732 2746 7744
rect 2777 7735 2835 7741
rect 2777 7732 2789 7735
rect 2740 7704 2789 7732
rect 2740 7692 2746 7704
rect 2777 7701 2789 7704
rect 2823 7701 2835 7735
rect 6822 7732 6828 7744
rect 6783 7704 6828 7732
rect 2777 7695 2835 7701
rect 6822 7692 6828 7704
rect 6880 7692 6886 7744
rect 9125 7735 9183 7741
rect 9125 7701 9137 7735
rect 9171 7732 9183 7735
rect 9214 7732 9220 7744
rect 9171 7704 9220 7732
rect 9171 7701 9183 7704
rect 9125 7695 9183 7701
rect 9214 7692 9220 7704
rect 9272 7692 9278 7744
rect 12069 7735 12127 7741
rect 12069 7701 12081 7735
rect 12115 7732 12127 7735
rect 12342 7732 12348 7744
rect 12115 7704 12348 7732
rect 12115 7701 12127 7704
rect 12069 7695 12127 7701
rect 12342 7692 12348 7704
rect 12400 7692 12406 7744
rect 12636 7732 12664 7772
rect 16390 7760 16396 7772
rect 16448 7760 16454 7812
rect 13633 7735 13691 7741
rect 13633 7732 13645 7735
rect 12636 7704 13645 7732
rect 13633 7701 13645 7704
rect 13679 7732 13691 7735
rect 14461 7735 14519 7741
rect 14461 7732 14473 7735
rect 13679 7704 14473 7732
rect 13679 7701 13691 7704
rect 13633 7695 13691 7701
rect 14461 7701 14473 7704
rect 14507 7701 14519 7735
rect 14461 7695 14519 7701
rect 14550 7692 14556 7744
rect 14608 7732 14614 7744
rect 14737 7735 14795 7741
rect 14737 7732 14749 7735
rect 14608 7704 14749 7732
rect 14608 7692 14614 7704
rect 14737 7701 14749 7704
rect 14783 7701 14795 7735
rect 14737 7695 14795 7701
rect 14826 7692 14832 7744
rect 14884 7732 14890 7744
rect 15102 7732 15108 7744
rect 14884 7704 15108 7732
rect 14884 7692 14890 7704
rect 15102 7692 15108 7704
rect 15160 7692 15166 7744
rect 15841 7735 15899 7741
rect 15841 7701 15853 7735
rect 15887 7732 15899 7735
rect 15930 7732 15936 7744
rect 15887 7704 15936 7732
rect 15887 7701 15899 7704
rect 15841 7695 15899 7701
rect 15930 7692 15936 7704
rect 15988 7692 15994 7744
rect 1104 7642 16836 7664
rect 1104 7590 3604 7642
rect 3656 7590 3668 7642
rect 3720 7590 3732 7642
rect 3784 7590 3796 7642
rect 3848 7590 8848 7642
rect 8900 7590 8912 7642
rect 8964 7590 8976 7642
rect 9028 7590 9040 7642
rect 9092 7590 14092 7642
rect 14144 7590 14156 7642
rect 14208 7590 14220 7642
rect 14272 7590 14284 7642
rect 14336 7590 16836 7642
rect 1104 7568 16836 7590
rect 3418 7488 3424 7540
rect 3476 7528 3482 7540
rect 4430 7528 4436 7540
rect 3476 7500 4436 7528
rect 3476 7488 3482 7500
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 11882 7528 11888 7540
rect 11843 7500 11888 7528
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 11974 7488 11980 7540
rect 12032 7528 12038 7540
rect 12526 7528 12532 7540
rect 12032 7500 12388 7528
rect 12487 7500 12532 7528
rect 12032 7488 12038 7500
rect 3712 7432 4936 7460
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 2682 7392 2688 7404
rect 1719 7364 2688 7392
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 2958 7352 2964 7404
rect 3016 7392 3022 7404
rect 3145 7395 3203 7401
rect 3145 7392 3157 7395
rect 3016 7364 3157 7392
rect 3016 7352 3022 7364
rect 3145 7361 3157 7364
rect 3191 7392 3203 7395
rect 3712 7392 3740 7432
rect 4525 7395 4583 7401
rect 4525 7392 4537 7395
rect 3191 7364 3740 7392
rect 3191 7361 3203 7364
rect 3145 7355 3203 7361
rect 1394 7324 1400 7336
rect 1355 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7284 1458 7336
rect 3418 7324 3424 7336
rect 3379 7296 3424 7324
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 3605 7327 3663 7333
rect 3605 7293 3617 7327
rect 3651 7324 3663 7327
rect 3712 7324 3740 7364
rect 4172 7364 4537 7392
rect 3651 7296 3740 7324
rect 3789 7327 3847 7333
rect 3651 7293 3663 7296
rect 3605 7287 3663 7293
rect 3789 7293 3801 7327
rect 3835 7324 3847 7327
rect 4062 7324 4068 7336
rect 3835 7296 4068 7324
rect 3835 7293 3847 7296
rect 3789 7287 3847 7293
rect 4062 7284 4068 7296
rect 4120 7284 4126 7336
rect 2406 7216 2412 7268
rect 2464 7216 2470 7268
rect 3510 7256 3516 7268
rect 3471 7228 3516 7256
rect 3510 7216 3516 7228
rect 3568 7216 3574 7268
rect 4172 7265 4200 7364
rect 4525 7361 4537 7364
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 4430 7324 4436 7336
rect 4391 7296 4436 7324
rect 4430 7284 4436 7296
rect 4488 7284 4494 7336
rect 4908 7333 4936 7432
rect 7926 7420 7932 7472
rect 7984 7460 7990 7472
rect 8205 7463 8263 7469
rect 8205 7460 8217 7463
rect 7984 7432 8217 7460
rect 7984 7420 7990 7432
rect 8205 7429 8217 7432
rect 8251 7429 8263 7463
rect 8205 7423 8263 7429
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7392 5135 7395
rect 9766 7392 9772 7404
rect 5123 7364 9772 7392
rect 5123 7361 5135 7364
rect 5077 7355 5135 7361
rect 9766 7352 9772 7364
rect 9824 7352 9830 7404
rect 12250 7392 12256 7404
rect 12084 7364 12256 7392
rect 4893 7327 4951 7333
rect 4893 7293 4905 7327
rect 4939 7293 4951 7327
rect 4893 7287 4951 7293
rect 5353 7327 5411 7333
rect 5353 7293 5365 7327
rect 5399 7324 5411 7327
rect 6086 7324 6092 7336
rect 5399 7296 6092 7324
rect 5399 7293 5411 7296
rect 5353 7287 5411 7293
rect 6086 7284 6092 7296
rect 6144 7284 6150 7336
rect 6457 7327 6515 7333
rect 6457 7293 6469 7327
rect 6503 7293 6515 7327
rect 6457 7287 6515 7293
rect 10137 7327 10195 7333
rect 10137 7293 10149 7327
rect 10183 7324 10195 7327
rect 10226 7324 10232 7336
rect 10183 7296 10232 7324
rect 10183 7293 10195 7296
rect 10137 7287 10195 7293
rect 4157 7259 4215 7265
rect 4157 7256 4169 7259
rect 3804 7228 4169 7256
rect 3234 7148 3240 7200
rect 3292 7188 3298 7200
rect 3528 7188 3556 7216
rect 3804 7188 3832 7228
rect 4157 7225 4169 7228
rect 4203 7225 4215 7259
rect 4157 7219 4215 7225
rect 4249 7259 4307 7265
rect 4249 7225 4261 7259
rect 4295 7256 4307 7259
rect 4801 7259 4859 7265
rect 4801 7256 4813 7259
rect 4295 7228 4813 7256
rect 4295 7225 4307 7228
rect 4249 7219 4307 7225
rect 4801 7225 4813 7228
rect 4847 7256 4859 7259
rect 5718 7256 5724 7268
rect 4847 7228 5724 7256
rect 4847 7225 4859 7228
rect 4801 7219 4859 7225
rect 5718 7216 5724 7228
rect 5776 7216 5782 7268
rect 3292 7160 3337 7188
rect 3528 7160 3832 7188
rect 3881 7191 3939 7197
rect 3292 7148 3298 7160
rect 3881 7157 3893 7191
rect 3927 7188 3939 7191
rect 4338 7188 4344 7200
rect 3927 7160 4344 7188
rect 3927 7157 3939 7160
rect 3881 7151 3939 7157
rect 4338 7148 4344 7160
rect 4396 7148 4402 7200
rect 4706 7188 4712 7200
rect 4667 7160 4712 7188
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 5169 7191 5227 7197
rect 5169 7157 5181 7191
rect 5215 7188 5227 7191
rect 5258 7188 5264 7200
rect 5215 7160 5264 7188
rect 5215 7157 5227 7160
rect 5169 7151 5227 7157
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 6472 7188 6500 7287
rect 10226 7284 10232 7296
rect 10284 7284 10290 7336
rect 10778 7324 10784 7336
rect 10739 7296 10784 7324
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 10962 7324 10968 7336
rect 10923 7296 10968 7324
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11238 7324 11244 7336
rect 11199 7296 11244 7324
rect 11238 7284 11244 7296
rect 11296 7284 11302 7336
rect 12084 7333 12112 7364
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 12360 7392 12388 7500
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 13446 7488 13452 7540
rect 13504 7528 13510 7540
rect 14461 7531 14519 7537
rect 13504 7500 14412 7528
rect 13504 7488 13510 7500
rect 14185 7463 14243 7469
rect 14185 7429 14197 7463
rect 14231 7460 14243 7463
rect 14384 7460 14412 7500
rect 14461 7497 14473 7531
rect 14507 7528 14519 7531
rect 14642 7528 14648 7540
rect 14507 7500 14648 7528
rect 14507 7497 14519 7500
rect 14461 7491 14519 7497
rect 14642 7488 14648 7500
rect 14700 7488 14706 7540
rect 16390 7528 16396 7540
rect 16351 7500 16396 7528
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 14231 7432 14320 7460
rect 14384 7432 14596 7460
rect 14231 7429 14243 7432
rect 14185 7423 14243 7429
rect 12360 7364 12572 7392
rect 11425 7327 11483 7333
rect 11425 7293 11437 7327
rect 11471 7324 11483 7327
rect 12069 7327 12127 7333
rect 12069 7324 12081 7327
rect 11471 7296 12081 7324
rect 11471 7293 11483 7296
rect 11425 7287 11483 7293
rect 12069 7293 12081 7296
rect 12115 7293 12127 7327
rect 12069 7287 12127 7293
rect 12342 7284 12348 7336
rect 12400 7324 12406 7336
rect 12544 7333 12572 7364
rect 13814 7352 13820 7404
rect 13872 7352 13878 7404
rect 13906 7352 13912 7404
rect 13964 7352 13970 7404
rect 14292 7401 14320 7432
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 12400 7296 12449 7324
rect 12400 7284 12406 7296
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 12437 7287 12495 7293
rect 12529 7327 12587 7333
rect 12529 7293 12541 7327
rect 12575 7293 12587 7327
rect 12529 7287 12587 7293
rect 12618 7284 12624 7336
rect 12676 7324 12682 7336
rect 13538 7324 13544 7336
rect 12676 7296 12769 7324
rect 13499 7296 13544 7324
rect 12676 7284 12682 7296
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 13689 7327 13747 7333
rect 13689 7293 13701 7327
rect 13735 7324 13747 7327
rect 13832 7324 13860 7352
rect 13735 7296 13860 7324
rect 13924 7324 13952 7352
rect 14006 7327 14064 7333
rect 14006 7324 14018 7327
rect 13924 7296 14018 7324
rect 13735 7293 13747 7296
rect 13689 7287 13747 7293
rect 14006 7293 14018 7296
rect 14052 7293 14064 7327
rect 14366 7324 14372 7336
rect 14006 7287 14064 7293
rect 14200 7296 14372 7324
rect 6730 7256 6736 7268
rect 6691 7228 6736 7256
rect 6730 7216 6736 7228
rect 6788 7216 6794 7268
rect 6822 7216 6828 7268
rect 6880 7256 6886 7268
rect 6880 7228 7222 7256
rect 6880 7216 6886 7228
rect 9214 7216 9220 7268
rect 9272 7216 9278 7268
rect 9858 7256 9864 7268
rect 9819 7228 9864 7256
rect 9858 7216 9864 7228
rect 9916 7216 9922 7268
rect 10318 7256 10324 7268
rect 10279 7228 10324 7256
rect 10318 7216 10324 7228
rect 10376 7216 10382 7268
rect 11974 7216 11980 7268
rect 12032 7256 12038 7268
rect 12161 7259 12219 7265
rect 12161 7256 12173 7259
rect 12032 7228 12173 7256
rect 12032 7216 12038 7228
rect 12161 7225 12173 7228
rect 12207 7225 12219 7259
rect 12161 7219 12219 7225
rect 12253 7259 12311 7265
rect 12253 7225 12265 7259
rect 12299 7256 12311 7259
rect 12636 7256 12664 7284
rect 12299 7228 12664 7256
rect 13817 7259 13875 7265
rect 12299 7225 12311 7228
rect 12253 7219 12311 7225
rect 7098 7188 7104 7200
rect 6472 7160 7104 7188
rect 7098 7148 7104 7160
rect 7156 7188 7162 7200
rect 7466 7188 7472 7200
rect 7156 7160 7472 7188
rect 7156 7148 7162 7160
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 8202 7148 8208 7200
rect 8260 7188 8266 7200
rect 8389 7191 8447 7197
rect 8389 7188 8401 7191
rect 8260 7160 8401 7188
rect 8260 7148 8266 7160
rect 8389 7157 8401 7160
rect 8435 7157 8447 7191
rect 12360 7188 12388 7228
rect 13817 7225 13829 7259
rect 13863 7225 13875 7259
rect 13817 7219 13875 7225
rect 13909 7259 13967 7265
rect 13909 7225 13921 7259
rect 13955 7256 13967 7259
rect 14200 7256 14228 7296
rect 14366 7284 14372 7296
rect 14424 7284 14430 7336
rect 14568 7333 14596 7432
rect 14645 7395 14703 7401
rect 14645 7361 14657 7395
rect 14691 7392 14703 7395
rect 14918 7392 14924 7404
rect 14691 7364 14924 7392
rect 14691 7361 14703 7364
rect 14645 7355 14703 7361
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 14553 7327 14611 7333
rect 14553 7293 14565 7327
rect 14599 7293 14611 7327
rect 14553 7287 14611 7293
rect 13955 7228 14228 7256
rect 14277 7259 14335 7265
rect 13955 7225 13967 7228
rect 13909 7219 13967 7225
rect 14277 7225 14289 7259
rect 14323 7256 14335 7259
rect 14921 7259 14979 7265
rect 14921 7256 14933 7259
rect 14323 7228 14933 7256
rect 14323 7225 14335 7228
rect 14277 7219 14335 7225
rect 14921 7225 14933 7228
rect 14967 7225 14979 7259
rect 14921 7219 14979 7225
rect 12434 7188 12440 7200
rect 12360 7160 12440 7188
rect 8389 7151 8447 7157
rect 12434 7148 12440 7160
rect 12492 7148 12498 7200
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13832 7188 13860 7219
rect 15930 7216 15936 7268
rect 15988 7216 15994 7268
rect 15010 7188 15016 7200
rect 13832 7160 15016 7188
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 1104 7098 16836 7120
rect 1104 7046 6226 7098
rect 6278 7046 6290 7098
rect 6342 7046 6354 7098
rect 6406 7046 6418 7098
rect 6470 7046 11470 7098
rect 11522 7046 11534 7098
rect 11586 7046 11598 7098
rect 11650 7046 11662 7098
rect 11714 7046 16836 7098
rect 1104 7024 16836 7046
rect 3237 6987 3295 6993
rect 3237 6953 3249 6987
rect 3283 6984 3295 6987
rect 3510 6984 3516 6996
rect 3283 6956 3516 6984
rect 3283 6953 3295 6956
rect 3237 6947 3295 6953
rect 3510 6944 3516 6956
rect 3568 6944 3574 6996
rect 5718 6984 5724 6996
rect 5679 6956 5724 6984
rect 5718 6944 5724 6956
rect 5776 6944 5782 6996
rect 8202 6984 8208 6996
rect 8036 6956 8208 6984
rect 2498 6876 2504 6928
rect 2556 6876 2562 6928
rect 5258 6876 5264 6928
rect 5316 6876 5322 6928
rect 6457 6919 6515 6925
rect 6457 6885 6469 6919
rect 6503 6916 6515 6919
rect 6638 6916 6644 6928
rect 6503 6888 6644 6916
rect 6503 6885 6515 6888
rect 6457 6879 6515 6885
rect 6638 6876 6644 6888
rect 6696 6876 6702 6928
rect 7926 6916 7932 6928
rect 7887 6888 7932 6916
rect 7926 6876 7932 6888
rect 7984 6876 7990 6928
rect 8036 6925 8064 6956
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 13538 6984 13544 6996
rect 11624 6956 13544 6984
rect 8021 6919 8079 6925
rect 8021 6885 8033 6919
rect 8067 6885 8079 6919
rect 8021 6879 8079 6885
rect 6273 6851 6331 6857
rect 6273 6817 6285 6851
rect 6319 6817 6331 6851
rect 6273 6811 6331 6817
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 6914 6848 6920 6860
rect 6595 6820 6920 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 1394 6740 1400 6792
rect 1452 6780 1458 6792
rect 1489 6783 1547 6789
rect 1489 6780 1501 6783
rect 1452 6752 1501 6780
rect 1452 6740 1458 6752
rect 1489 6749 1501 6752
rect 1535 6749 1547 6783
rect 1489 6743 1547 6749
rect 1765 6783 1823 6789
rect 1765 6749 1777 6783
rect 1811 6780 1823 6783
rect 3234 6780 3240 6792
rect 1811 6752 3240 6780
rect 1811 6749 1823 6752
rect 1765 6743 1823 6749
rect 1504 6656 1532 6743
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6780 4031 6783
rect 4249 6783 4307 6789
rect 4019 6752 4108 6780
rect 4019 6749 4031 6752
rect 3973 6743 4031 6749
rect 2774 6672 2780 6724
rect 2832 6672 2838 6724
rect 1486 6644 1492 6656
rect 1399 6616 1492 6644
rect 1486 6604 1492 6616
rect 1544 6644 1550 6656
rect 2792 6644 2820 6672
rect 4080 6644 4108 6752
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 4338 6780 4344 6792
rect 4295 6752 4344 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 4338 6740 4344 6752
rect 4396 6740 4402 6792
rect 4706 6740 4712 6792
rect 4764 6780 4770 6792
rect 5258 6780 5264 6792
rect 4764 6752 5264 6780
rect 4764 6740 4770 6752
rect 5258 6740 5264 6752
rect 5316 6780 5322 6792
rect 6288 6780 6316 6811
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 7745 6851 7803 6857
rect 7745 6817 7757 6851
rect 7791 6817 7803 6851
rect 8137 6851 8195 6857
rect 8137 6848 8149 6851
rect 7745 6811 7803 6817
rect 8128 6817 8149 6848
rect 8183 6817 8195 6851
rect 8128 6811 8195 6817
rect 7760 6780 7788 6811
rect 5316 6752 7788 6780
rect 5316 6740 5322 6752
rect 6273 6715 6331 6721
rect 6273 6681 6285 6715
rect 6319 6712 6331 6715
rect 6730 6712 6736 6724
rect 6319 6684 6736 6712
rect 6319 6681 6331 6684
rect 6273 6675 6331 6681
rect 6730 6672 6736 6684
rect 6788 6672 6794 6724
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 8128 6712 8156 6811
rect 10318 6808 10324 6860
rect 10376 6848 10382 6860
rect 10413 6851 10471 6857
rect 10413 6848 10425 6851
rect 10376 6820 10425 6848
rect 10376 6808 10382 6820
rect 10413 6817 10425 6820
rect 10459 6817 10471 6851
rect 10413 6811 10471 6817
rect 10505 6851 10563 6857
rect 10505 6817 10517 6851
rect 10551 6848 10563 6851
rect 11333 6851 11391 6857
rect 11333 6848 11345 6851
rect 10551 6820 11345 6848
rect 10551 6817 10563 6820
rect 10505 6811 10563 6817
rect 11333 6817 11345 6820
rect 11379 6848 11391 6851
rect 11624 6848 11652 6956
rect 13538 6944 13544 6956
rect 13596 6944 13602 6996
rect 12434 6916 12440 6928
rect 11716 6888 12440 6916
rect 11716 6857 11744 6888
rect 12434 6876 12440 6888
rect 12492 6916 12498 6928
rect 12621 6919 12679 6925
rect 12621 6916 12633 6919
rect 12492 6888 12633 6916
rect 12492 6876 12498 6888
rect 12621 6885 12633 6888
rect 12667 6885 12679 6919
rect 13556 6916 13584 6944
rect 13556 6888 13860 6916
rect 12621 6879 12679 6885
rect 11379 6820 11652 6848
rect 11701 6851 11759 6857
rect 11379 6817 11391 6820
rect 11333 6811 11391 6817
rect 11701 6817 11713 6851
rect 11747 6817 11759 6851
rect 11701 6811 11759 6817
rect 10428 6780 10456 6811
rect 11882 6808 11888 6860
rect 11940 6848 11946 6860
rect 12069 6851 12127 6857
rect 12069 6848 12081 6851
rect 11940 6820 12081 6848
rect 11940 6808 11946 6820
rect 12069 6817 12081 6820
rect 12115 6848 12127 6851
rect 12345 6851 12403 6857
rect 12345 6848 12357 6851
rect 12115 6820 12357 6848
rect 12115 6817 12127 6820
rect 12069 6811 12127 6817
rect 12345 6817 12357 6820
rect 12391 6817 12403 6851
rect 12345 6811 12403 6817
rect 12713 6851 12771 6857
rect 12713 6817 12725 6851
rect 12759 6848 12771 6851
rect 12894 6848 12900 6860
rect 12759 6820 12900 6848
rect 12759 6817 12771 6820
rect 12713 6811 12771 6817
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 13354 6808 13360 6860
rect 13412 6848 13418 6860
rect 13832 6857 13860 6888
rect 13725 6851 13783 6857
rect 13725 6848 13737 6851
rect 13412 6820 13737 6848
rect 13412 6808 13418 6820
rect 13725 6817 13737 6820
rect 13771 6817 13783 6851
rect 13725 6811 13783 6817
rect 13817 6851 13875 6857
rect 13817 6817 13829 6851
rect 13863 6817 13875 6851
rect 14093 6851 14151 6857
rect 14093 6848 14105 6851
rect 13817 6811 13875 6817
rect 13924 6820 14105 6848
rect 11517 6783 11575 6789
rect 10428 6752 10548 6780
rect 7248 6684 8156 6712
rect 8297 6715 8355 6721
rect 7248 6672 7254 6684
rect 8297 6681 8309 6715
rect 8343 6712 8355 6715
rect 9858 6712 9864 6724
rect 8343 6684 9864 6712
rect 8343 6681 8355 6684
rect 8297 6675 8355 6681
rect 9858 6672 9864 6684
rect 9916 6672 9922 6724
rect 7466 6644 7472 6656
rect 1544 6616 7472 6644
rect 1544 6604 1550 6616
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 10520 6644 10548 6752
rect 11517 6749 11529 6783
rect 11563 6780 11575 6783
rect 11977 6783 12035 6789
rect 11563 6752 11836 6780
rect 11563 6749 11575 6752
rect 11517 6743 11575 6749
rect 11808 6721 11836 6752
rect 11977 6749 11989 6783
rect 12023 6780 12035 6783
rect 12437 6783 12495 6789
rect 12437 6780 12449 6783
rect 12023 6752 12449 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 12437 6749 12449 6752
rect 12483 6780 12495 6783
rect 12526 6780 12532 6792
rect 12483 6752 12532 6780
rect 12483 6749 12495 6752
rect 12437 6743 12495 6749
rect 12526 6740 12532 6752
rect 12584 6740 12590 6792
rect 13446 6740 13452 6792
rect 13504 6780 13510 6792
rect 13924 6780 13952 6820
rect 14093 6817 14105 6820
rect 14139 6848 14151 6851
rect 15286 6848 15292 6860
rect 14139 6820 15292 6848
rect 14139 6817 14151 6820
rect 14093 6811 14151 6817
rect 15286 6808 15292 6820
rect 15344 6808 15350 6860
rect 13504 6752 13952 6780
rect 14001 6783 14059 6789
rect 13504 6740 13510 6752
rect 14001 6749 14013 6783
rect 14047 6780 14059 6783
rect 14642 6780 14648 6792
rect 14047 6752 14648 6780
rect 14047 6749 14059 6752
rect 14001 6743 14059 6749
rect 11403 6715 11461 6721
rect 11403 6681 11415 6715
rect 11449 6712 11461 6715
rect 11793 6715 11851 6721
rect 11449 6684 11744 6712
rect 11449 6681 11461 6684
rect 11403 6675 11461 6681
rect 11514 6644 11520 6656
rect 10520 6616 11520 6644
rect 11514 6604 11520 6616
rect 11572 6644 11578 6656
rect 11609 6647 11667 6653
rect 11609 6644 11621 6647
rect 11572 6616 11621 6644
rect 11572 6604 11578 6616
rect 11609 6613 11621 6616
rect 11655 6613 11667 6647
rect 11716 6644 11744 6684
rect 11793 6681 11805 6715
rect 11839 6681 11851 6715
rect 11793 6675 11851 6681
rect 11882 6672 11888 6724
rect 11940 6712 11946 6724
rect 14016 6712 14044 6743
rect 14642 6740 14648 6752
rect 14700 6740 14706 6792
rect 11940 6684 14044 6712
rect 11940 6672 11946 6684
rect 12250 6644 12256 6656
rect 11716 6616 12256 6644
rect 11609 6607 11667 6613
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 13541 6647 13599 6653
rect 13541 6613 13553 6647
rect 13587 6644 13599 6647
rect 13814 6644 13820 6656
rect 13587 6616 13820 6644
rect 13587 6613 13599 6616
rect 13541 6607 13599 6613
rect 13814 6604 13820 6616
rect 13872 6604 13878 6656
rect 1104 6554 16836 6576
rect 1104 6502 3604 6554
rect 3656 6502 3668 6554
rect 3720 6502 3732 6554
rect 3784 6502 3796 6554
rect 3848 6502 8848 6554
rect 8900 6502 8912 6554
rect 8964 6502 8976 6554
rect 9028 6502 9040 6554
rect 9092 6502 14092 6554
rect 14144 6502 14156 6554
rect 14208 6502 14220 6554
rect 14272 6502 14284 6554
rect 14336 6502 16836 6554
rect 1104 6480 16836 6502
rect 2498 6440 2504 6452
rect 2459 6412 2504 6440
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 10689 6443 10747 6449
rect 10689 6409 10701 6443
rect 10735 6440 10747 6443
rect 10778 6440 10784 6452
rect 10735 6412 10784 6440
rect 10735 6409 10747 6412
rect 10689 6403 10747 6409
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 12069 6443 12127 6449
rect 12069 6409 12081 6443
rect 12115 6440 12127 6443
rect 12115 6412 12480 6440
rect 12115 6409 12127 6412
rect 12069 6403 12127 6409
rect 8202 6332 8208 6384
rect 8260 6372 8266 6384
rect 11701 6375 11759 6381
rect 11701 6372 11713 6375
rect 8260 6344 8800 6372
rect 8260 6332 8266 6344
rect 7852 6276 8340 6304
rect 7852 6248 7880 6276
rect 2317 6239 2375 6245
rect 2317 6205 2329 6239
rect 2363 6236 2375 6239
rect 2590 6236 2596 6248
rect 2363 6208 2596 6236
rect 2363 6205 2375 6208
rect 2317 6199 2375 6205
rect 2590 6196 2596 6208
rect 2648 6196 2654 6248
rect 3418 6196 3424 6248
rect 3476 6236 3482 6248
rect 4062 6236 4068 6248
rect 3476 6208 4068 6236
rect 3476 6196 3482 6208
rect 4062 6196 4068 6208
rect 4120 6236 4126 6248
rect 5169 6239 5227 6245
rect 5169 6236 5181 6239
rect 4120 6208 5181 6236
rect 4120 6196 4126 6208
rect 5169 6205 5181 6208
rect 5215 6205 5227 6239
rect 5169 6199 5227 6205
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6236 6883 6239
rect 7006 6236 7012 6248
rect 6871 6208 7012 6236
rect 6871 6205 6883 6208
rect 6825 6199 6883 6205
rect 5184 6168 5212 6199
rect 7006 6196 7012 6208
rect 7064 6236 7070 6248
rect 7834 6236 7840 6248
rect 7064 6208 7840 6236
rect 7064 6196 7070 6208
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 8202 6236 8208 6248
rect 8163 6208 8208 6236
rect 8202 6196 8208 6208
rect 8260 6196 8266 6248
rect 8312 6245 8340 6276
rect 8772 6245 8800 6344
rect 10244 6344 11713 6372
rect 10244 6313 10272 6344
rect 11701 6341 11713 6344
rect 11747 6341 11759 6375
rect 12452 6372 12480 6412
rect 12526 6400 12532 6452
rect 12584 6440 12590 6452
rect 13354 6440 13360 6452
rect 12584 6412 13360 6440
rect 12584 6400 12590 6412
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 15286 6440 15292 6452
rect 15247 6412 15292 6440
rect 15286 6400 15292 6412
rect 15344 6400 15350 6452
rect 15746 6400 15752 6452
rect 15804 6440 15810 6452
rect 16301 6443 16359 6449
rect 16301 6440 16313 6443
rect 15804 6412 16313 6440
rect 15804 6400 15810 6412
rect 16301 6409 16313 6412
rect 16347 6409 16359 6443
rect 16301 6403 16359 6409
rect 13446 6372 13452 6384
rect 12452 6344 13452 6372
rect 11701 6335 11759 6341
rect 13446 6332 13452 6344
rect 13504 6332 13510 6384
rect 10229 6307 10287 6313
rect 10229 6273 10241 6307
rect 10275 6273 10287 6307
rect 11974 6304 11980 6316
rect 11887 6276 11980 6304
rect 10229 6267 10287 6273
rect 11974 6264 11980 6276
rect 12032 6304 12038 6316
rect 12894 6304 12900 6316
rect 12032 6276 12900 6304
rect 12032 6264 12038 6276
rect 12894 6264 12900 6276
rect 12952 6264 12958 6316
rect 13814 6304 13820 6316
rect 13775 6276 13820 6304
rect 13814 6264 13820 6276
rect 13872 6264 13878 6316
rect 14458 6264 14464 6316
rect 14516 6304 14522 6316
rect 15654 6304 15660 6316
rect 14516 6276 15660 6304
rect 14516 6264 14522 6276
rect 15654 6264 15660 6276
rect 15712 6304 15718 6316
rect 15712 6276 15792 6304
rect 15712 6264 15718 6276
rect 8297 6239 8355 6245
rect 8297 6205 8309 6239
rect 8343 6205 8355 6239
rect 8297 6199 8355 6205
rect 8573 6239 8631 6245
rect 8573 6205 8585 6239
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 8757 6239 8815 6245
rect 8757 6205 8769 6239
rect 8803 6205 8815 6239
rect 8757 6199 8815 6205
rect 7190 6168 7196 6180
rect 5184 6140 7196 6168
rect 7190 6128 7196 6140
rect 7248 6128 7254 6180
rect 8386 6128 8392 6180
rect 8444 6168 8450 6180
rect 8588 6168 8616 6199
rect 9766 6196 9772 6248
rect 9824 6236 9830 6248
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 9824 6208 9965 6236
rect 9824 6196 9830 6208
rect 9953 6205 9965 6208
rect 9999 6205 10011 6239
rect 9953 6199 10011 6205
rect 10137 6239 10195 6245
rect 10137 6205 10149 6239
rect 10183 6205 10195 6239
rect 10318 6236 10324 6248
rect 10279 6208 10324 6236
rect 10137 6199 10195 6205
rect 8444 6140 8489 6168
rect 8588 6140 8892 6168
rect 8444 6128 8450 6140
rect 8864 6112 8892 6140
rect 5258 6100 5264 6112
rect 5219 6072 5264 6100
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 6638 6060 6644 6112
rect 6696 6100 6702 6112
rect 6917 6103 6975 6109
rect 6917 6100 6929 6103
rect 6696 6072 6929 6100
rect 6696 6060 6702 6072
rect 6917 6069 6929 6072
rect 6963 6100 6975 6103
rect 7558 6100 7564 6112
rect 6963 6072 7564 6100
rect 6963 6069 6975 6072
rect 6917 6063 6975 6069
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 8021 6103 8079 6109
rect 8021 6069 8033 6103
rect 8067 6100 8079 6103
rect 8478 6100 8484 6112
rect 8067 6072 8484 6100
rect 8067 6069 8079 6072
rect 8021 6063 8079 6069
rect 8478 6060 8484 6072
rect 8536 6060 8542 6112
rect 8846 6100 8852 6112
rect 8807 6072 8852 6100
rect 8846 6060 8852 6072
rect 8904 6060 8910 6112
rect 10152 6100 10180 6199
rect 10318 6196 10324 6208
rect 10376 6196 10382 6248
rect 10502 6236 10508 6248
rect 10463 6208 10508 6236
rect 10502 6196 10508 6208
rect 10560 6236 10566 6248
rect 10781 6239 10839 6245
rect 10781 6236 10793 6239
rect 10560 6208 10793 6236
rect 10560 6196 10566 6208
rect 10781 6205 10793 6208
rect 10827 6205 10839 6239
rect 10962 6236 10968 6248
rect 10923 6208 10968 6236
rect 10781 6199 10839 6205
rect 10962 6196 10968 6208
rect 11020 6196 11026 6248
rect 12069 6239 12127 6245
rect 12069 6205 12081 6239
rect 12115 6236 12127 6239
rect 12158 6236 12164 6248
rect 12115 6208 12164 6236
rect 12115 6205 12127 6208
rect 12069 6199 12127 6205
rect 12158 6196 12164 6208
rect 12216 6196 12222 6248
rect 13446 6236 13452 6248
rect 13407 6208 13452 6236
rect 13446 6196 13452 6208
rect 13504 6196 13510 6248
rect 15764 6245 15792 6276
rect 13541 6239 13599 6245
rect 13541 6205 13553 6239
rect 13587 6205 13599 6239
rect 13541 6199 13599 6205
rect 15749 6239 15807 6245
rect 15749 6205 15761 6239
rect 15795 6205 15807 6239
rect 16482 6236 16488 6248
rect 16443 6208 16488 6236
rect 15749 6199 15807 6205
rect 11057 6103 11115 6109
rect 11057 6100 11069 6103
rect 10152 6072 11069 6100
rect 11057 6069 11069 6072
rect 11103 6100 11115 6103
rect 12342 6100 12348 6112
rect 11103 6072 12348 6100
rect 11103 6069 11115 6072
rect 11057 6063 11115 6069
rect 12342 6060 12348 6072
rect 12400 6060 12406 6112
rect 13556 6100 13584 6199
rect 16482 6196 16488 6208
rect 16540 6196 16546 6248
rect 14550 6128 14556 6180
rect 14608 6128 14614 6180
rect 13814 6100 13820 6112
rect 13556 6072 13820 6100
rect 13814 6060 13820 6072
rect 13872 6100 13878 6112
rect 14826 6100 14832 6112
rect 13872 6072 14832 6100
rect 13872 6060 13878 6072
rect 14826 6060 14832 6072
rect 14884 6060 14890 6112
rect 15930 6100 15936 6112
rect 15891 6072 15936 6100
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 1104 6010 16836 6032
rect 1104 5958 6226 6010
rect 6278 5958 6290 6010
rect 6342 5958 6354 6010
rect 6406 5958 6418 6010
rect 6470 5958 11470 6010
rect 11522 5958 11534 6010
rect 11586 5958 11598 6010
rect 11650 5958 11662 6010
rect 11714 5958 16836 6010
rect 1104 5936 16836 5958
rect 1578 5896 1584 5908
rect 1539 5868 1584 5896
rect 1578 5856 1584 5868
rect 1636 5856 1642 5908
rect 3881 5899 3939 5905
rect 3881 5865 3893 5899
rect 3927 5896 3939 5899
rect 4154 5896 4160 5908
rect 3927 5868 4160 5896
rect 3927 5865 3939 5868
rect 3881 5859 3939 5865
rect 4154 5856 4160 5868
rect 4212 5896 4218 5908
rect 5258 5896 5264 5908
rect 4212 5868 5264 5896
rect 4212 5856 4218 5868
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 7466 5896 7472 5908
rect 7379 5868 7472 5896
rect 7466 5856 7472 5868
rect 7524 5896 7530 5908
rect 10226 5896 10232 5908
rect 7524 5868 10232 5896
rect 7524 5856 7530 5868
rect 10226 5856 10232 5868
rect 10284 5856 10290 5908
rect 12894 5856 12900 5908
rect 12952 5896 12958 5908
rect 13725 5899 13783 5905
rect 13725 5896 13737 5899
rect 12952 5868 13737 5896
rect 12952 5856 12958 5868
rect 13725 5865 13737 5868
rect 13771 5865 13783 5899
rect 13725 5859 13783 5865
rect 14550 5856 14556 5908
rect 14608 5896 14614 5908
rect 14645 5899 14703 5905
rect 14645 5896 14657 5899
rect 14608 5868 14657 5896
rect 14608 5856 14614 5868
rect 14645 5865 14657 5868
rect 14691 5865 14703 5899
rect 14645 5859 14703 5865
rect 14826 5856 14832 5908
rect 14884 5896 14890 5908
rect 14884 5868 16528 5896
rect 14884 5856 14890 5868
rect 3421 5831 3479 5837
rect 3421 5797 3433 5831
rect 3467 5828 3479 5831
rect 3467 5800 4200 5828
rect 3467 5797 3479 5800
rect 3421 5791 3479 5797
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 4172 5769 4200 5800
rect 6362 5788 6368 5840
rect 6420 5788 6426 5840
rect 3329 5763 3387 5769
rect 3329 5729 3341 5763
rect 3375 5729 3387 5763
rect 3329 5723 3387 5729
rect 3513 5763 3571 5769
rect 3513 5729 3525 5763
rect 3559 5729 3571 5763
rect 3513 5723 3571 5729
rect 3697 5763 3755 5769
rect 3697 5729 3709 5763
rect 3743 5760 3755 5763
rect 3881 5763 3939 5769
rect 3881 5760 3893 5763
rect 3743 5732 3893 5760
rect 3743 5729 3755 5732
rect 3697 5723 3755 5729
rect 3881 5729 3893 5732
rect 3927 5729 3939 5763
rect 3881 5723 3939 5729
rect 3973 5763 4031 5769
rect 3973 5729 3985 5763
rect 4019 5729 4031 5763
rect 3973 5723 4031 5729
rect 4157 5763 4215 5769
rect 4157 5729 4169 5763
rect 4203 5760 4215 5763
rect 4246 5760 4252 5772
rect 4203 5732 4252 5760
rect 4203 5729 4215 5732
rect 4157 5723 4215 5729
rect 3344 5692 3372 5723
rect 3418 5692 3424 5704
rect 3344 5664 3424 5692
rect 3418 5652 3424 5664
rect 3476 5652 3482 5704
rect 3528 5692 3556 5723
rect 3988 5692 4016 5723
rect 4246 5720 4252 5732
rect 4304 5720 4310 5772
rect 7374 5720 7380 5772
rect 7432 5760 7438 5772
rect 7484 5760 7512 5856
rect 10045 5831 10103 5837
rect 10045 5797 10057 5831
rect 10091 5828 10103 5831
rect 10502 5828 10508 5840
rect 10091 5800 10508 5828
rect 10091 5797 10103 5800
rect 10045 5791 10103 5797
rect 10502 5788 10508 5800
rect 10560 5788 10566 5840
rect 12250 5828 12256 5840
rect 12211 5800 12256 5828
rect 12250 5788 12256 5800
rect 12308 5788 12314 5840
rect 13262 5788 13268 5840
rect 13320 5788 13326 5840
rect 15930 5828 15936 5840
rect 15778 5800 15936 5828
rect 15930 5788 15936 5800
rect 15988 5788 15994 5840
rect 16209 5831 16267 5837
rect 16209 5797 16221 5831
rect 16255 5828 16267 5831
rect 16298 5828 16304 5840
rect 16255 5800 16304 5828
rect 16255 5797 16267 5800
rect 16209 5791 16267 5797
rect 16298 5788 16304 5800
rect 16356 5788 16362 5840
rect 7432 5732 7525 5760
rect 7432 5720 7438 5732
rect 8846 5720 8852 5772
rect 8904 5760 8910 5772
rect 9309 5763 9367 5769
rect 9309 5760 9321 5763
rect 8904 5732 9321 5760
rect 8904 5720 8910 5732
rect 9309 5729 9321 5732
rect 9355 5729 9367 5763
rect 9309 5723 9367 5729
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5729 9735 5763
rect 10134 5760 10140 5772
rect 10095 5732 10140 5760
rect 9677 5723 9735 5729
rect 4614 5692 4620 5704
rect 3528 5664 4620 5692
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 7098 5692 7104 5704
rect 7059 5664 7104 5692
rect 7098 5652 7104 5664
rect 7156 5652 7162 5704
rect 7558 5652 7564 5704
rect 7616 5692 7622 5704
rect 8386 5692 8392 5704
rect 7616 5664 8392 5692
rect 7616 5652 7622 5664
rect 8386 5652 8392 5664
rect 8444 5692 8450 5704
rect 9401 5695 9459 5701
rect 9401 5692 9413 5695
rect 8444 5664 9413 5692
rect 8444 5652 8450 5664
rect 9401 5661 9413 5664
rect 9447 5661 9459 5695
rect 9401 5655 9459 5661
rect 9214 5584 9220 5636
rect 9272 5624 9278 5636
rect 9692 5624 9720 5723
rect 10134 5720 10140 5732
rect 10192 5720 10198 5772
rect 14458 5760 14464 5772
rect 14419 5732 14464 5760
rect 14458 5720 14464 5732
rect 14516 5720 14522 5772
rect 16500 5769 16528 5868
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5729 16543 5763
rect 16485 5723 16543 5729
rect 9950 5692 9956 5704
rect 9911 5664 9956 5692
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 11977 5695 12035 5701
rect 11977 5692 11989 5695
rect 10284 5664 11989 5692
rect 10284 5652 10290 5664
rect 11977 5661 11989 5664
rect 12023 5692 12035 5695
rect 13814 5692 13820 5704
rect 12023 5664 13820 5692
rect 12023 5661 12035 5664
rect 11977 5655 12035 5661
rect 13814 5652 13820 5664
rect 13872 5652 13878 5704
rect 9272 5596 9720 5624
rect 9272 5584 9278 5596
rect 3142 5556 3148 5568
rect 3103 5528 3148 5556
rect 3142 5516 3148 5528
rect 3200 5516 3206 5568
rect 4154 5556 4160 5568
rect 4115 5528 4160 5556
rect 4154 5516 4160 5528
rect 4212 5516 4218 5568
rect 5442 5516 5448 5568
rect 5500 5556 5506 5568
rect 5629 5559 5687 5565
rect 5629 5556 5641 5559
rect 5500 5528 5641 5556
rect 5500 5516 5506 5528
rect 5629 5525 5641 5528
rect 5675 5525 5687 5559
rect 5629 5519 5687 5525
rect 14737 5559 14795 5565
rect 14737 5525 14749 5559
rect 14783 5556 14795 5559
rect 14826 5556 14832 5568
rect 14783 5528 14832 5556
rect 14783 5525 14795 5528
rect 14737 5519 14795 5525
rect 14826 5516 14832 5528
rect 14884 5516 14890 5568
rect 1104 5466 16836 5488
rect 1104 5414 3604 5466
rect 3656 5414 3668 5466
rect 3720 5414 3732 5466
rect 3784 5414 3796 5466
rect 3848 5414 8848 5466
rect 8900 5414 8912 5466
rect 8964 5414 8976 5466
rect 9028 5414 9040 5466
rect 9092 5414 14092 5466
rect 14144 5414 14156 5466
rect 14208 5414 14220 5466
rect 14272 5414 14284 5466
rect 14336 5414 16836 5466
rect 1104 5392 16836 5414
rect 6273 5355 6331 5361
rect 6273 5321 6285 5355
rect 6319 5352 6331 5355
rect 6362 5352 6368 5364
rect 6319 5324 6368 5352
rect 6319 5321 6331 5324
rect 6273 5315 6331 5321
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 6457 5355 6515 5361
rect 6457 5321 6469 5355
rect 6503 5352 6515 5355
rect 7098 5352 7104 5364
rect 6503 5324 7104 5352
rect 6503 5321 6515 5324
rect 6457 5315 6515 5321
rect 7098 5312 7104 5324
rect 7156 5312 7162 5364
rect 9217 5355 9275 5361
rect 9217 5321 9229 5355
rect 9263 5352 9275 5355
rect 9309 5355 9367 5361
rect 9309 5352 9321 5355
rect 9263 5324 9321 5352
rect 9263 5321 9275 5324
rect 9217 5315 9275 5321
rect 9309 5321 9321 5324
rect 9355 5352 9367 5355
rect 10134 5352 10140 5364
rect 9355 5324 10140 5352
rect 9355 5321 9367 5324
rect 9309 5315 9367 5321
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 13173 5355 13231 5361
rect 13173 5321 13185 5355
rect 13219 5352 13231 5355
rect 13262 5352 13268 5364
rect 13219 5324 13268 5352
rect 13219 5321 13231 5324
rect 13173 5315 13231 5321
rect 13262 5312 13268 5324
rect 13320 5312 13326 5364
rect 3881 5287 3939 5293
rect 3881 5253 3893 5287
rect 3927 5284 3939 5287
rect 4338 5284 4344 5296
rect 3927 5256 4344 5284
rect 3927 5253 3939 5256
rect 3881 5247 3939 5253
rect 4338 5244 4344 5256
rect 4396 5244 4402 5296
rect 4433 5287 4491 5293
rect 4433 5253 4445 5287
rect 4479 5284 4491 5287
rect 8113 5287 8171 5293
rect 4479 5256 7512 5284
rect 4479 5253 4491 5256
rect 4433 5247 4491 5253
rect 1486 5176 1492 5228
rect 1544 5216 1550 5228
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 1544 5188 1593 5216
rect 1544 5176 1550 5188
rect 1581 5185 1593 5188
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5216 1915 5219
rect 3142 5216 3148 5228
rect 1903 5188 3148 5216
rect 1903 5185 1915 5188
rect 1857 5179 1915 5185
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 3789 5219 3847 5225
rect 3789 5185 3801 5219
rect 3835 5216 3847 5219
rect 4154 5216 4160 5228
rect 3835 5188 4160 5216
rect 3835 5185 3847 5188
rect 3789 5179 3847 5185
rect 4154 5176 4160 5188
rect 4212 5216 4218 5228
rect 6914 5216 6920 5228
rect 4212 5188 4752 5216
rect 6875 5188 6920 5216
rect 4212 5176 4218 5188
rect 4308 5151 4366 5157
rect 4308 5117 4320 5151
rect 4354 5148 4366 5151
rect 4614 5148 4620 5160
rect 4354 5120 4620 5148
rect 4354 5117 4366 5120
rect 4308 5111 4366 5117
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 4724 5157 4752 5188
rect 6914 5176 6920 5188
rect 6972 5216 6978 5228
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 6972 5188 7389 5216
rect 6972 5176 6978 5188
rect 7377 5185 7389 5188
rect 7423 5185 7435 5219
rect 7484 5216 7512 5256
rect 8113 5253 8125 5287
rect 8159 5284 8171 5287
rect 11241 5287 11299 5293
rect 11241 5284 11253 5287
rect 8159 5256 9260 5284
rect 8159 5253 8171 5256
rect 8113 5247 8171 5253
rect 9232 5228 9260 5256
rect 9968 5256 11253 5284
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 7484 5188 8309 5216
rect 7377 5179 7435 5185
rect 8297 5185 8309 5188
rect 8343 5185 8355 5219
rect 8297 5179 8355 5185
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5216 8447 5219
rect 8478 5216 8484 5228
rect 8435 5188 8484 5216
rect 8435 5185 8447 5188
rect 8389 5179 8447 5185
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5117 4767 5151
rect 4709 5111 4767 5117
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5117 5043 5151
rect 6086 5148 6092 5160
rect 6047 5120 6092 5148
rect 4985 5111 5043 5117
rect 2590 5040 2596 5092
rect 2648 5040 2654 5092
rect 5000 5080 5028 5111
rect 6086 5108 6092 5120
rect 6144 5108 6150 5160
rect 6641 5151 6699 5157
rect 6641 5117 6653 5151
rect 6687 5117 6699 5151
rect 6641 5111 6699 5117
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5117 6883 5151
rect 7006 5148 7012 5160
rect 6967 5120 7012 5148
rect 6825 5111 6883 5117
rect 4264 5052 5028 5080
rect 4264 5024 4292 5052
rect 5442 5040 5448 5092
rect 5500 5080 5506 5092
rect 6656 5080 6684 5111
rect 5500 5052 6684 5080
rect 6840 5080 6868 5111
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 7190 5148 7196 5160
rect 7151 5120 7196 5148
rect 7190 5108 7196 5120
rect 7248 5108 7254 5160
rect 7282 5108 7288 5160
rect 7340 5148 7346 5160
rect 7469 5151 7527 5157
rect 7340 5120 7385 5148
rect 7340 5108 7346 5120
rect 7469 5117 7481 5151
rect 7515 5117 7527 5151
rect 8312 5148 8340 5179
rect 8478 5176 8484 5188
rect 8536 5216 8542 5228
rect 8536 5188 9076 5216
rect 8536 5176 8542 5188
rect 9048 5157 9076 5188
rect 9214 5176 9220 5228
rect 9272 5176 9278 5228
rect 9968 5225 9996 5256
rect 11241 5253 11253 5256
rect 11287 5253 11299 5287
rect 11241 5247 11299 5253
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5185 10011 5219
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 9953 5179 10011 5185
rect 10060 5188 10425 5216
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 8312 5120 8861 5148
rect 7469 5111 7527 5117
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 9033 5151 9091 5157
rect 9033 5117 9045 5151
rect 9079 5117 9091 5151
rect 9674 5148 9680 5160
rect 9635 5120 9680 5148
rect 9033 5111 9091 5117
rect 7098 5080 7104 5092
rect 6840 5052 7104 5080
rect 5500 5040 5506 5052
rect 3329 5015 3387 5021
rect 3329 4981 3341 5015
rect 3375 5012 3387 5015
rect 4246 5012 4252 5024
rect 3375 4984 4252 5012
rect 3375 4981 3387 4984
rect 3329 4975 3387 4981
rect 4246 4972 4252 4984
rect 4304 4972 4310 5024
rect 4522 4972 4528 5024
rect 4580 5012 4586 5024
rect 4580 4984 4625 5012
rect 4580 4972 4586 4984
rect 4706 4972 4712 5024
rect 4764 5012 4770 5024
rect 4893 5015 4951 5021
rect 4893 5012 4905 5015
rect 4764 4984 4905 5012
rect 4764 4972 4770 4984
rect 4893 4981 4905 4984
rect 4939 5012 4951 5015
rect 5460 5012 5488 5040
rect 4939 4984 5488 5012
rect 6656 5012 6684 5052
rect 7098 5040 7104 5052
rect 7156 5080 7162 5092
rect 7484 5080 7512 5111
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 9858 5148 9864 5160
rect 9819 5120 9864 5148
rect 9858 5108 9864 5120
rect 9916 5108 9922 5160
rect 10060 5157 10088 5188
rect 10413 5185 10425 5188
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 11532 5188 12020 5216
rect 10045 5151 10103 5157
rect 10045 5117 10057 5151
rect 10091 5117 10103 5151
rect 10226 5148 10232 5160
rect 10187 5120 10232 5148
rect 10045 5111 10103 5117
rect 10226 5108 10232 5120
rect 10284 5108 10290 5160
rect 10502 5148 10508 5160
rect 10463 5120 10508 5148
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 11330 5108 11336 5160
rect 11388 5148 11394 5160
rect 11532 5157 11560 5188
rect 11517 5151 11575 5157
rect 11517 5148 11529 5151
rect 11388 5120 11529 5148
rect 11388 5108 11394 5120
rect 11517 5117 11529 5120
rect 11563 5117 11575 5151
rect 11882 5148 11888 5160
rect 11843 5120 11888 5148
rect 11517 5111 11575 5117
rect 11882 5108 11888 5120
rect 11940 5108 11946 5160
rect 11992 5157 12020 5188
rect 11977 5151 12035 5157
rect 11977 5117 11989 5151
rect 12023 5117 12035 5151
rect 11977 5111 12035 5117
rect 12161 5151 12219 5157
rect 12161 5117 12173 5151
rect 12207 5117 12219 5151
rect 12986 5148 12992 5160
rect 12947 5120 12992 5148
rect 12161 5111 12219 5117
rect 7156 5052 7512 5080
rect 9493 5083 9551 5089
rect 7156 5040 7162 5052
rect 9493 5049 9505 5083
rect 9539 5080 9551 5083
rect 10962 5080 10968 5092
rect 9539 5052 10968 5080
rect 9539 5049 9551 5052
rect 9493 5043 9551 5049
rect 10962 5040 10968 5052
rect 11020 5040 11026 5092
rect 11238 5080 11244 5092
rect 11199 5052 11244 5080
rect 11238 5040 11244 5052
rect 11296 5040 11302 5092
rect 11425 5083 11483 5089
rect 11425 5049 11437 5083
rect 11471 5080 11483 5083
rect 12066 5080 12072 5092
rect 11471 5052 12072 5080
rect 11471 5049 11483 5052
rect 11425 5043 11483 5049
rect 12066 5040 12072 5052
rect 12124 5080 12130 5092
rect 12176 5080 12204 5111
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 12124 5052 12204 5080
rect 12124 5040 12130 5052
rect 6914 5012 6920 5024
rect 6656 4984 6920 5012
rect 4939 4981 4951 4984
rect 4893 4975 4951 4981
rect 6914 4972 6920 4984
rect 6972 5012 6978 5024
rect 7282 5012 7288 5024
rect 6972 4984 7288 5012
rect 6972 4972 6978 4984
rect 7282 4972 7288 4984
rect 7340 4972 7346 5024
rect 8757 5015 8815 5021
rect 8757 4981 8769 5015
rect 8803 5012 8815 5015
rect 9309 5015 9367 5021
rect 9309 5012 9321 5015
rect 8803 4984 9321 5012
rect 8803 4981 8815 4984
rect 8757 4975 8815 4981
rect 9309 4981 9321 4984
rect 9355 4981 9367 5015
rect 11790 5012 11796 5024
rect 11751 4984 11796 5012
rect 9309 4975 9367 4981
rect 11790 4972 11796 4984
rect 11848 4972 11854 5024
rect 12161 5015 12219 5021
rect 12161 4981 12173 5015
rect 12207 5012 12219 5015
rect 12710 5012 12716 5024
rect 12207 4984 12716 5012
rect 12207 4981 12219 4984
rect 12161 4975 12219 4981
rect 12710 4972 12716 4984
rect 12768 4972 12774 5024
rect 1104 4922 16836 4944
rect 1104 4870 6226 4922
rect 6278 4870 6290 4922
rect 6342 4870 6354 4922
rect 6406 4870 6418 4922
rect 6470 4870 11470 4922
rect 11522 4870 11534 4922
rect 11586 4870 11598 4922
rect 11650 4870 11662 4922
rect 11714 4870 16836 4922
rect 1104 4848 16836 4870
rect 5534 4768 5540 4820
rect 5592 4768 5598 4820
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 9858 4808 9864 4820
rect 9723 4780 9864 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 11238 4768 11244 4820
rect 11296 4768 11302 4820
rect 16301 4811 16359 4817
rect 16301 4808 16313 4811
rect 12406 4780 16313 4808
rect 3973 4743 4031 4749
rect 3973 4709 3985 4743
rect 4019 4740 4031 4743
rect 4019 4712 4476 4740
rect 4019 4709 4031 4712
rect 3973 4703 4031 4709
rect 4065 4675 4123 4681
rect 4065 4641 4077 4675
rect 4111 4672 4123 4675
rect 4338 4672 4344 4684
rect 4111 4644 4344 4672
rect 4111 4641 4123 4644
rect 4065 4635 4123 4641
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 4448 4681 4476 4712
rect 4433 4675 4491 4681
rect 4433 4641 4445 4675
rect 4479 4672 4491 4675
rect 4522 4672 4528 4684
rect 4479 4644 4528 4672
rect 4479 4641 4491 4644
rect 4433 4635 4491 4641
rect 4522 4632 4528 4644
rect 4580 4632 4586 4684
rect 5555 4681 5583 4768
rect 9493 4743 9551 4749
rect 9493 4709 9505 4743
rect 9539 4740 9551 4743
rect 10045 4743 10103 4749
rect 9539 4712 9904 4740
rect 9539 4709 9551 4712
rect 9493 4703 9551 4709
rect 5718 4681 5724 4684
rect 5261 4675 5319 4681
rect 5261 4641 5273 4675
rect 5307 4641 5319 4675
rect 5261 4635 5319 4641
rect 5440 4675 5498 4681
rect 5440 4641 5452 4675
rect 5486 4641 5498 4675
rect 5555 4675 5614 4681
rect 5555 4644 5568 4675
rect 5440 4635 5498 4641
rect 5556 4641 5568 4644
rect 5602 4641 5614 4675
rect 5556 4635 5614 4641
rect 5675 4675 5724 4681
rect 5675 4641 5687 4675
rect 5721 4641 5724 4675
rect 5675 4635 5724 4641
rect 5276 4536 5304 4635
rect 5460 4604 5488 4635
rect 5718 4632 5724 4635
rect 5776 4632 5782 4684
rect 5994 4672 6000 4684
rect 5955 4644 6000 4672
rect 5994 4632 6000 4644
rect 6052 4632 6058 4684
rect 6178 4672 6184 4684
rect 6139 4644 6184 4672
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 9214 4672 9220 4684
rect 9175 4644 9220 4672
rect 9214 4632 9220 4644
rect 9272 4632 9278 4684
rect 9398 4672 9404 4684
rect 9359 4644 9404 4672
rect 9398 4632 9404 4644
rect 9456 4632 9462 4684
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4641 9643 4675
rect 9876 4672 9904 4712
rect 10045 4709 10057 4743
rect 10091 4740 10103 4743
rect 10318 4740 10324 4752
rect 10091 4712 10324 4740
rect 10091 4709 10103 4712
rect 10045 4703 10103 4709
rect 10318 4700 10324 4712
rect 10376 4700 10382 4752
rect 11256 4740 11284 4768
rect 11977 4743 12035 4749
rect 11977 4740 11989 4743
rect 11072 4712 11989 4740
rect 10137 4675 10195 4681
rect 10137 4672 10149 4675
rect 9876 4644 10149 4672
rect 9585 4635 9643 4641
rect 10137 4641 10149 4644
rect 10183 4672 10195 4675
rect 10226 4672 10232 4684
rect 10183 4644 10232 4672
rect 10183 4641 10195 4644
rect 10137 4635 10195 4641
rect 6365 4607 6423 4613
rect 6365 4604 6377 4607
rect 5460 4576 6377 4604
rect 6365 4573 6377 4576
rect 6411 4604 6423 4607
rect 9600 4604 9628 4635
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 10413 4675 10471 4681
rect 10413 4672 10425 4675
rect 10336 4644 10425 4672
rect 6411 4576 9628 4604
rect 6411 4573 6423 4576
rect 6365 4567 6423 4573
rect 5718 4536 5724 4548
rect 5276 4508 5724 4536
rect 5718 4496 5724 4508
rect 5776 4496 5782 4548
rect 5905 4539 5963 4545
rect 5905 4505 5917 4539
rect 5951 4536 5963 4539
rect 10336 4536 10364 4644
rect 10413 4641 10425 4644
rect 10459 4672 10471 4675
rect 10502 4672 10508 4684
rect 10459 4644 10508 4672
rect 10459 4641 10471 4644
rect 10413 4635 10471 4641
rect 10502 4632 10508 4644
rect 10560 4632 10566 4684
rect 11072 4681 11100 4712
rect 11977 4709 11989 4712
rect 12023 4709 12035 4743
rect 11977 4703 12035 4709
rect 11057 4675 11115 4681
rect 11057 4641 11069 4675
rect 11103 4641 11115 4675
rect 11238 4672 11244 4684
rect 11199 4644 11244 4672
rect 11057 4635 11115 4641
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 11790 4672 11796 4684
rect 11751 4644 11796 4672
rect 11790 4632 11796 4644
rect 11848 4632 11854 4684
rect 12066 4632 12072 4684
rect 12124 4672 12130 4684
rect 12161 4675 12219 4681
rect 12161 4672 12173 4675
rect 12124 4644 12173 4672
rect 12124 4632 12130 4644
rect 12161 4641 12173 4644
rect 12207 4672 12219 4675
rect 12406 4672 12434 4780
rect 16301 4777 16313 4780
rect 16347 4777 16359 4811
rect 16301 4771 16359 4777
rect 14734 4740 14740 4752
rect 12610 4712 14740 4740
rect 12610 4681 12638 4712
rect 14734 4700 14740 4712
rect 14792 4700 14798 4752
rect 12207 4644 12434 4672
rect 12557 4675 12638 4681
rect 12207 4641 12219 4644
rect 12161 4635 12219 4641
rect 12557 4641 12569 4675
rect 12603 4641 12638 4675
rect 12710 4672 12716 4684
rect 12671 4644 12716 4672
rect 12557 4635 12638 4641
rect 11330 4564 11336 4616
rect 11388 4604 11394 4616
rect 12345 4607 12403 4613
rect 12345 4604 12357 4607
rect 11388 4576 12357 4604
rect 11388 4564 11394 4576
rect 12345 4573 12357 4576
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 12492 4576 12537 4604
rect 12492 4564 12498 4576
rect 5951 4508 10364 4536
rect 5951 4505 5963 4508
rect 5905 4499 5963 4505
rect 11882 4496 11888 4548
rect 11940 4536 11946 4548
rect 12610 4536 12638 4635
rect 12710 4632 12716 4644
rect 12768 4632 12774 4684
rect 12986 4632 12992 4684
rect 13044 4672 13050 4684
rect 14001 4675 14059 4681
rect 14001 4672 14013 4675
rect 13044 4644 14013 4672
rect 13044 4632 13050 4644
rect 14001 4641 14013 4644
rect 14047 4672 14059 4675
rect 14458 4672 14464 4684
rect 14047 4644 14464 4672
rect 14047 4641 14059 4644
rect 14001 4635 14059 4641
rect 14458 4632 14464 4644
rect 14516 4672 14522 4684
rect 15473 4675 15531 4681
rect 15473 4672 15485 4675
rect 14516 4644 15485 4672
rect 14516 4632 14522 4644
rect 15473 4641 15485 4644
rect 15519 4641 15531 4675
rect 16482 4672 16488 4684
rect 16443 4644 16488 4672
rect 15473 4635 15531 4641
rect 16482 4632 16488 4644
rect 16540 4632 16546 4684
rect 15194 4536 15200 4548
rect 11940 4508 12638 4536
rect 13648 4508 15200 4536
rect 11940 4496 11946 4508
rect 4617 4471 4675 4477
rect 4617 4437 4629 4471
rect 4663 4468 4675 4471
rect 5074 4468 5080 4480
rect 4663 4440 5080 4468
rect 4663 4437 4675 4440
rect 4617 4431 4675 4437
rect 5074 4428 5080 4440
rect 5132 4468 5138 4480
rect 5994 4468 6000 4480
rect 5132 4440 6000 4468
rect 5132 4428 5138 4440
rect 5994 4428 6000 4440
rect 6052 4428 6058 4480
rect 9398 4428 9404 4480
rect 9456 4468 9462 4480
rect 9950 4468 9956 4480
rect 9456 4440 9956 4468
rect 9456 4428 9462 4440
rect 9950 4428 9956 4440
rect 10008 4468 10014 4480
rect 13648 4468 13676 4508
rect 15194 4496 15200 4508
rect 15252 4496 15258 4548
rect 13814 4468 13820 4480
rect 10008 4440 13676 4468
rect 13775 4440 13820 4468
rect 10008 4428 10014 4440
rect 13814 4428 13820 4440
rect 13872 4428 13878 4480
rect 15562 4428 15568 4480
rect 15620 4468 15626 4480
rect 15657 4471 15715 4477
rect 15657 4468 15669 4471
rect 15620 4440 15669 4468
rect 15620 4428 15626 4440
rect 15657 4437 15669 4440
rect 15703 4437 15715 4471
rect 15657 4431 15715 4437
rect 1104 4378 16836 4400
rect 1104 4326 3604 4378
rect 3656 4326 3668 4378
rect 3720 4326 3732 4378
rect 3784 4326 3796 4378
rect 3848 4326 8848 4378
rect 8900 4326 8912 4378
rect 8964 4326 8976 4378
rect 9028 4326 9040 4378
rect 9092 4326 14092 4378
rect 14144 4326 14156 4378
rect 14208 4326 14220 4378
rect 14272 4326 14284 4378
rect 14336 4326 16836 4378
rect 1104 4304 16836 4326
rect 6178 4264 6184 4276
rect 5552 4236 6184 4264
rect 5552 4196 5580 4236
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 9674 4264 9680 4276
rect 6748 4236 9680 4264
rect 5368 4168 5580 4196
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5368 4128 5396 4168
rect 5626 4156 5632 4208
rect 5684 4156 5690 4208
rect 5718 4156 5724 4208
rect 5776 4196 5782 4208
rect 6748 4196 6776 4236
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 10134 4224 10140 4276
rect 10192 4264 10198 4276
rect 12986 4264 12992 4276
rect 10192 4236 12992 4264
rect 10192 4224 10198 4236
rect 12986 4224 12992 4236
rect 13044 4224 13050 4276
rect 14826 4273 14832 4276
rect 14816 4267 14832 4273
rect 14816 4233 14828 4267
rect 14816 4227 14832 4233
rect 14826 4224 14832 4227
rect 14884 4224 14890 4276
rect 12434 4196 12440 4208
rect 5776 4168 6776 4196
rect 5776 4156 5782 4168
rect 12406 4156 12440 4196
rect 12492 4156 12498 4208
rect 5644 4128 5672 4156
rect 4948 4100 5396 4128
rect 5460 4100 5672 4128
rect 4948 4088 4954 4100
rect 5074 4060 5080 4072
rect 5035 4032 5080 4060
rect 5074 4020 5080 4032
rect 5132 4020 5138 4072
rect 5184 4069 5212 4100
rect 5460 4069 5488 4100
rect 7006 4088 7012 4140
rect 7064 4128 7070 4140
rect 11333 4131 11391 4137
rect 7064 4100 7144 4128
rect 7064 4088 7070 4100
rect 5169 4063 5227 4069
rect 5169 4029 5181 4063
rect 5215 4029 5227 4063
rect 5169 4023 5227 4029
rect 5445 4063 5503 4069
rect 5445 4029 5457 4063
rect 5491 4029 5503 4063
rect 5626 4060 5632 4072
rect 5587 4032 5632 4060
rect 5445 4023 5503 4029
rect 1578 3952 1584 4004
rect 1636 3992 1642 4004
rect 5460 3992 5488 4023
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 6638 4060 6644 4072
rect 6599 4032 6644 4060
rect 6638 4020 6644 4032
rect 6696 4020 6702 4072
rect 6730 4020 6736 4072
rect 6788 4060 6794 4072
rect 7116 4069 7144 4100
rect 11333 4097 11345 4131
rect 11379 4128 11391 4131
rect 12406 4128 12434 4156
rect 11379 4100 12434 4128
rect 12713 4131 12771 4137
rect 11379 4097 11391 4100
rect 11333 4091 11391 4097
rect 12713 4097 12725 4131
rect 12759 4128 12771 4131
rect 13722 4128 13728 4140
rect 12759 4100 13728 4128
rect 12759 4097 12771 4100
rect 12713 4091 12771 4097
rect 13722 4088 13728 4100
rect 13780 4128 13786 4140
rect 14550 4128 14556 4140
rect 13780 4100 14556 4128
rect 13780 4088 13786 4100
rect 14550 4088 14556 4100
rect 14608 4088 14614 4140
rect 7101 4063 7159 4069
rect 6788 4032 6833 4060
rect 6788 4020 6794 4032
rect 7101 4029 7113 4063
rect 7147 4029 7159 4063
rect 7374 4060 7380 4072
rect 7335 4032 7380 4060
rect 7101 4023 7159 4029
rect 7374 4020 7380 4032
rect 7432 4020 7438 4072
rect 11238 4060 11244 4072
rect 11199 4032 11244 4060
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 12066 4060 12072 4072
rect 12027 4032 12072 4060
rect 12066 4020 12072 4032
rect 12124 4020 12130 4072
rect 12253 4063 12311 4069
rect 12253 4060 12265 4063
rect 12176 4032 12265 4060
rect 1636 3964 5488 3992
rect 1636 3952 1642 3964
rect 6822 3952 6828 4004
rect 6880 3992 6886 4004
rect 6917 3995 6975 4001
rect 6917 3992 6929 3995
rect 6880 3964 6929 3992
rect 6880 3952 6886 3964
rect 6917 3961 6929 3964
rect 6963 3961 6975 3995
rect 6917 3955 6975 3961
rect 7012 3995 7070 4001
rect 7012 3961 7024 3995
rect 7058 3992 7070 3995
rect 7640 3995 7698 4001
rect 7640 3992 7652 3995
rect 7058 3964 7144 3992
rect 7058 3961 7070 3964
rect 7012 3955 7070 3961
rect 7116 3936 7144 3964
rect 7300 3964 7652 3992
rect 4430 3884 4436 3936
rect 4488 3924 4494 3936
rect 5258 3924 5264 3936
rect 4488 3896 5264 3924
rect 4488 3884 4494 3896
rect 5258 3884 5264 3896
rect 5316 3924 5322 3936
rect 6638 3924 6644 3936
rect 5316 3896 6644 3924
rect 5316 3884 5322 3896
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 7098 3884 7104 3936
rect 7156 3884 7162 3936
rect 7300 3933 7328 3964
rect 7640 3961 7652 3964
rect 7686 3961 7698 3995
rect 7640 3955 7698 3961
rect 8662 3952 8668 4004
rect 8720 3952 8726 4004
rect 7285 3927 7343 3933
rect 7285 3893 7297 3927
rect 7331 3893 7343 3927
rect 7285 3887 7343 3893
rect 9125 3927 9183 3933
rect 9125 3893 9137 3927
rect 9171 3924 9183 3927
rect 10042 3924 10048 3936
rect 9171 3896 10048 3924
rect 9171 3893 9183 3896
rect 9125 3887 9183 3893
rect 10042 3884 10048 3896
rect 10100 3924 10106 3936
rect 12176 3924 12204 4032
rect 12253 4029 12265 4032
rect 12299 4029 12311 4063
rect 12253 4023 12311 4029
rect 12434 4020 12440 4072
rect 12492 4060 12498 4072
rect 12492 4032 12537 4060
rect 12492 4020 12498 4032
rect 12342 3992 12348 4004
rect 12303 3964 12348 3992
rect 12342 3952 12348 3964
rect 12400 3952 12406 4004
rect 12989 3995 13047 4001
rect 12989 3961 13001 3995
rect 13035 3961 13047 3995
rect 12989 3955 13047 3961
rect 10100 3896 12204 3924
rect 12621 3927 12679 3933
rect 10100 3884 10106 3896
rect 12621 3893 12633 3927
rect 12667 3924 12679 3927
rect 13004 3924 13032 3955
rect 13832 3936 13860 3978
rect 15562 3952 15568 4004
rect 15620 3952 15626 4004
rect 12667 3896 13032 3924
rect 12667 3893 12679 3896
rect 12621 3887 12679 3893
rect 13814 3884 13820 3936
rect 13872 3884 13878 3936
rect 14458 3924 14464 3936
rect 14419 3896 14464 3924
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 16301 3927 16359 3933
rect 16301 3893 16313 3927
rect 16347 3924 16359 3927
rect 16390 3924 16396 3936
rect 16347 3896 16396 3924
rect 16347 3893 16359 3896
rect 16301 3887 16359 3893
rect 16390 3884 16396 3896
rect 16448 3884 16454 3936
rect 1104 3834 16836 3856
rect 1104 3782 6226 3834
rect 6278 3782 6290 3834
rect 6342 3782 6354 3834
rect 6406 3782 6418 3834
rect 6470 3782 11470 3834
rect 11522 3782 11534 3834
rect 11586 3782 11598 3834
rect 11650 3782 11662 3834
rect 11714 3782 16836 3834
rect 1104 3760 16836 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 4338 3680 4344 3732
rect 4396 3720 4402 3732
rect 4433 3723 4491 3729
rect 4433 3720 4445 3723
rect 4396 3692 4445 3720
rect 4396 3680 4402 3692
rect 4433 3689 4445 3692
rect 4479 3689 4491 3723
rect 4433 3683 4491 3689
rect 4617 3723 4675 3729
rect 4617 3689 4629 3723
rect 4663 3720 4675 3723
rect 5166 3720 5172 3732
rect 4663 3692 5172 3720
rect 4663 3689 4675 3692
rect 4617 3683 4675 3689
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 7006 3680 7012 3732
rect 7064 3720 7070 3732
rect 7193 3723 7251 3729
rect 7193 3720 7205 3723
rect 7064 3692 7205 3720
rect 7064 3680 7070 3692
rect 7193 3689 7205 3692
rect 7239 3689 7251 3723
rect 7193 3683 7251 3689
rect 8573 3723 8631 3729
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 8662 3720 8668 3732
rect 8619 3692 8668 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 11882 3680 11888 3732
rect 11940 3720 11946 3732
rect 12069 3723 12127 3729
rect 12069 3720 12081 3723
rect 11940 3692 12081 3720
rect 11940 3680 11946 3692
rect 12069 3689 12081 3692
rect 12115 3689 12127 3723
rect 12069 3683 12127 3689
rect 6086 3652 6092 3664
rect 3160 3624 6092 3652
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 2317 3587 2375 3593
rect 2317 3553 2329 3587
rect 2363 3584 2375 3587
rect 2590 3584 2596 3596
rect 2363 3556 2596 3584
rect 2363 3553 2375 3556
rect 2317 3547 2375 3553
rect 2590 3544 2596 3556
rect 2648 3584 2654 3596
rect 3160 3593 3188 3624
rect 6086 3612 6092 3624
rect 6144 3652 6150 3664
rect 11900 3652 11928 3680
rect 6144 3624 8432 3652
rect 6144 3612 6150 3624
rect 3145 3587 3203 3593
rect 3145 3584 3157 3587
rect 2648 3556 3157 3584
rect 2648 3544 2654 3556
rect 3145 3553 3157 3556
rect 3191 3553 3203 3587
rect 3145 3547 3203 3553
rect 3418 3544 3424 3596
rect 3476 3584 3482 3596
rect 4614 3593 4620 3596
rect 4558 3587 4620 3593
rect 4558 3584 4570 3587
rect 3476 3556 4570 3584
rect 3476 3544 3482 3556
rect 4558 3553 4570 3556
rect 4604 3553 4620 3587
rect 4558 3547 4620 3553
rect 4614 3544 4620 3547
rect 4672 3584 4678 3596
rect 5166 3584 5172 3596
rect 4672 3556 4706 3584
rect 5127 3556 5172 3584
rect 4672 3544 4678 3556
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 5353 3587 5411 3593
rect 5353 3553 5365 3587
rect 5399 3553 5411 3587
rect 6914 3584 6920 3596
rect 6875 3556 6920 3584
rect 5353 3547 5411 3553
rect 4982 3476 4988 3528
rect 5040 3516 5046 3528
rect 5077 3519 5135 3525
rect 5077 3516 5089 3519
rect 5040 3488 5089 3516
rect 5040 3476 5046 3488
rect 5077 3485 5089 3488
rect 5123 3516 5135 3519
rect 5261 3519 5319 3525
rect 5261 3516 5273 3519
rect 5123 3488 5273 3516
rect 5123 3485 5135 3488
rect 5077 3479 5135 3485
rect 5261 3485 5273 3488
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 4614 3408 4620 3460
rect 4672 3448 4678 3460
rect 5368 3448 5396 3547
rect 6914 3544 6920 3556
rect 6972 3544 6978 3596
rect 7098 3584 7104 3596
rect 7059 3556 7104 3584
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 7190 3544 7196 3596
rect 7248 3584 7254 3596
rect 8404 3593 8432 3624
rect 10980 3624 11928 3652
rect 7285 3587 7343 3593
rect 7285 3584 7297 3587
rect 7248 3556 7297 3584
rect 7248 3544 7254 3556
rect 7285 3553 7297 3556
rect 7331 3553 7343 3587
rect 7285 3547 7343 3553
rect 8389 3587 8447 3593
rect 8389 3553 8401 3587
rect 8435 3584 8447 3587
rect 10134 3584 10140 3596
rect 8435 3556 10140 3584
rect 8435 3553 8447 3556
rect 8389 3547 8447 3553
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 10980 3593 11008 3624
rect 12342 3612 12348 3664
rect 12400 3652 12406 3664
rect 12400 3624 13032 3652
rect 12400 3612 12406 3624
rect 10965 3587 11023 3593
rect 10965 3553 10977 3587
rect 11011 3553 11023 3587
rect 10965 3547 11023 3553
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 13004 3593 13032 3624
rect 15764 3624 16344 3652
rect 11333 3587 11391 3593
rect 11333 3584 11345 3587
rect 11204 3556 11345 3584
rect 11204 3544 11210 3556
rect 11333 3553 11345 3556
rect 11379 3584 11391 3587
rect 11977 3587 12035 3593
rect 11977 3584 11989 3587
rect 11379 3556 11989 3584
rect 11379 3553 11391 3556
rect 11333 3547 11391 3553
rect 11977 3553 11989 3556
rect 12023 3553 12035 3587
rect 12529 3587 12587 3593
rect 12529 3584 12541 3587
rect 11977 3547 12035 3553
rect 12406 3556 12541 3584
rect 6638 3476 6644 3528
rect 6696 3516 6702 3528
rect 11793 3519 11851 3525
rect 6696 3488 11376 3516
rect 6696 3476 6702 3488
rect 4672 3420 5396 3448
rect 4672 3408 4678 3420
rect 7282 3408 7288 3460
rect 7340 3448 7346 3460
rect 7469 3451 7527 3457
rect 7469 3448 7481 3451
rect 7340 3420 7481 3448
rect 7340 3408 7346 3420
rect 7469 3417 7481 3420
rect 7515 3448 7527 3451
rect 9398 3448 9404 3460
rect 7515 3420 9404 3448
rect 7515 3417 7527 3420
rect 7469 3411 7527 3417
rect 9398 3408 9404 3420
rect 9456 3408 9462 3460
rect 11057 3451 11115 3457
rect 11057 3417 11069 3451
rect 11103 3448 11115 3451
rect 11238 3448 11244 3460
rect 11103 3420 11244 3448
rect 11103 3417 11115 3420
rect 11057 3411 11115 3417
rect 11238 3408 11244 3420
rect 11296 3408 11302 3460
rect 11348 3448 11376 3488
rect 11793 3485 11805 3519
rect 11839 3516 11851 3519
rect 12406 3516 12434 3556
rect 12529 3553 12541 3556
rect 12575 3584 12587 3587
rect 12897 3587 12955 3593
rect 12897 3584 12909 3587
rect 12575 3556 12909 3584
rect 12575 3553 12587 3556
rect 12529 3547 12587 3553
rect 12897 3553 12909 3556
rect 12943 3553 12955 3587
rect 12897 3547 12955 3553
rect 12989 3587 13047 3593
rect 12989 3553 13001 3587
rect 13035 3584 13047 3587
rect 14458 3584 14464 3596
rect 13035 3556 14464 3584
rect 13035 3553 13047 3556
rect 12989 3547 13047 3553
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 15562 3584 15568 3596
rect 15523 3556 15568 3584
rect 15562 3544 15568 3556
rect 15620 3544 15626 3596
rect 15764 3593 15792 3624
rect 16316 3596 16344 3624
rect 15749 3587 15807 3593
rect 15749 3553 15761 3587
rect 15795 3553 15807 3587
rect 15749 3547 15807 3553
rect 16298 3544 16304 3596
rect 16356 3584 16362 3596
rect 16356 3556 16401 3584
rect 16356 3544 16362 3556
rect 16390 3516 16396 3528
rect 11839 3488 12434 3516
rect 16303 3488 16396 3516
rect 11839 3485 11851 3488
rect 11793 3479 11851 3485
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 12158 3448 12164 3460
rect 11348 3420 12164 3448
rect 12158 3408 12164 3420
rect 12216 3408 12222 3460
rect 15562 3408 15568 3460
rect 15620 3448 15626 3460
rect 16408 3448 16436 3476
rect 15620 3420 16436 3448
rect 15620 3408 15626 3420
rect 2406 3340 2412 3392
rect 2464 3380 2470 3392
rect 2501 3383 2559 3389
rect 2501 3380 2513 3383
rect 2464 3352 2513 3380
rect 2464 3340 2470 3352
rect 2501 3349 2513 3352
rect 2547 3349 2559 3383
rect 2501 3343 2559 3349
rect 3329 3383 3387 3389
rect 3329 3349 3341 3383
rect 3375 3380 3387 3383
rect 4246 3380 4252 3392
rect 3375 3352 4252 3380
rect 3375 3349 3387 3352
rect 3329 3343 3387 3349
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 4985 3383 5043 3389
rect 4985 3349 4997 3383
rect 5031 3380 5043 3383
rect 6178 3380 6184 3392
rect 5031 3352 6184 3380
rect 5031 3349 5043 3352
rect 4985 3343 5043 3349
rect 6178 3340 6184 3352
rect 6236 3340 6242 3392
rect 8386 3340 8392 3392
rect 8444 3380 8450 3392
rect 12434 3380 12440 3392
rect 8444 3352 12440 3380
rect 8444 3340 8450 3352
rect 12434 3340 12440 3352
rect 12492 3380 12498 3392
rect 15289 3383 15347 3389
rect 15289 3380 15301 3383
rect 12492 3352 15301 3380
rect 12492 3340 12498 3352
rect 15289 3349 15301 3352
rect 15335 3349 15347 3383
rect 15289 3343 15347 3349
rect 1104 3290 16836 3312
rect 1104 3238 3604 3290
rect 3656 3238 3668 3290
rect 3720 3238 3732 3290
rect 3784 3238 3796 3290
rect 3848 3238 8848 3290
rect 8900 3238 8912 3290
rect 8964 3238 8976 3290
rect 9028 3238 9040 3290
rect 9092 3238 14092 3290
rect 14144 3238 14156 3290
rect 14208 3238 14220 3290
rect 14272 3238 14284 3290
rect 14336 3238 16836 3290
rect 1104 3216 16836 3238
rect 1486 3136 1492 3188
rect 1544 3136 1550 3188
rect 5353 3179 5411 3185
rect 5353 3145 5365 3179
rect 5399 3176 5411 3179
rect 5626 3176 5632 3188
rect 5399 3148 5632 3176
rect 5399 3145 5411 3148
rect 5353 3139 5411 3145
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 6178 3176 6184 3188
rect 6139 3148 6184 3176
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 7098 3136 7104 3188
rect 7156 3176 7162 3188
rect 7561 3179 7619 3185
rect 7561 3176 7573 3179
rect 7156 3148 7573 3176
rect 7156 3136 7162 3148
rect 7561 3145 7573 3148
rect 7607 3145 7619 3179
rect 10594 3176 10600 3188
rect 10555 3148 10600 3176
rect 7561 3139 7619 3145
rect 10594 3136 10600 3148
rect 10652 3136 10658 3188
rect 11330 3176 11336 3188
rect 11291 3148 11336 3176
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 13170 3136 13176 3188
rect 13228 3176 13234 3188
rect 13357 3179 13415 3185
rect 13357 3176 13369 3179
rect 13228 3148 13369 3176
rect 13228 3136 13234 3148
rect 13357 3145 13369 3148
rect 13403 3145 13415 3179
rect 13357 3139 13415 3145
rect 16298 3136 16304 3188
rect 16356 3176 16362 3188
rect 16485 3179 16543 3185
rect 16485 3176 16497 3179
rect 16356 3148 16497 3176
rect 16356 3136 16362 3148
rect 16485 3145 16497 3148
rect 16531 3145 16543 3179
rect 16485 3139 16543 3145
rect 1397 3043 1455 3049
rect 1397 3009 1409 3043
rect 1443 3040 1455 3043
rect 1504 3040 1532 3136
rect 4798 3068 4804 3120
rect 4856 3108 4862 3120
rect 5166 3108 5172 3120
rect 4856 3080 5172 3108
rect 4856 3068 4862 3080
rect 5166 3068 5172 3080
rect 5224 3108 5230 3120
rect 5261 3111 5319 3117
rect 5261 3108 5273 3111
rect 5224 3080 5273 3108
rect 5224 3068 5230 3080
rect 5261 3077 5273 3080
rect 5307 3077 5319 3111
rect 5261 3071 5319 3077
rect 7089 3080 7512 3108
rect 7089 3049 7117 3080
rect 3513 3043 3571 3049
rect 3513 3040 3525 3043
rect 1443 3012 3525 3040
rect 1443 3009 1455 3012
rect 1397 3003 1455 3009
rect 3513 3009 3525 3012
rect 3559 3009 3571 3043
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 3513 3003 3571 3009
rect 5092 3012 6837 3040
rect 3418 2972 3424 2984
rect 3379 2944 3424 2972
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 1673 2907 1731 2913
rect 1673 2873 1685 2907
rect 1719 2873 1731 2907
rect 1673 2867 1731 2873
rect 1688 2836 1716 2867
rect 2406 2864 2412 2916
rect 2464 2864 2470 2916
rect 3786 2904 3792 2916
rect 3747 2876 3792 2904
rect 3786 2864 3792 2876
rect 3844 2864 3850 2916
rect 4246 2864 4252 2916
rect 4304 2864 4310 2916
rect 5092 2836 5120 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 7089 3043 7148 3049
rect 7089 3009 7102 3043
rect 7136 3009 7148 3043
rect 7089 3003 7148 3009
rect 5537 2975 5595 2981
rect 5537 2941 5549 2975
rect 5583 2941 5595 2975
rect 5537 2935 5595 2941
rect 5552 2904 5580 2935
rect 5626 2932 5632 2984
rect 5684 2972 5690 2984
rect 5905 2975 5963 2981
rect 5905 2972 5917 2975
rect 5684 2944 5917 2972
rect 5684 2932 5690 2944
rect 5905 2941 5917 2944
rect 5951 2941 5963 2975
rect 5905 2935 5963 2941
rect 6273 2975 6331 2981
rect 6273 2941 6285 2975
rect 6319 2941 6331 2975
rect 6996 2975 7054 2981
rect 6996 2972 7008 2975
rect 6273 2935 6331 2941
rect 6840 2944 7008 2972
rect 5997 2907 6055 2913
rect 5997 2904 6009 2907
rect 5552 2876 6009 2904
rect 5997 2873 6009 2876
rect 6043 2904 6055 2907
rect 6288 2904 6316 2935
rect 6840 2916 6868 2944
rect 6996 2941 7008 2944
rect 7042 2941 7054 2975
rect 6996 2935 7054 2941
rect 7089 2916 7117 3003
rect 7282 3000 7288 3052
rect 7340 3040 7346 3052
rect 7340 3012 7385 3040
rect 7340 3000 7346 3012
rect 7190 2932 7196 2984
rect 7248 2972 7254 2984
rect 7484 2981 7512 3080
rect 8754 3068 8760 3120
rect 8812 3108 8818 3120
rect 9953 3111 10011 3117
rect 9953 3108 9965 3111
rect 8812 3080 9965 3108
rect 8812 3068 8818 3080
rect 9953 3077 9965 3080
rect 9999 3108 10011 3111
rect 11146 3108 11152 3120
rect 9999 3080 11152 3108
rect 9999 3077 10011 3080
rect 9953 3071 10011 3077
rect 11146 3068 11152 3080
rect 11204 3068 11210 3120
rect 12434 3068 12440 3120
rect 12492 3108 12498 3120
rect 12989 3111 13047 3117
rect 12492 3080 12848 3108
rect 12492 3068 12498 3080
rect 11425 3043 11483 3049
rect 9140 3012 10088 3040
rect 7469 2975 7527 2981
rect 7248 2944 7293 2972
rect 7248 2932 7254 2944
rect 7469 2941 7481 2975
rect 7515 2941 7527 2975
rect 8386 2972 8392 2984
rect 8299 2944 8392 2972
rect 7469 2935 7527 2941
rect 8386 2932 8392 2944
rect 8444 2932 8450 2984
rect 8570 2972 8576 2984
rect 8531 2944 8576 2972
rect 8570 2932 8576 2944
rect 8628 2932 8634 2984
rect 8665 2975 8723 2981
rect 8665 2941 8677 2975
rect 8711 2941 8723 2975
rect 8665 2935 8723 2941
rect 6043 2876 6316 2904
rect 6043 2873 6055 2876
rect 5997 2867 6055 2873
rect 1688 2808 5120 2836
rect 6288 2836 6316 2876
rect 6822 2864 6828 2916
rect 6880 2864 6886 2916
rect 7089 2876 7104 2916
rect 7098 2864 7104 2876
rect 7156 2864 7162 2916
rect 7208 2904 7236 2932
rect 8404 2904 8432 2932
rect 7208 2876 8432 2904
rect 8680 2904 8708 2935
rect 8754 2932 8760 2984
rect 8812 2972 8818 2984
rect 8938 2972 8944 2984
rect 8812 2944 8857 2972
rect 8899 2944 8944 2972
rect 8812 2932 8818 2944
rect 8938 2932 8944 2944
rect 8996 2932 9002 2984
rect 9140 2972 9168 3012
rect 10060 2984 10088 3012
rect 11425 3009 11437 3043
rect 11471 3040 11483 3043
rect 11471 3012 11744 3040
rect 11471 3009 11483 3012
rect 11425 3003 11483 3009
rect 9398 2972 9404 2984
rect 9048 2944 9168 2972
rect 9359 2944 9404 2972
rect 9048 2904 9076 2944
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 10042 2972 10048 2984
rect 10003 2944 10048 2972
rect 10042 2932 10048 2944
rect 10100 2932 10106 2984
rect 10134 2932 10140 2984
rect 10192 2972 10198 2984
rect 10192 2944 10237 2972
rect 10192 2932 10198 2944
rect 10318 2932 10324 2984
rect 10376 2972 10382 2984
rect 10413 2975 10471 2981
rect 10413 2972 10425 2975
rect 10376 2944 10425 2972
rect 10376 2932 10382 2944
rect 10413 2941 10425 2944
rect 10459 2941 10471 2975
rect 10413 2935 10471 2941
rect 10965 2975 11023 2981
rect 10965 2941 10977 2975
rect 11011 2941 11023 2975
rect 10965 2935 11023 2941
rect 11057 2975 11115 2981
rect 11057 2941 11069 2975
rect 11103 2972 11115 2975
rect 11440 2972 11468 3003
rect 11716 2981 11744 3012
rect 12084 3012 12756 3040
rect 11103 2944 11468 2972
rect 11517 2975 11575 2981
rect 11103 2941 11115 2944
rect 11057 2935 11115 2941
rect 11517 2941 11529 2975
rect 11563 2941 11575 2975
rect 11517 2935 11575 2941
rect 11701 2975 11759 2981
rect 11701 2941 11713 2975
rect 11747 2972 11759 2975
rect 11790 2972 11796 2984
rect 11747 2944 11796 2972
rect 11747 2941 11759 2944
rect 11701 2935 11759 2941
rect 8680 2876 9076 2904
rect 9125 2907 9183 2913
rect 9125 2873 9137 2907
rect 9171 2904 9183 2907
rect 9217 2907 9275 2913
rect 9217 2904 9229 2907
rect 9171 2876 9229 2904
rect 9171 2873 9183 2876
rect 9125 2867 9183 2873
rect 9217 2873 9229 2876
rect 9263 2873 9275 2907
rect 10980 2904 11008 2935
rect 11532 2904 11560 2935
rect 11790 2932 11796 2944
rect 11848 2932 11854 2984
rect 11882 2932 11888 2984
rect 11940 2972 11946 2984
rect 12084 2981 12112 3012
rect 12069 2975 12127 2981
rect 11940 2944 11985 2972
rect 11940 2932 11946 2944
rect 12069 2941 12081 2975
rect 12115 2941 12127 2975
rect 12069 2935 12127 2941
rect 12158 2932 12164 2984
rect 12216 2972 12222 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12216 2944 12449 2972
rect 12216 2932 12222 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 11900 2904 11928 2932
rect 12728 2916 12756 3012
rect 12820 2981 12848 3080
rect 12989 3077 13001 3111
rect 13035 3108 13047 3111
rect 14090 3108 14096 3120
rect 13035 3080 14096 3108
rect 13035 3077 13047 3080
rect 12989 3071 13047 3077
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 14550 3000 14556 3052
rect 14608 3040 14614 3052
rect 14737 3043 14795 3049
rect 14737 3040 14749 3043
rect 14608 3012 14749 3040
rect 14608 3000 14614 3012
rect 14737 3009 14749 3012
rect 14783 3009 14795 3043
rect 14737 3003 14795 3009
rect 15013 3043 15071 3049
rect 15013 3009 15025 3043
rect 15059 3040 15071 3043
rect 15562 3040 15568 3052
rect 15059 3012 15568 3040
rect 15059 3009 15071 3012
rect 15013 3003 15071 3009
rect 15562 3000 15568 3012
rect 15620 3000 15626 3052
rect 12805 2975 12863 2981
rect 12805 2941 12817 2975
rect 12851 2941 12863 2975
rect 12805 2935 12863 2941
rect 13354 2932 13360 2984
rect 13412 2972 13418 2984
rect 13541 2975 13599 2981
rect 13541 2972 13553 2975
rect 13412 2944 13553 2972
rect 13412 2932 13418 2944
rect 13541 2941 13553 2944
rect 13587 2941 13599 2975
rect 13541 2935 13599 2941
rect 9217 2867 9275 2873
rect 9324 2876 10456 2904
rect 10980 2876 11928 2904
rect 9324 2836 9352 2876
rect 9582 2836 9588 2848
rect 6288 2808 9352 2836
rect 9543 2808 9588 2836
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 10226 2796 10232 2848
rect 10284 2836 10290 2848
rect 10321 2839 10379 2845
rect 10321 2836 10333 2839
rect 10284 2808 10333 2836
rect 10284 2796 10290 2808
rect 10321 2805 10333 2808
rect 10367 2805 10379 2839
rect 10428 2836 10456 2876
rect 11974 2864 11980 2916
rect 12032 2904 12038 2916
rect 12621 2907 12679 2913
rect 12621 2904 12633 2907
rect 12032 2876 12633 2904
rect 12032 2864 12038 2876
rect 12621 2873 12633 2876
rect 12667 2873 12679 2907
rect 12621 2867 12679 2873
rect 12710 2864 12716 2916
rect 12768 2904 12774 2916
rect 12768 2876 12813 2904
rect 12768 2864 12774 2876
rect 15746 2864 15752 2916
rect 15804 2864 15810 2916
rect 12253 2839 12311 2845
rect 12253 2836 12265 2839
rect 10428 2808 12265 2836
rect 10321 2799 10379 2805
rect 12253 2805 12265 2808
rect 12299 2805 12311 2839
rect 12253 2799 12311 2805
rect 1104 2746 16836 2768
rect 1104 2694 6226 2746
rect 6278 2694 6290 2746
rect 6342 2694 6354 2746
rect 6406 2694 6418 2746
rect 6470 2694 11470 2746
rect 11522 2694 11534 2746
rect 11586 2694 11598 2746
rect 11650 2694 11662 2746
rect 11714 2694 16836 2746
rect 1104 2672 16836 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 3418 2632 3424 2644
rect 1627 2604 3424 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 3786 2592 3792 2644
rect 3844 2632 3850 2644
rect 3881 2635 3939 2641
rect 3881 2632 3893 2635
rect 3844 2604 3893 2632
rect 3844 2592 3850 2604
rect 3881 2601 3893 2604
rect 3927 2601 3939 2635
rect 3881 2595 3939 2601
rect 5261 2635 5319 2641
rect 5261 2601 5273 2635
rect 5307 2632 5319 2635
rect 5718 2632 5724 2644
rect 5307 2604 5724 2632
rect 5307 2601 5319 2604
rect 5261 2595 5319 2601
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2601 6423 2635
rect 6365 2595 6423 2601
rect 7009 2635 7067 2641
rect 7009 2601 7021 2635
rect 7055 2632 7067 2635
rect 7098 2632 7104 2644
rect 7055 2604 7104 2632
rect 7055 2601 7067 2604
rect 7009 2595 7067 2601
rect 4157 2567 4215 2573
rect 4157 2533 4169 2567
rect 4203 2564 4215 2567
rect 4982 2564 4988 2576
rect 4203 2536 4752 2564
rect 4943 2536 4988 2564
rect 4203 2533 4215 2536
rect 4157 2527 4215 2533
rect 4724 2508 4752 2536
rect 4982 2524 4988 2536
rect 5040 2524 5046 2576
rect 6380 2564 6408 2595
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 7374 2592 7380 2644
rect 7432 2632 7438 2644
rect 7834 2632 7840 2644
rect 7432 2604 7840 2632
rect 7432 2592 7438 2604
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8294 2632 8300 2644
rect 8255 2604 8300 2632
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 8680 2604 11284 2632
rect 6733 2567 6791 2573
rect 6733 2564 6745 2567
rect 6380 2536 6745 2564
rect 6733 2533 6745 2536
rect 6779 2533 6791 2567
rect 6733 2527 6791 2533
rect 6822 2524 6828 2576
rect 6880 2564 6886 2576
rect 7469 2567 7527 2573
rect 7469 2564 7481 2567
rect 6880 2536 7481 2564
rect 6880 2524 6886 2536
rect 7469 2533 7481 2536
rect 7515 2533 7527 2567
rect 7469 2527 7527 2533
rect 474 2456 480 2508
rect 532 2496 538 2508
rect 1397 2499 1455 2505
rect 1397 2496 1409 2499
rect 532 2468 1409 2496
rect 532 2456 538 2468
rect 1397 2465 1409 2468
rect 1443 2465 1455 2499
rect 1854 2496 1860 2508
rect 1815 2468 1860 2496
rect 1397 2459 1455 2465
rect 1854 2456 1860 2468
rect 1912 2456 1918 2508
rect 3418 2456 3424 2508
rect 3476 2496 3482 2508
rect 3513 2499 3571 2505
rect 3513 2496 3525 2499
rect 3476 2468 3525 2496
rect 3476 2456 3482 2468
rect 3513 2465 3525 2468
rect 3559 2465 3571 2499
rect 4062 2496 4068 2508
rect 4023 2468 4068 2496
rect 3513 2459 3571 2465
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2465 4307 2499
rect 4430 2496 4436 2508
rect 4391 2468 4436 2496
rect 4249 2459 4307 2465
rect 4264 2428 4292 2459
rect 4430 2456 4436 2468
rect 4488 2456 4494 2508
rect 4706 2496 4712 2508
rect 4667 2468 4712 2496
rect 4706 2456 4712 2468
rect 4764 2456 4770 2508
rect 4801 2499 4859 2505
rect 4801 2465 4813 2499
rect 4847 2465 4859 2499
rect 4801 2459 4859 2465
rect 4614 2428 4620 2440
rect 4264 2400 4620 2428
rect 4614 2388 4620 2400
rect 4672 2428 4678 2440
rect 4816 2428 4844 2459
rect 5074 2456 5080 2508
rect 5132 2496 5138 2508
rect 5721 2499 5779 2505
rect 5132 2468 5177 2496
rect 5132 2456 5138 2468
rect 5721 2465 5733 2499
rect 5767 2465 5779 2499
rect 5721 2459 5779 2465
rect 6089 2499 6147 2505
rect 6089 2465 6101 2499
rect 6135 2496 6147 2499
rect 6181 2499 6239 2505
rect 6181 2496 6193 2499
rect 6135 2468 6193 2496
rect 6135 2465 6147 2468
rect 6089 2459 6147 2465
rect 6181 2465 6193 2468
rect 6227 2465 6239 2499
rect 7377 2499 7435 2505
rect 7377 2496 7389 2499
rect 6181 2459 6239 2465
rect 6932 2468 7389 2496
rect 5736 2428 5764 2459
rect 4672 2400 5764 2428
rect 5813 2431 5871 2437
rect 4672 2388 4678 2400
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 6932 2428 6960 2468
rect 7377 2465 7389 2468
rect 7423 2496 7435 2499
rect 7745 2499 7803 2505
rect 7423 2468 7512 2496
rect 7423 2465 7435 2468
rect 7377 2459 7435 2465
rect 7484 2437 7512 2468
rect 7745 2465 7757 2499
rect 7791 2465 7803 2499
rect 7745 2459 7803 2465
rect 5859 2400 6960 2428
rect 7285 2431 7343 2437
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 7285 2397 7297 2431
rect 7331 2428 7343 2431
rect 7469 2431 7527 2437
rect 7331 2400 7420 2428
rect 7331 2397 7343 2400
rect 7285 2391 7343 2397
rect 4890 2360 4896 2372
rect 2746 2332 4896 2360
rect 2041 2295 2099 2301
rect 2041 2261 2053 2295
rect 2087 2292 2099 2295
rect 2746 2292 2774 2332
rect 4890 2320 4896 2332
rect 4948 2320 4954 2372
rect 4985 2363 5043 2369
rect 4985 2329 4997 2363
rect 5031 2360 5043 2363
rect 5626 2360 5632 2372
rect 5031 2332 5632 2360
rect 5031 2329 5043 2332
rect 4985 2323 5043 2329
rect 5626 2320 5632 2332
rect 5684 2320 5690 2372
rect 6914 2360 6920 2372
rect 6875 2332 6920 2360
rect 6914 2320 6920 2332
rect 6972 2320 6978 2372
rect 7006 2320 7012 2372
rect 7064 2360 7070 2372
rect 7392 2360 7420 2400
rect 7469 2397 7481 2431
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 7760 2428 7788 2459
rect 8294 2456 8300 2508
rect 8352 2496 8358 2508
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 8352 2468 8493 2496
rect 8352 2456 8358 2468
rect 8481 2465 8493 2468
rect 8527 2465 8539 2499
rect 8481 2459 8539 2465
rect 8570 2456 8576 2508
rect 8628 2496 8634 2508
rect 8680 2505 8708 2604
rect 8757 2567 8815 2573
rect 8757 2533 8769 2567
rect 8803 2564 8815 2567
rect 8938 2564 8944 2576
rect 8803 2536 8944 2564
rect 8803 2533 8815 2536
rect 8757 2527 8815 2533
rect 8665 2499 8723 2505
rect 8665 2496 8677 2499
rect 8628 2468 8677 2496
rect 8628 2456 8634 2468
rect 8665 2465 8677 2468
rect 8711 2465 8723 2499
rect 8665 2459 8723 2465
rect 8772 2428 8800 2527
rect 8938 2524 8944 2536
rect 8996 2524 9002 2576
rect 9493 2567 9551 2573
rect 9493 2533 9505 2567
rect 9539 2564 9551 2567
rect 9582 2564 9588 2576
rect 9539 2536 9588 2564
rect 9539 2533 9551 2536
rect 9493 2527 9551 2533
rect 9582 2524 9588 2536
rect 9640 2524 9646 2576
rect 10226 2524 10232 2576
rect 10284 2524 10290 2576
rect 11256 2573 11284 2604
rect 11790 2592 11796 2644
rect 11848 2632 11854 2644
rect 11885 2635 11943 2641
rect 11885 2632 11897 2635
rect 11848 2604 11897 2632
rect 11848 2592 11854 2604
rect 11885 2601 11897 2604
rect 11931 2601 11943 2635
rect 11885 2595 11943 2601
rect 12069 2635 12127 2641
rect 12069 2601 12081 2635
rect 12115 2632 12127 2635
rect 12621 2635 12679 2641
rect 12621 2632 12633 2635
rect 12115 2604 12633 2632
rect 12115 2601 12127 2604
rect 12069 2595 12127 2601
rect 12621 2601 12633 2604
rect 12667 2632 12679 2635
rect 12710 2632 12716 2644
rect 12667 2604 12716 2632
rect 12667 2601 12679 2604
rect 12621 2595 12679 2601
rect 11241 2567 11299 2573
rect 11241 2533 11253 2567
rect 11287 2564 11299 2567
rect 11287 2536 11836 2564
rect 11287 2533 11299 2536
rect 11241 2527 11299 2533
rect 11514 2456 11520 2508
rect 11572 2496 11578 2508
rect 11701 2499 11759 2505
rect 11701 2496 11713 2499
rect 11572 2468 11713 2496
rect 11572 2456 11578 2468
rect 11701 2465 11713 2468
rect 11747 2465 11759 2499
rect 11808 2496 11836 2536
rect 11974 2496 11980 2508
rect 12032 2505 12038 2508
rect 12032 2499 12068 2505
rect 11808 2468 11980 2496
rect 11701 2459 11759 2465
rect 11974 2456 11980 2468
rect 12056 2465 12068 2499
rect 12032 2459 12068 2465
rect 12437 2499 12495 2505
rect 12437 2465 12449 2499
rect 12483 2496 12495 2499
rect 12636 2496 12664 2595
rect 12710 2592 12716 2604
rect 12768 2592 12774 2644
rect 14553 2635 14611 2641
rect 14553 2601 14565 2635
rect 14599 2601 14611 2635
rect 15194 2632 15200 2644
rect 15155 2604 15200 2632
rect 14553 2595 14611 2601
rect 14568 2564 14596 2595
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 15746 2632 15752 2644
rect 15707 2604 15752 2632
rect 15746 2592 15752 2604
rect 15804 2592 15810 2644
rect 16022 2632 16028 2644
rect 15983 2604 16028 2632
rect 16022 2592 16028 2604
rect 16080 2592 16086 2644
rect 13662 2536 14596 2564
rect 14752 2536 15608 2564
rect 12483 2468 12664 2496
rect 14369 2499 14427 2505
rect 12483 2465 12495 2468
rect 12437 2459 12495 2465
rect 14369 2465 14381 2499
rect 14415 2496 14427 2499
rect 14550 2496 14556 2508
rect 14415 2468 14556 2496
rect 14415 2465 14427 2468
rect 14369 2459 14427 2465
rect 12032 2456 12066 2459
rect 14550 2456 14556 2468
rect 14608 2456 14614 2508
rect 14642 2456 14648 2508
rect 14700 2496 14706 2508
rect 14752 2505 14780 2536
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 14700 2468 14749 2496
rect 14700 2456 14706 2468
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 14737 2459 14795 2465
rect 15194 2456 15200 2508
rect 15252 2496 15258 2508
rect 15580 2505 15608 2536
rect 15381 2499 15439 2505
rect 15381 2496 15393 2499
rect 15252 2468 15393 2496
rect 15252 2456 15258 2468
rect 15381 2465 15393 2468
rect 15427 2465 15439 2499
rect 15381 2459 15439 2465
rect 15565 2499 15623 2505
rect 15565 2465 15577 2499
rect 15611 2465 15623 2499
rect 15565 2459 15623 2465
rect 16209 2499 16267 2505
rect 16209 2465 16221 2499
rect 16255 2465 16267 2499
rect 16482 2496 16488 2508
rect 16443 2468 16488 2496
rect 16209 2459 16267 2465
rect 7760 2400 8800 2428
rect 8941 2431 8999 2437
rect 7760 2360 7788 2400
rect 8941 2397 8953 2431
rect 8987 2428 8999 2431
rect 9217 2431 9275 2437
rect 9217 2428 9229 2431
rect 8987 2400 9229 2428
rect 8987 2397 8999 2400
rect 8941 2391 8999 2397
rect 9217 2397 9229 2400
rect 9263 2397 9275 2431
rect 12038 2428 12066 2456
rect 12529 2431 12587 2437
rect 12529 2428 12541 2431
rect 12038 2400 12541 2428
rect 9217 2391 9275 2397
rect 12529 2397 12541 2400
rect 12575 2397 12587 2431
rect 14090 2428 14096 2440
rect 14051 2400 14096 2428
rect 12529 2391 12587 2397
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 16224 2428 16252 2459
rect 16482 2456 16488 2468
rect 16540 2456 16546 2508
rect 16574 2428 16580 2440
rect 16224 2400 16580 2428
rect 16574 2388 16580 2400
rect 16632 2388 16638 2440
rect 7064 2332 7328 2360
rect 7392 2332 7788 2360
rect 7064 2320 7070 2332
rect 2087 2264 2774 2292
rect 3697 2295 3755 2301
rect 2087 2261 2099 2264
rect 2041 2255 2099 2261
rect 3697 2261 3709 2295
rect 3743 2292 3755 2295
rect 3970 2292 3976 2304
rect 3743 2264 3976 2292
rect 3743 2261 3755 2264
rect 3697 2255 3755 2261
rect 3970 2252 3976 2264
rect 4028 2252 4034 2304
rect 6089 2295 6147 2301
rect 6089 2261 6101 2295
rect 6135 2292 6147 2295
rect 7190 2292 7196 2304
rect 6135 2264 7196 2292
rect 6135 2261 6147 2264
rect 6089 2255 6147 2261
rect 7190 2252 7196 2264
rect 7248 2252 7254 2304
rect 7300 2301 7328 2332
rect 8018 2320 8024 2372
rect 8076 2360 8082 2372
rect 8076 2332 9352 2360
rect 8076 2320 8082 2332
rect 7285 2295 7343 2301
rect 7285 2261 7297 2295
rect 7331 2292 7343 2295
rect 7653 2295 7711 2301
rect 7653 2292 7665 2295
rect 7331 2264 7665 2292
rect 7331 2261 7343 2264
rect 7285 2255 7343 2261
rect 7653 2261 7665 2264
rect 7699 2261 7711 2295
rect 7653 2255 7711 2261
rect 7834 2252 7840 2304
rect 7892 2292 7898 2304
rect 8941 2295 8999 2301
rect 8941 2292 8953 2295
rect 7892 2264 8953 2292
rect 7892 2252 7898 2264
rect 8941 2261 8953 2264
rect 8987 2261 8999 2295
rect 9324 2292 9352 2332
rect 15838 2320 15844 2372
rect 15896 2360 15902 2372
rect 16301 2363 16359 2369
rect 16301 2360 16313 2363
rect 15896 2332 16313 2360
rect 15896 2320 15902 2332
rect 16301 2329 16313 2332
rect 16347 2329 16359 2363
rect 16301 2323 16359 2329
rect 11517 2295 11575 2301
rect 11517 2292 11529 2295
rect 9324 2264 11529 2292
rect 8941 2255 8999 2261
rect 11517 2261 11529 2264
rect 11563 2261 11575 2295
rect 11517 2255 11575 2261
rect 1104 2202 16836 2224
rect 1104 2150 3604 2202
rect 3656 2150 3668 2202
rect 3720 2150 3732 2202
rect 3784 2150 3796 2202
rect 3848 2150 8848 2202
rect 8900 2150 8912 2202
rect 8964 2150 8976 2202
rect 9028 2150 9040 2202
rect 9092 2150 14092 2202
rect 14144 2150 14156 2202
rect 14208 2150 14220 2202
rect 14272 2150 14284 2202
rect 14336 2150 16836 2202
rect 1104 2128 16836 2150
rect 3970 2048 3976 2100
rect 4028 2088 4034 2100
rect 7742 2088 7748 2100
rect 4028 2060 7748 2088
rect 4028 2048 4034 2060
rect 7742 2048 7748 2060
rect 7800 2048 7806 2100
<< via1 >>
rect 6226 17926 6278 17978
rect 6290 17926 6342 17978
rect 6354 17926 6406 17978
rect 6418 17926 6470 17978
rect 11470 17926 11522 17978
rect 11534 17926 11586 17978
rect 11598 17926 11650 17978
rect 11662 17926 11714 17978
rect 5080 17824 5132 17876
rect 6920 17799 6972 17808
rect 6920 17765 6929 17799
rect 6929 17765 6963 17799
rect 6963 17765 6972 17799
rect 6920 17756 6972 17765
rect 17040 17756 17092 17808
rect 480 17688 532 17740
rect 2320 17731 2372 17740
rect 2320 17697 2329 17731
rect 2329 17697 2363 17731
rect 2363 17697 2372 17731
rect 2320 17688 2372 17697
rect 3700 17688 3752 17740
rect 5540 17731 5592 17740
rect 5540 17697 5549 17731
rect 5549 17697 5583 17731
rect 5583 17697 5592 17731
rect 5540 17688 5592 17697
rect 6552 17688 6604 17740
rect 8760 17688 8812 17740
rect 10140 17731 10192 17740
rect 10140 17697 10149 17731
rect 10149 17697 10183 17731
rect 10183 17697 10192 17731
rect 10140 17688 10192 17697
rect 11980 17731 12032 17740
rect 11980 17697 11989 17731
rect 11989 17697 12023 17731
rect 12023 17697 12032 17731
rect 11980 17688 12032 17697
rect 13820 17688 13872 17740
rect 15200 17688 15252 17740
rect 16120 17731 16172 17740
rect 16120 17697 16129 17731
rect 16129 17697 16163 17731
rect 16163 17697 16172 17731
rect 16120 17688 16172 17697
rect 4436 17620 4488 17672
rect 12440 17620 12492 17672
rect 4252 17552 4304 17604
rect 1584 17527 1636 17536
rect 1584 17493 1593 17527
rect 1593 17493 1627 17527
rect 1627 17493 1636 17527
rect 1584 17484 1636 17493
rect 3976 17484 4028 17536
rect 4344 17484 4396 17536
rect 4896 17552 4948 17604
rect 5724 17527 5776 17536
rect 5724 17493 5733 17527
rect 5733 17493 5767 17527
rect 5767 17493 5776 17527
rect 5724 17484 5776 17493
rect 8668 17484 8720 17536
rect 12164 17527 12216 17536
rect 12164 17493 12173 17527
rect 12173 17493 12207 17527
rect 12207 17493 12216 17527
rect 12164 17484 12216 17493
rect 15016 17484 15068 17536
rect 15200 17527 15252 17536
rect 15200 17493 15209 17527
rect 15209 17493 15243 17527
rect 15243 17493 15252 17527
rect 15200 17484 15252 17493
rect 15936 17527 15988 17536
rect 15936 17493 15945 17527
rect 15945 17493 15979 17527
rect 15979 17493 15988 17527
rect 15936 17484 15988 17493
rect 3604 17382 3656 17434
rect 3668 17382 3720 17434
rect 3732 17382 3784 17434
rect 3796 17382 3848 17434
rect 8848 17382 8900 17434
rect 8912 17382 8964 17434
rect 8976 17382 9028 17434
rect 9040 17382 9092 17434
rect 14092 17382 14144 17434
rect 14156 17382 14208 17434
rect 14220 17382 14272 17434
rect 14284 17382 14336 17434
rect 4436 17323 4488 17332
rect 4436 17289 4445 17323
rect 4445 17289 4479 17323
rect 4479 17289 4488 17323
rect 4436 17280 4488 17289
rect 5080 17323 5132 17332
rect 5080 17289 5089 17323
rect 5089 17289 5123 17323
rect 5123 17289 5132 17323
rect 5080 17280 5132 17289
rect 6552 17323 6604 17332
rect 6552 17289 6561 17323
rect 6561 17289 6595 17323
rect 6595 17289 6604 17323
rect 6552 17280 6604 17289
rect 2688 17212 2740 17264
rect 4252 17212 4304 17264
rect 3976 17187 4028 17196
rect 1400 17119 1452 17128
rect 1400 17085 1409 17119
rect 1409 17085 1443 17119
rect 1443 17085 1452 17119
rect 1400 17076 1452 17085
rect 3976 17153 3985 17187
rect 3985 17153 4019 17187
rect 4019 17153 4028 17187
rect 3976 17144 4028 17153
rect 4068 17076 4120 17128
rect 5172 17076 5224 17128
rect 10784 17144 10836 17196
rect 15200 17280 15252 17332
rect 12624 17255 12676 17264
rect 12624 17221 12633 17255
rect 12633 17221 12667 17255
rect 12667 17221 12676 17255
rect 12624 17212 12676 17221
rect 6000 17008 6052 17060
rect 7196 17076 7248 17128
rect 8392 17119 8444 17128
rect 8392 17085 8401 17119
rect 8401 17085 8435 17119
rect 8435 17085 8444 17119
rect 8392 17076 8444 17085
rect 12440 17144 12492 17196
rect 13176 17187 13228 17196
rect 13176 17153 13185 17187
rect 13185 17153 13219 17187
rect 13219 17153 13228 17187
rect 13176 17144 13228 17153
rect 8576 17051 8628 17060
rect 8576 17017 8585 17051
rect 8585 17017 8619 17051
rect 8619 17017 8628 17051
rect 8576 17008 8628 17017
rect 9864 17051 9916 17060
rect 9864 17017 9873 17051
rect 9873 17017 9907 17051
rect 9907 17017 9916 17051
rect 10968 17076 11020 17128
rect 9864 17008 9916 17017
rect 5632 16940 5684 16992
rect 10784 17008 10836 17060
rect 10876 16940 10928 16992
rect 11060 17008 11112 17060
rect 12532 17008 12584 17060
rect 12900 17051 12952 17060
rect 12900 17017 12909 17051
rect 12909 17017 12943 17051
rect 12943 17017 12952 17051
rect 12900 17008 12952 17017
rect 15936 17076 15988 17128
rect 12072 16983 12124 16992
rect 12072 16949 12081 16983
rect 12081 16949 12115 16983
rect 12115 16949 12124 16983
rect 12072 16940 12124 16949
rect 6226 16838 6278 16890
rect 6290 16838 6342 16890
rect 6354 16838 6406 16890
rect 6418 16838 6470 16890
rect 11470 16838 11522 16890
rect 11534 16838 11586 16890
rect 11598 16838 11650 16890
rect 11662 16838 11714 16890
rect 4896 16779 4948 16788
rect 4896 16745 4905 16779
rect 4905 16745 4939 16779
rect 4939 16745 4948 16779
rect 4896 16736 4948 16745
rect 5080 16736 5132 16788
rect 6000 16779 6052 16788
rect 6000 16745 6009 16779
rect 6009 16745 6043 16779
rect 6043 16745 6052 16779
rect 6000 16736 6052 16745
rect 10784 16779 10836 16788
rect 10784 16745 10793 16779
rect 10793 16745 10827 16779
rect 10827 16745 10836 16779
rect 10784 16736 10836 16745
rect 8392 16668 8444 16720
rect 5080 16643 5132 16652
rect 5080 16609 5089 16643
rect 5089 16609 5123 16643
rect 5123 16609 5132 16643
rect 5080 16600 5132 16609
rect 5908 16643 5960 16652
rect 5908 16609 5917 16643
rect 5917 16609 5951 16643
rect 5951 16609 5960 16643
rect 5908 16600 5960 16609
rect 6092 16600 6144 16652
rect 7196 16643 7248 16652
rect 7196 16609 7205 16643
rect 7205 16609 7239 16643
rect 7239 16609 7248 16643
rect 7196 16600 7248 16609
rect 8116 16643 8168 16652
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 12624 16668 12676 16720
rect 12532 16600 12584 16652
rect 13360 16643 13412 16652
rect 13360 16609 13369 16643
rect 13369 16609 13403 16643
rect 13403 16609 13412 16643
rect 13360 16600 13412 16609
rect 13820 16532 13872 16584
rect 4712 16439 4764 16448
rect 4712 16405 4721 16439
rect 4721 16405 4755 16439
rect 4755 16405 4764 16439
rect 4712 16396 4764 16405
rect 10692 16439 10744 16448
rect 10692 16405 10701 16439
rect 10701 16405 10735 16439
rect 10735 16405 10744 16439
rect 10692 16396 10744 16405
rect 3604 16294 3656 16346
rect 3668 16294 3720 16346
rect 3732 16294 3784 16346
rect 3796 16294 3848 16346
rect 8848 16294 8900 16346
rect 8912 16294 8964 16346
rect 8976 16294 9028 16346
rect 9040 16294 9092 16346
rect 14092 16294 14144 16346
rect 14156 16294 14208 16346
rect 14220 16294 14272 16346
rect 14284 16294 14336 16346
rect 1584 16056 1636 16108
rect 4068 16192 4120 16244
rect 5632 16235 5684 16244
rect 5632 16201 5641 16235
rect 5641 16201 5675 16235
rect 5675 16201 5684 16235
rect 5632 16192 5684 16201
rect 8116 16192 8168 16244
rect 13820 16235 13872 16244
rect 4712 16124 4764 16176
rect 6828 16056 6880 16108
rect 9496 16124 9548 16176
rect 3976 15988 4028 16040
rect 5080 15988 5132 16040
rect 5632 15988 5684 16040
rect 8576 15988 8628 16040
rect 9496 16031 9548 16040
rect 9496 15997 9505 16031
rect 9505 15997 9539 16031
rect 9539 15997 9548 16031
rect 9496 15988 9548 15997
rect 9864 15988 9916 16040
rect 10692 16124 10744 16176
rect 13820 16201 13829 16235
rect 13829 16201 13863 16235
rect 13863 16201 13872 16235
rect 13820 16192 13872 16201
rect 14924 16124 14976 16176
rect 13360 16056 13412 16108
rect 13452 15988 13504 16040
rect 13912 15988 13964 16040
rect 1768 15895 1820 15904
rect 1768 15861 1777 15895
rect 1777 15861 1811 15895
rect 1811 15861 1820 15895
rect 1768 15852 1820 15861
rect 3240 15852 3292 15904
rect 8116 15852 8168 15904
rect 10508 15895 10560 15904
rect 10508 15861 10517 15895
rect 10517 15861 10551 15895
rect 10551 15861 10560 15895
rect 10508 15852 10560 15861
rect 13728 15895 13780 15904
rect 13728 15861 13737 15895
rect 13737 15861 13771 15895
rect 13771 15861 13780 15895
rect 13728 15852 13780 15861
rect 6226 15750 6278 15802
rect 6290 15750 6342 15802
rect 6354 15750 6406 15802
rect 6418 15750 6470 15802
rect 11470 15750 11522 15802
rect 11534 15750 11586 15802
rect 11598 15750 11650 15802
rect 11662 15750 11714 15802
rect 2504 15648 2556 15700
rect 8576 15648 8628 15700
rect 13728 15648 13780 15700
rect 3240 15623 3292 15632
rect 3240 15589 3249 15623
rect 3249 15589 3283 15623
rect 3283 15589 3292 15623
rect 3240 15580 3292 15589
rect 10508 15580 10560 15632
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 1768 15555 1820 15564
rect 1768 15521 1777 15555
rect 1777 15521 1811 15555
rect 1811 15521 1820 15555
rect 1768 15512 1820 15521
rect 2320 15555 2372 15564
rect 2320 15521 2329 15555
rect 2329 15521 2363 15555
rect 2363 15521 2372 15555
rect 2320 15512 2372 15521
rect 8576 15555 8628 15564
rect 8576 15521 8585 15555
rect 8585 15521 8619 15555
rect 8619 15521 8628 15555
rect 8576 15512 8628 15521
rect 13360 15555 13412 15564
rect 13360 15521 13369 15555
rect 13369 15521 13403 15555
rect 13403 15521 13412 15555
rect 13360 15512 13412 15521
rect 13452 15512 13504 15564
rect 12440 15444 12492 15496
rect 13176 15444 13228 15496
rect 13636 15376 13688 15428
rect 13912 15512 13964 15564
rect 15752 15555 15804 15564
rect 15752 15521 15761 15555
rect 15761 15521 15795 15555
rect 15795 15521 15804 15555
rect 15752 15512 15804 15521
rect 16488 15555 16540 15564
rect 16488 15521 16497 15555
rect 16497 15521 16531 15555
rect 16531 15521 16540 15555
rect 16488 15512 16540 15521
rect 4436 15308 4488 15360
rect 15844 15351 15896 15360
rect 15844 15317 15853 15351
rect 15853 15317 15887 15351
rect 15887 15317 15896 15351
rect 15844 15308 15896 15317
rect 3604 15206 3656 15258
rect 3668 15206 3720 15258
rect 3732 15206 3784 15258
rect 3796 15206 3848 15258
rect 8848 15206 8900 15258
rect 8912 15206 8964 15258
rect 8976 15206 9028 15258
rect 9040 15206 9092 15258
rect 14092 15206 14144 15258
rect 14156 15206 14208 15258
rect 14220 15206 14272 15258
rect 14284 15206 14336 15258
rect 3976 15147 4028 15156
rect 3976 15113 3985 15147
rect 3985 15113 4019 15147
rect 4019 15113 4028 15147
rect 3976 15104 4028 15113
rect 9496 15104 9548 15156
rect 13912 15104 13964 15156
rect 15752 15104 15804 15156
rect 4068 15036 4120 15088
rect 1492 14943 1544 14952
rect 1492 14909 1501 14943
rect 1501 14909 1535 14943
rect 1535 14909 1544 14943
rect 1492 14900 1544 14909
rect 2412 14968 2464 15020
rect 4436 15011 4488 15020
rect 4436 14977 4445 15011
rect 4445 14977 4479 15011
rect 4479 14977 4488 15011
rect 4436 14968 4488 14977
rect 4528 14968 4580 15020
rect 5908 15036 5960 15088
rect 10048 15036 10100 15088
rect 5816 14968 5868 15020
rect 6552 15011 6604 15020
rect 6552 14977 6561 15011
rect 6561 14977 6595 15011
rect 6595 14977 6604 15011
rect 6552 14968 6604 14977
rect 12164 15011 12216 15020
rect 12164 14977 12173 15011
rect 12173 14977 12207 15011
rect 12207 14977 12216 15011
rect 12164 14968 12216 14977
rect 12440 14968 12492 15020
rect 2504 14943 2556 14952
rect 2504 14909 2513 14943
rect 2513 14909 2547 14943
rect 2547 14909 2556 14943
rect 2504 14900 2556 14909
rect 6920 14900 6972 14952
rect 2320 14832 2372 14884
rect 5540 14832 5592 14884
rect 2596 14807 2648 14816
rect 2596 14773 2605 14807
rect 2605 14773 2639 14807
rect 2639 14773 2648 14807
rect 2596 14764 2648 14773
rect 5356 14764 5408 14816
rect 6000 14832 6052 14884
rect 11336 14832 11388 14884
rect 6920 14764 6972 14816
rect 10416 14764 10468 14816
rect 13636 14900 13688 14952
rect 13912 14832 13964 14884
rect 15200 14900 15252 14952
rect 12348 14764 12400 14816
rect 15752 14764 15804 14816
rect 6226 14662 6278 14714
rect 6290 14662 6342 14714
rect 6354 14662 6406 14714
rect 6418 14662 6470 14714
rect 11470 14662 11522 14714
rect 11534 14662 11586 14714
rect 11598 14662 11650 14714
rect 11662 14662 11714 14714
rect 4344 14603 4396 14612
rect 4344 14569 4353 14603
rect 4353 14569 4387 14603
rect 4387 14569 4396 14603
rect 4344 14560 4396 14569
rect 6092 14560 6144 14612
rect 5540 14492 5592 14544
rect 2596 14467 2648 14476
rect 2596 14433 2605 14467
rect 2605 14433 2639 14467
rect 2639 14433 2648 14467
rect 2596 14424 2648 14433
rect 1492 14356 1544 14408
rect 2320 14356 2372 14408
rect 2412 14356 2464 14408
rect 4528 14399 4580 14408
rect 4528 14365 4537 14399
rect 4537 14365 4571 14399
rect 4571 14365 4580 14399
rect 4528 14356 4580 14365
rect 5632 14356 5684 14408
rect 6184 14467 6236 14476
rect 6184 14433 6193 14467
rect 6193 14433 6227 14467
rect 6227 14433 6236 14467
rect 8576 14560 8628 14612
rect 6184 14424 6236 14433
rect 6920 14424 6972 14476
rect 7564 14424 7616 14476
rect 8024 14467 8076 14476
rect 8024 14433 8033 14467
rect 8033 14433 8067 14467
rect 8067 14433 8076 14467
rect 8024 14424 8076 14433
rect 8300 14424 8352 14476
rect 9220 14467 9272 14476
rect 9220 14433 9229 14467
rect 9229 14433 9263 14467
rect 9263 14433 9272 14467
rect 9220 14424 9272 14433
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 10416 14467 10468 14476
rect 10416 14433 10425 14467
rect 10425 14433 10459 14467
rect 10459 14433 10468 14467
rect 10416 14424 10468 14433
rect 11888 14467 11940 14476
rect 6000 14331 6052 14340
rect 6000 14297 6009 14331
rect 6009 14297 6043 14331
rect 6043 14297 6052 14331
rect 6000 14288 6052 14297
rect 6644 14399 6696 14408
rect 6644 14365 6653 14399
rect 6653 14365 6687 14399
rect 6687 14365 6696 14399
rect 6644 14356 6696 14365
rect 3148 14220 3200 14272
rect 5908 14220 5960 14272
rect 6920 14288 6972 14340
rect 10600 14263 10652 14272
rect 10600 14229 10609 14263
rect 10609 14229 10643 14263
rect 10643 14229 10652 14263
rect 10600 14220 10652 14229
rect 11888 14433 11897 14467
rect 11897 14433 11931 14467
rect 11931 14433 11940 14467
rect 11888 14424 11940 14433
rect 11336 14356 11388 14408
rect 16488 14467 16540 14476
rect 16488 14433 16497 14467
rect 16497 14433 16531 14467
rect 16531 14433 16540 14467
rect 16488 14424 16540 14433
rect 16304 14263 16356 14272
rect 16304 14229 16313 14263
rect 16313 14229 16347 14263
rect 16347 14229 16356 14263
rect 16304 14220 16356 14229
rect 3604 14118 3656 14170
rect 3668 14118 3720 14170
rect 3732 14118 3784 14170
rect 3796 14118 3848 14170
rect 8848 14118 8900 14170
rect 8912 14118 8964 14170
rect 8976 14118 9028 14170
rect 9040 14118 9092 14170
rect 14092 14118 14144 14170
rect 14156 14118 14208 14170
rect 14220 14118 14272 14170
rect 14284 14118 14336 14170
rect 9220 14016 9272 14068
rect 13912 14016 13964 14068
rect 14832 14016 14884 14068
rect 8208 13948 8260 14000
rect 13728 13948 13780 14000
rect 5632 13812 5684 13864
rect 7288 13855 7340 13864
rect 7288 13821 7297 13855
rect 7297 13821 7331 13855
rect 7331 13821 7340 13855
rect 7288 13812 7340 13821
rect 8024 13812 8076 13864
rect 10600 13812 10652 13864
rect 11796 13855 11848 13864
rect 11796 13821 11805 13855
rect 11805 13821 11839 13855
rect 11839 13821 11848 13855
rect 11796 13812 11848 13821
rect 12072 13812 12124 13864
rect 13728 13855 13780 13864
rect 13728 13821 13737 13855
rect 13737 13821 13771 13855
rect 13771 13821 13780 13855
rect 14096 13855 14148 13864
rect 13728 13812 13780 13821
rect 14096 13821 14105 13855
rect 14105 13821 14139 13855
rect 14139 13821 14148 13855
rect 14096 13812 14148 13821
rect 15844 13948 15896 14000
rect 15384 13812 15436 13864
rect 14832 13744 14884 13796
rect 4252 13676 4304 13728
rect 4804 13719 4856 13728
rect 4804 13685 4813 13719
rect 4813 13685 4847 13719
rect 4847 13685 4856 13719
rect 8300 13719 8352 13728
rect 4804 13676 4856 13685
rect 8300 13685 8309 13719
rect 8309 13685 8343 13719
rect 8343 13685 8352 13719
rect 8300 13676 8352 13685
rect 12072 13719 12124 13728
rect 12072 13685 12081 13719
rect 12081 13685 12115 13719
rect 12115 13685 12124 13719
rect 12072 13676 12124 13685
rect 6226 13574 6278 13626
rect 6290 13574 6342 13626
rect 6354 13574 6406 13626
rect 6418 13574 6470 13626
rect 11470 13574 11522 13626
rect 11534 13574 11586 13626
rect 11598 13574 11650 13626
rect 11662 13574 11714 13626
rect 5724 13472 5776 13524
rect 8668 13515 8720 13524
rect 8668 13481 8677 13515
rect 8677 13481 8711 13515
rect 8711 13481 8720 13515
rect 8668 13472 8720 13481
rect 11888 13472 11940 13524
rect 12072 13472 12124 13524
rect 14096 13515 14148 13524
rect 14096 13481 14105 13515
rect 14105 13481 14139 13515
rect 14139 13481 14148 13515
rect 14096 13472 14148 13481
rect 4252 13404 4304 13456
rect 2412 13379 2464 13388
rect 2412 13345 2421 13379
rect 2421 13345 2455 13379
rect 2455 13345 2464 13379
rect 2412 13336 2464 13345
rect 3884 13379 3936 13388
rect 3884 13345 3893 13379
rect 3893 13345 3927 13379
rect 3927 13345 3936 13379
rect 3884 13336 3936 13345
rect 10508 13404 10560 13456
rect 16212 13404 16264 13456
rect 5172 13379 5224 13388
rect 5172 13345 5181 13379
rect 5181 13345 5215 13379
rect 5215 13345 5224 13379
rect 5172 13336 5224 13345
rect 6460 13336 6512 13388
rect 8576 13379 8628 13388
rect 8576 13345 8585 13379
rect 8585 13345 8619 13379
rect 8619 13345 8628 13379
rect 8576 13336 8628 13345
rect 9864 13336 9916 13388
rect 10600 13379 10652 13388
rect 10600 13345 10609 13379
rect 10609 13345 10643 13379
rect 10643 13345 10652 13379
rect 10600 13336 10652 13345
rect 13912 13336 13964 13388
rect 6000 13311 6052 13320
rect 6000 13277 6009 13311
rect 6009 13277 6043 13311
rect 6043 13277 6052 13311
rect 6000 13268 6052 13277
rect 6552 13268 6604 13320
rect 8668 13268 8720 13320
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 10784 13200 10836 13252
rect 12440 13268 12492 13320
rect 15108 13268 15160 13320
rect 3240 13132 3292 13184
rect 4436 13132 4488 13184
rect 10140 13175 10192 13184
rect 10140 13141 10149 13175
rect 10149 13141 10183 13175
rect 10183 13141 10192 13175
rect 10140 13132 10192 13141
rect 3604 13030 3656 13082
rect 3668 13030 3720 13082
rect 3732 13030 3784 13082
rect 3796 13030 3848 13082
rect 8848 13030 8900 13082
rect 8912 13030 8964 13082
rect 8976 13030 9028 13082
rect 9040 13030 9092 13082
rect 14092 13030 14144 13082
rect 14156 13030 14208 13082
rect 14220 13030 14272 13082
rect 14284 13030 14336 13082
rect 6460 12971 6512 12980
rect 6460 12937 6469 12971
rect 6469 12937 6503 12971
rect 6503 12937 6512 12971
rect 6460 12928 6512 12937
rect 6552 12928 6604 12980
rect 6828 12928 6880 12980
rect 7196 12928 7248 12980
rect 7564 12971 7616 12980
rect 4804 12903 4856 12912
rect 4804 12869 4813 12903
rect 4813 12869 4847 12903
rect 4847 12869 4856 12903
rect 4804 12860 4856 12869
rect 7564 12937 7573 12971
rect 7573 12937 7607 12971
rect 7607 12937 7616 12971
rect 7564 12928 7616 12937
rect 8576 12928 8628 12980
rect 8484 12860 8536 12912
rect 11796 12928 11848 12980
rect 13912 12928 13964 12980
rect 15384 12971 15436 12980
rect 12164 12860 12216 12912
rect 2780 12792 2832 12844
rect 3148 12792 3200 12844
rect 4436 12835 4488 12844
rect 3240 12767 3292 12776
rect 3240 12733 3249 12767
rect 3249 12733 3283 12767
rect 3283 12733 3292 12767
rect 3240 12724 3292 12733
rect 3976 12724 4028 12776
rect 4436 12801 4445 12835
rect 4445 12801 4479 12835
rect 4479 12801 4488 12835
rect 4436 12792 4488 12801
rect 5908 12792 5960 12844
rect 6644 12835 6696 12844
rect 6644 12801 6653 12835
rect 6653 12801 6687 12835
rect 6687 12801 6696 12835
rect 6644 12792 6696 12801
rect 7104 12792 7156 12844
rect 8668 12792 8720 12844
rect 10140 12792 10192 12844
rect 6736 12767 6788 12776
rect 6736 12733 6745 12767
rect 6745 12733 6779 12767
rect 6779 12733 6788 12767
rect 6920 12767 6972 12776
rect 6736 12724 6788 12733
rect 6920 12733 6929 12767
rect 6929 12733 6963 12767
rect 6963 12733 6972 12767
rect 6920 12724 6972 12733
rect 8208 12724 8260 12776
rect 10784 12767 10836 12776
rect 10784 12733 10793 12767
rect 10793 12733 10827 12767
rect 10827 12733 10836 12767
rect 10784 12724 10836 12733
rect 10876 12767 10928 12776
rect 10876 12733 10885 12767
rect 10885 12733 10919 12767
rect 10919 12733 10928 12767
rect 11336 12792 11388 12844
rect 12808 12792 12860 12844
rect 15384 12937 15393 12971
rect 15393 12937 15427 12971
rect 15427 12937 15436 12971
rect 15384 12928 15436 12937
rect 10876 12724 10928 12733
rect 2228 12656 2280 12708
rect 6092 12656 6144 12708
rect 7380 12656 7432 12708
rect 4988 12588 5040 12640
rect 6920 12588 6972 12640
rect 8300 12656 8352 12708
rect 14004 12767 14056 12776
rect 7840 12588 7892 12640
rect 8024 12631 8076 12640
rect 8024 12597 8033 12631
rect 8033 12597 8067 12631
rect 8067 12597 8076 12631
rect 8024 12588 8076 12597
rect 10324 12588 10376 12640
rect 11336 12656 11388 12708
rect 14004 12733 14013 12767
rect 14013 12733 14047 12767
rect 14047 12733 14056 12767
rect 14004 12724 14056 12733
rect 11244 12588 11296 12640
rect 11796 12588 11848 12640
rect 15108 12792 15160 12844
rect 14280 12724 14332 12776
rect 14832 12724 14884 12776
rect 16304 12724 16356 12776
rect 15752 12631 15804 12640
rect 15752 12597 15761 12631
rect 15761 12597 15795 12631
rect 15795 12597 15804 12631
rect 15752 12588 15804 12597
rect 6226 12486 6278 12538
rect 6290 12486 6342 12538
rect 6354 12486 6406 12538
rect 6418 12486 6470 12538
rect 11470 12486 11522 12538
rect 11534 12486 11586 12538
rect 11598 12486 11650 12538
rect 11662 12486 11714 12538
rect 7196 12384 7248 12436
rect 9864 12427 9916 12436
rect 9864 12393 9873 12427
rect 9873 12393 9907 12427
rect 9907 12393 9916 12427
rect 10600 12427 10652 12436
rect 9864 12384 9916 12393
rect 10600 12393 10609 12427
rect 10609 12393 10643 12427
rect 10643 12393 10652 12427
rect 10600 12384 10652 12393
rect 11336 12427 11388 12436
rect 2136 12316 2188 12368
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 2780 12248 2832 12300
rect 5356 12248 5408 12300
rect 6736 12248 6788 12300
rect 7104 12248 7156 12300
rect 7840 12291 7892 12300
rect 6920 12180 6972 12232
rect 7196 12180 7248 12232
rect 7840 12257 7849 12291
rect 7849 12257 7883 12291
rect 7883 12257 7892 12291
rect 7840 12248 7892 12257
rect 8484 12316 8536 12368
rect 10232 12316 10284 12368
rect 1584 12155 1636 12164
rect 1584 12121 1593 12155
rect 1593 12121 1627 12155
rect 1627 12121 1636 12155
rect 1584 12112 1636 12121
rect 8300 12223 8352 12232
rect 8300 12189 8309 12223
rect 8309 12189 8343 12223
rect 8343 12189 8352 12223
rect 8300 12180 8352 12189
rect 8392 12180 8444 12232
rect 9680 12180 9732 12232
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10324 12291 10376 12300
rect 10048 12248 10100 12257
rect 10324 12257 10333 12291
rect 10333 12257 10367 12291
rect 10367 12257 10376 12291
rect 10324 12248 10376 12257
rect 10876 12316 10928 12368
rect 10784 12291 10836 12300
rect 10784 12257 10793 12291
rect 10793 12257 10827 12291
rect 10827 12257 10836 12291
rect 10784 12248 10836 12257
rect 11152 12248 11204 12300
rect 11336 12393 11345 12427
rect 11345 12393 11379 12427
rect 11379 12393 11388 12427
rect 11336 12384 11388 12393
rect 11980 12427 12032 12436
rect 11980 12393 11989 12427
rect 11989 12393 12023 12427
rect 12023 12393 12032 12427
rect 11980 12384 12032 12393
rect 12072 12384 12124 12436
rect 12348 12384 12400 12436
rect 15752 12384 15804 12436
rect 10876 12223 10928 12232
rect 10876 12189 10885 12223
rect 10885 12189 10919 12223
rect 10919 12189 10928 12223
rect 10876 12180 10928 12189
rect 13176 12316 13228 12368
rect 14832 12316 14884 12368
rect 11796 12291 11848 12300
rect 11796 12257 11805 12291
rect 11805 12257 11839 12291
rect 11839 12257 11848 12291
rect 11796 12248 11848 12257
rect 11980 12291 12032 12300
rect 11980 12257 11989 12291
rect 11989 12257 12023 12291
rect 12023 12257 12032 12291
rect 11980 12248 12032 12257
rect 12072 12248 12124 12300
rect 12808 12291 12860 12300
rect 12808 12257 12817 12291
rect 12817 12257 12851 12291
rect 12851 12257 12860 12291
rect 12808 12248 12860 12257
rect 15568 12248 15620 12300
rect 9404 12112 9456 12164
rect 9496 12112 9548 12164
rect 10232 12155 10284 12164
rect 10232 12121 10241 12155
rect 10241 12121 10275 12155
rect 10275 12121 10284 12155
rect 10232 12112 10284 12121
rect 11152 12112 11204 12164
rect 13268 12180 13320 12232
rect 11980 12112 12032 12164
rect 14556 12112 14608 12164
rect 1768 12087 1820 12096
rect 1768 12053 1777 12087
rect 1777 12053 1811 12087
rect 1811 12053 1820 12087
rect 1768 12044 1820 12053
rect 6092 12044 6144 12096
rect 6184 12087 6236 12096
rect 6184 12053 6193 12087
rect 6193 12053 6227 12087
rect 6227 12053 6236 12087
rect 6184 12044 6236 12053
rect 7656 12044 7708 12096
rect 7932 12087 7984 12096
rect 7932 12053 7941 12087
rect 7941 12053 7975 12087
rect 7975 12053 7984 12087
rect 7932 12044 7984 12053
rect 8208 12044 8260 12096
rect 12348 12044 12400 12096
rect 13820 12044 13872 12096
rect 3604 11942 3656 11994
rect 3668 11942 3720 11994
rect 3732 11942 3784 11994
rect 3796 11942 3848 11994
rect 8848 11942 8900 11994
rect 8912 11942 8964 11994
rect 8976 11942 9028 11994
rect 9040 11942 9092 11994
rect 14092 11942 14144 11994
rect 14156 11942 14208 11994
rect 14220 11942 14272 11994
rect 14284 11942 14336 11994
rect 7932 11840 7984 11892
rect 6644 11815 6696 11824
rect 6644 11781 6653 11815
rect 6653 11781 6687 11815
rect 6687 11781 6696 11815
rect 6644 11772 6696 11781
rect 8852 11772 8904 11824
rect 8944 11772 8996 11824
rect 9772 11840 9824 11892
rect 10140 11840 10192 11892
rect 12256 11840 12308 11892
rect 12900 11840 12952 11892
rect 8576 11704 8628 11756
rect 1768 11636 1820 11688
rect 2412 11636 2464 11688
rect 4988 11679 5040 11688
rect 4988 11645 4997 11679
rect 4997 11645 5031 11679
rect 5031 11645 5040 11679
rect 4988 11636 5040 11645
rect 6552 11679 6604 11688
rect 6552 11645 6561 11679
rect 6561 11645 6595 11679
rect 6595 11645 6604 11679
rect 6552 11636 6604 11645
rect 6736 11679 6788 11688
rect 6736 11645 6745 11679
rect 6745 11645 6779 11679
rect 6779 11645 6788 11679
rect 6736 11636 6788 11645
rect 7196 11636 7248 11688
rect 8484 11636 8536 11688
rect 9864 11772 9916 11824
rect 12440 11772 12492 11824
rect 13268 11840 13320 11892
rect 13728 11883 13780 11892
rect 13728 11849 13737 11883
rect 13737 11849 13771 11883
rect 13771 11849 13780 11883
rect 13728 11840 13780 11849
rect 15200 11840 15252 11892
rect 13084 11772 13136 11824
rect 11152 11704 11204 11756
rect 2228 11611 2280 11620
rect 2228 11577 2237 11611
rect 2237 11577 2271 11611
rect 2271 11577 2280 11611
rect 2228 11568 2280 11577
rect 7656 11568 7708 11620
rect 10692 11636 10744 11688
rect 11980 11704 12032 11756
rect 12808 11704 12860 11756
rect 12072 11679 12124 11688
rect 12072 11645 12081 11679
rect 12081 11645 12115 11679
rect 12115 11645 12124 11679
rect 12072 11636 12124 11645
rect 12256 11679 12308 11688
rect 12256 11645 12265 11679
rect 12265 11645 12299 11679
rect 12299 11645 12308 11679
rect 12256 11636 12308 11645
rect 12440 11636 12492 11688
rect 12716 11636 12768 11688
rect 13268 11636 13320 11688
rect 14280 11704 14332 11756
rect 15108 11704 15160 11756
rect 14832 11679 14884 11688
rect 14832 11645 14841 11679
rect 14841 11645 14875 11679
rect 14875 11645 14884 11679
rect 14832 11636 14884 11645
rect 15752 11679 15804 11688
rect 15752 11645 15761 11679
rect 15761 11645 15795 11679
rect 15795 11645 15804 11679
rect 15752 11636 15804 11645
rect 9680 11568 9732 11620
rect 14556 11611 14608 11620
rect 14556 11577 14565 11611
rect 14565 11577 14599 11611
rect 14599 11577 14608 11611
rect 14556 11568 14608 11577
rect 4344 11500 4396 11552
rect 9220 11500 9272 11552
rect 14004 11500 14056 11552
rect 14096 11543 14148 11552
rect 14096 11509 14105 11543
rect 14105 11509 14139 11543
rect 14139 11509 14148 11543
rect 14096 11500 14148 11509
rect 14280 11500 14332 11552
rect 15752 11500 15804 11552
rect 16028 11500 16080 11552
rect 6226 11398 6278 11450
rect 6290 11398 6342 11450
rect 6354 11398 6406 11450
rect 6418 11398 6470 11450
rect 11470 11398 11522 11450
rect 11534 11398 11586 11450
rect 11598 11398 11650 11450
rect 11662 11398 11714 11450
rect 3332 11228 3384 11280
rect 5080 11296 5132 11348
rect 7840 11296 7892 11348
rect 1584 11203 1636 11212
rect 1584 11169 1593 11203
rect 1593 11169 1627 11203
rect 1627 11169 1636 11203
rect 1584 11160 1636 11169
rect 2688 11160 2740 11212
rect 4344 11160 4396 11212
rect 7748 11203 7800 11212
rect 2136 11024 2188 11076
rect 2320 11024 2372 11076
rect 3148 11092 3200 11144
rect 7748 11169 7757 11203
rect 7757 11169 7791 11203
rect 7791 11169 7800 11203
rect 7748 11160 7800 11169
rect 8300 11160 8352 11212
rect 9036 11228 9088 11280
rect 8668 11160 8720 11212
rect 8944 11203 8996 11212
rect 8944 11169 8953 11203
rect 8953 11169 8987 11203
rect 8987 11169 8996 11203
rect 8944 11160 8996 11169
rect 9220 11296 9272 11348
rect 9588 11228 9640 11280
rect 10876 11296 10928 11348
rect 13360 11296 13412 11348
rect 16212 11296 16264 11348
rect 9680 11160 9732 11212
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 10416 11160 10468 11212
rect 11152 11203 11204 11212
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 11152 11169 11161 11203
rect 11161 11169 11195 11203
rect 11195 11169 11204 11203
rect 11152 11160 11204 11169
rect 11428 11203 11480 11212
rect 11428 11169 11442 11203
rect 11442 11169 11476 11203
rect 11476 11169 11480 11203
rect 11428 11160 11480 11169
rect 11520 11135 11572 11144
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 13268 11228 13320 11280
rect 15844 11228 15896 11280
rect 13176 11203 13228 11212
rect 13176 11169 13185 11203
rect 13185 11169 13219 11203
rect 13219 11169 13228 11203
rect 13176 11160 13228 11169
rect 11520 11092 11572 11101
rect 12348 11092 12400 11144
rect 13820 11160 13872 11212
rect 14556 11203 14608 11212
rect 7472 11024 7524 11076
rect 8392 11024 8444 11076
rect 9772 11024 9824 11076
rect 11428 11024 11480 11076
rect 11796 11067 11848 11076
rect 11796 11033 11805 11067
rect 11805 11033 11839 11067
rect 11839 11033 11848 11067
rect 11796 11024 11848 11033
rect 11980 11024 12032 11076
rect 14556 11169 14565 11203
rect 14565 11169 14599 11203
rect 14599 11169 14608 11203
rect 14556 11160 14608 11169
rect 15108 11160 15160 11212
rect 16488 11203 16540 11212
rect 16488 11169 16497 11203
rect 16497 11169 16531 11203
rect 16531 11169 16540 11203
rect 16488 11160 16540 11169
rect 14924 11067 14976 11076
rect 14924 11033 14933 11067
rect 14933 11033 14967 11067
rect 14967 11033 14976 11067
rect 14924 11024 14976 11033
rect 6460 10956 6512 11008
rect 8208 10999 8260 11008
rect 8208 10965 8217 10999
rect 8217 10965 8251 10999
rect 8251 10965 8260 10999
rect 8208 10956 8260 10965
rect 8484 10956 8536 11008
rect 11612 10999 11664 11008
rect 11612 10965 11621 10999
rect 11621 10965 11655 10999
rect 11655 10965 11664 10999
rect 11612 10956 11664 10965
rect 13268 10999 13320 11008
rect 13268 10965 13277 10999
rect 13277 10965 13311 10999
rect 13311 10965 13320 10999
rect 13268 10956 13320 10965
rect 3604 10854 3656 10906
rect 3668 10854 3720 10906
rect 3732 10854 3784 10906
rect 3796 10854 3848 10906
rect 8848 10854 8900 10906
rect 8912 10854 8964 10906
rect 8976 10854 9028 10906
rect 9040 10854 9092 10906
rect 14092 10854 14144 10906
rect 14156 10854 14208 10906
rect 14220 10854 14272 10906
rect 14284 10854 14336 10906
rect 6460 10795 6512 10804
rect 6460 10761 6469 10795
rect 6469 10761 6503 10795
rect 6503 10761 6512 10795
rect 6460 10752 6512 10761
rect 6644 10752 6696 10804
rect 6920 10795 6972 10804
rect 6920 10761 6929 10795
rect 6929 10761 6963 10795
rect 6963 10761 6972 10795
rect 7288 10795 7340 10804
rect 6920 10752 6972 10761
rect 7288 10761 7297 10795
rect 7297 10761 7331 10795
rect 7331 10761 7340 10795
rect 7288 10752 7340 10761
rect 7748 10752 7800 10804
rect 9220 10752 9272 10804
rect 3148 10659 3200 10668
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 4804 10684 4856 10736
rect 6000 10684 6052 10736
rect 8668 10684 8720 10736
rect 10140 10752 10192 10804
rect 11152 10752 11204 10804
rect 11612 10752 11664 10804
rect 12348 10752 12400 10804
rect 2136 10548 2188 10600
rect 2780 10591 2832 10600
rect 2780 10557 2789 10591
rect 2789 10557 2823 10591
rect 2823 10557 2832 10591
rect 6552 10616 6604 10668
rect 7932 10659 7984 10668
rect 7932 10625 7941 10659
rect 7941 10625 7975 10659
rect 7975 10625 7984 10659
rect 7932 10616 7984 10625
rect 8392 10659 8444 10668
rect 8392 10625 8401 10659
rect 8401 10625 8435 10659
rect 8435 10625 8444 10659
rect 9588 10684 9640 10736
rect 10232 10727 10284 10736
rect 10232 10693 10241 10727
rect 10241 10693 10275 10727
rect 10275 10693 10284 10727
rect 10232 10684 10284 10693
rect 8392 10616 8444 10625
rect 8852 10616 8904 10668
rect 11520 10684 11572 10736
rect 11704 10727 11756 10736
rect 11704 10693 11713 10727
rect 11713 10693 11747 10727
rect 11747 10693 11756 10727
rect 11704 10684 11756 10693
rect 10416 10616 10468 10668
rect 2780 10548 2832 10557
rect 4344 10591 4396 10600
rect 4344 10557 4353 10591
rect 4353 10557 4387 10591
rect 4387 10557 4396 10591
rect 4344 10548 4396 10557
rect 5080 10591 5132 10600
rect 5080 10557 5089 10591
rect 5089 10557 5123 10591
rect 5123 10557 5132 10591
rect 5080 10548 5132 10557
rect 2228 10480 2280 10532
rect 3240 10455 3292 10464
rect 3240 10421 3249 10455
rect 3249 10421 3283 10455
rect 3283 10421 3292 10455
rect 3240 10412 3292 10421
rect 6000 10591 6052 10600
rect 6000 10557 6009 10591
rect 6009 10557 6043 10591
rect 6043 10557 6052 10591
rect 6184 10591 6236 10600
rect 6000 10548 6052 10557
rect 6184 10557 6193 10591
rect 6193 10557 6227 10591
rect 6227 10557 6236 10591
rect 6184 10548 6236 10557
rect 7012 10591 7064 10600
rect 7012 10557 7021 10591
rect 7021 10557 7055 10591
rect 7055 10557 7064 10591
rect 7012 10548 7064 10557
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 8208 10548 8260 10600
rect 8576 10591 8628 10600
rect 8576 10557 8585 10591
rect 8585 10557 8619 10591
rect 8619 10557 8628 10591
rect 8576 10548 8628 10557
rect 9036 10548 9088 10600
rect 9220 10591 9272 10600
rect 9220 10557 9229 10591
rect 9229 10557 9263 10591
rect 9263 10557 9272 10591
rect 9220 10548 9272 10557
rect 9680 10591 9732 10600
rect 8484 10480 8536 10532
rect 9680 10557 9689 10591
rect 9689 10557 9723 10591
rect 9723 10557 9732 10591
rect 9680 10548 9732 10557
rect 9864 10548 9916 10600
rect 10876 10616 10928 10668
rect 11152 10591 11204 10600
rect 11152 10557 11161 10591
rect 11161 10557 11195 10591
rect 11195 10557 11204 10591
rect 11152 10548 11204 10557
rect 11428 10591 11480 10600
rect 11428 10557 11437 10591
rect 11437 10557 11471 10591
rect 11471 10557 11480 10591
rect 11428 10548 11480 10557
rect 12256 10616 12308 10668
rect 12440 10591 12492 10600
rect 4804 10455 4856 10464
rect 4804 10421 4813 10455
rect 4813 10421 4847 10455
rect 4847 10421 4856 10455
rect 4804 10412 4856 10421
rect 5540 10412 5592 10464
rect 6644 10412 6696 10464
rect 7748 10455 7800 10464
rect 7748 10421 7757 10455
rect 7757 10421 7791 10455
rect 7791 10421 7800 10455
rect 7748 10412 7800 10421
rect 9496 10480 9548 10532
rect 10692 10480 10744 10532
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12440 10548 12492 10557
rect 14464 10659 14516 10668
rect 14464 10625 14473 10659
rect 14473 10625 14507 10659
rect 14507 10625 14516 10659
rect 14464 10616 14516 10625
rect 12716 10548 12768 10600
rect 13084 10548 13136 10600
rect 13360 10548 13412 10600
rect 14648 10548 14700 10600
rect 15660 10591 15712 10600
rect 15660 10557 15669 10591
rect 15669 10557 15703 10591
rect 15703 10557 15712 10591
rect 15660 10548 15712 10557
rect 11152 10412 11204 10464
rect 11336 10455 11388 10464
rect 11336 10421 11345 10455
rect 11345 10421 11379 10455
rect 11379 10421 11388 10455
rect 11336 10412 11388 10421
rect 14924 10412 14976 10464
rect 15936 10412 15988 10464
rect 6226 10310 6278 10362
rect 6290 10310 6342 10362
rect 6354 10310 6406 10362
rect 6418 10310 6470 10362
rect 11470 10310 11522 10362
rect 11534 10310 11586 10362
rect 11598 10310 11650 10362
rect 11662 10310 11714 10362
rect 3240 10208 3292 10260
rect 6000 10208 6052 10260
rect 6736 10208 6788 10260
rect 7012 10208 7064 10260
rect 10232 10208 10284 10260
rect 6644 10140 6696 10192
rect 10784 10140 10836 10192
rect 11336 10140 11388 10192
rect 14924 10183 14976 10192
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 2136 10115 2188 10124
rect 2136 10081 2145 10115
rect 2145 10081 2179 10115
rect 2179 10081 2188 10115
rect 2136 10072 2188 10081
rect 3148 10072 3200 10124
rect 6552 10072 6604 10124
rect 12348 10072 12400 10124
rect 13360 10072 13412 10124
rect 2320 10047 2372 10056
rect 2320 10013 2329 10047
rect 2329 10013 2363 10047
rect 2363 10013 2372 10047
rect 2320 10004 2372 10013
rect 12716 10047 12768 10056
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 13084 10004 13136 10056
rect 13820 10115 13872 10124
rect 13820 10081 13829 10115
rect 13829 10081 13863 10115
rect 13863 10081 13872 10115
rect 14924 10149 14933 10183
rect 14933 10149 14967 10183
rect 14967 10149 14976 10183
rect 14924 10140 14976 10149
rect 15936 10140 15988 10192
rect 13820 10072 13872 10081
rect 14556 10072 14608 10124
rect 11060 9936 11112 9988
rect 12256 9936 12308 9988
rect 13912 9936 13964 9988
rect 12532 9911 12584 9920
rect 12532 9877 12541 9911
rect 12541 9877 12575 9911
rect 12575 9877 12584 9911
rect 12532 9868 12584 9877
rect 13820 9868 13872 9920
rect 14924 10004 14976 10056
rect 3604 9766 3656 9818
rect 3668 9766 3720 9818
rect 3732 9766 3784 9818
rect 3796 9766 3848 9818
rect 8848 9766 8900 9818
rect 8912 9766 8964 9818
rect 8976 9766 9028 9818
rect 9040 9766 9092 9818
rect 14092 9766 14144 9818
rect 14156 9766 14208 9818
rect 14220 9766 14272 9818
rect 14284 9766 14336 9818
rect 5632 9596 5684 9648
rect 7840 9596 7892 9648
rect 11244 9639 11296 9648
rect 11244 9605 11253 9639
rect 11253 9605 11287 9639
rect 11287 9605 11296 9639
rect 11244 9596 11296 9605
rect 2780 9528 2832 9580
rect 2228 9503 2280 9512
rect 2228 9469 2237 9503
rect 2237 9469 2271 9503
rect 2271 9469 2280 9503
rect 2228 9460 2280 9469
rect 3608 9460 3660 9512
rect 3884 9503 3936 9512
rect 3884 9469 3893 9503
rect 3893 9469 3927 9503
rect 3927 9469 3936 9503
rect 3884 9460 3936 9469
rect 4712 9528 4764 9580
rect 7104 9528 7156 9580
rect 10968 9528 11020 9580
rect 5540 9460 5592 9512
rect 10048 9503 10100 9512
rect 10048 9469 10057 9503
rect 10057 9469 10091 9503
rect 10091 9469 10100 9503
rect 10048 9460 10100 9469
rect 10876 9503 10928 9512
rect 4804 9392 4856 9444
rect 6828 9392 6880 9444
rect 7012 9392 7064 9444
rect 9588 9392 9640 9444
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 10876 9460 10928 9469
rect 2044 9367 2096 9376
rect 2044 9333 2053 9367
rect 2053 9333 2087 9367
rect 2087 9333 2096 9367
rect 2044 9324 2096 9333
rect 4344 9324 4396 9376
rect 9772 9324 9824 9376
rect 10416 9324 10468 9376
rect 11060 9392 11112 9444
rect 11796 9460 11848 9512
rect 11888 9460 11940 9512
rect 12532 9664 12584 9716
rect 12716 9664 12768 9716
rect 14464 9707 14516 9716
rect 14464 9673 14473 9707
rect 14473 9673 14507 9707
rect 14507 9673 14516 9707
rect 14464 9664 14516 9673
rect 12348 9596 12400 9648
rect 13084 9596 13136 9648
rect 13820 9596 13872 9648
rect 12348 9503 12400 9512
rect 12348 9469 12357 9503
rect 12357 9469 12391 9503
rect 12391 9469 12400 9503
rect 12348 9460 12400 9469
rect 12072 9392 12124 9444
rect 11336 9324 11388 9376
rect 13176 9528 13228 9580
rect 13084 9503 13136 9512
rect 13084 9469 13093 9503
rect 13093 9469 13127 9503
rect 13127 9469 13136 9503
rect 13084 9460 13136 9469
rect 13268 9503 13320 9512
rect 13268 9469 13277 9503
rect 13277 9469 13311 9503
rect 13311 9469 13320 9503
rect 13268 9460 13320 9469
rect 13360 9392 13412 9444
rect 13636 9460 13688 9512
rect 13912 9503 13964 9512
rect 13912 9469 13922 9503
rect 13922 9469 13956 9503
rect 13956 9469 13964 9503
rect 13912 9460 13964 9469
rect 14464 9460 14516 9512
rect 15568 9503 15620 9512
rect 15568 9469 15577 9503
rect 15577 9469 15611 9503
rect 15611 9469 15620 9503
rect 15568 9460 15620 9469
rect 14556 9324 14608 9376
rect 15660 9324 15712 9376
rect 6226 9222 6278 9274
rect 6290 9222 6342 9274
rect 6354 9222 6406 9274
rect 6418 9222 6470 9274
rect 11470 9222 11522 9274
rect 11534 9222 11586 9274
rect 11598 9222 11650 9274
rect 11662 9222 11714 9274
rect 3608 9163 3660 9172
rect 3608 9129 3617 9163
rect 3617 9129 3651 9163
rect 3651 9129 3660 9163
rect 3608 9120 3660 9129
rect 3884 9120 3936 9172
rect 5540 9120 5592 9172
rect 6092 9120 6144 9172
rect 7012 9163 7064 9172
rect 7012 9129 7021 9163
rect 7021 9129 7055 9163
rect 7055 9129 7064 9163
rect 7012 9120 7064 9129
rect 3148 9052 3200 9104
rect 2044 9027 2096 9036
rect 2044 8993 2053 9027
rect 2053 8993 2087 9027
rect 2087 8993 2096 9027
rect 2044 8984 2096 8993
rect 4344 9095 4396 9104
rect 4344 9061 4353 9095
rect 4353 9061 4387 9095
rect 4387 9061 4396 9095
rect 4344 9052 4396 9061
rect 5632 9052 5684 9104
rect 9220 9120 9272 9172
rect 9588 9120 9640 9172
rect 4712 9027 4764 9036
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 4712 8993 4721 9027
rect 4721 8993 4755 9027
rect 4755 8993 4764 9027
rect 4712 8984 4764 8993
rect 5540 9027 5592 9036
rect 5540 8993 5549 9027
rect 5549 8993 5583 9027
rect 5583 8993 5592 9027
rect 5540 8984 5592 8993
rect 4896 8916 4948 8968
rect 6736 8984 6788 9036
rect 8484 8984 8536 9036
rect 2596 8780 2648 8832
rect 6552 8916 6604 8968
rect 7104 8959 7156 8968
rect 7104 8925 7113 8959
rect 7113 8925 7147 8959
rect 7147 8925 7156 8959
rect 7104 8916 7156 8925
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 10324 9027 10376 9036
rect 10324 8993 10333 9027
rect 10333 8993 10367 9027
rect 10367 8993 10376 9027
rect 10324 8984 10376 8993
rect 11796 9120 11848 9172
rect 11244 9052 11296 9104
rect 10784 9027 10836 9036
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 10784 8984 10836 8993
rect 11336 9027 11388 9036
rect 9772 8848 9824 8900
rect 10232 8848 10284 8900
rect 11336 8993 11345 9027
rect 11345 8993 11379 9027
rect 11379 8993 11388 9027
rect 12072 9052 12124 9104
rect 12624 9052 12676 9104
rect 14648 9120 14700 9172
rect 16304 9120 16356 9172
rect 12808 9095 12860 9104
rect 12808 9061 12817 9095
rect 12817 9061 12851 9095
rect 12851 9061 12860 9095
rect 12808 9052 12860 9061
rect 15660 9052 15712 9104
rect 11336 8984 11388 8993
rect 13176 9027 13228 9036
rect 13176 8993 13185 9027
rect 13185 8993 13219 9027
rect 13219 8993 13228 9027
rect 13176 8984 13228 8993
rect 13360 9027 13412 9036
rect 13360 8993 13369 9027
rect 13369 8993 13403 9027
rect 13403 8993 13412 9027
rect 13360 8984 13412 8993
rect 14924 8916 14976 8968
rect 13636 8848 13688 8900
rect 8576 8780 8628 8832
rect 9680 8823 9732 8832
rect 9680 8789 9689 8823
rect 9689 8789 9723 8823
rect 9723 8789 9732 8823
rect 9680 8780 9732 8789
rect 3604 8678 3656 8730
rect 3668 8678 3720 8730
rect 3732 8678 3784 8730
rect 3796 8678 3848 8730
rect 8848 8678 8900 8730
rect 8912 8678 8964 8730
rect 8976 8678 9028 8730
rect 9040 8678 9092 8730
rect 14092 8678 14144 8730
rect 14156 8678 14208 8730
rect 14220 8678 14272 8730
rect 14284 8678 14336 8730
rect 4896 8619 4948 8628
rect 4896 8585 4905 8619
rect 4905 8585 4939 8619
rect 4939 8585 4948 8619
rect 4896 8576 4948 8585
rect 6828 8619 6880 8628
rect 6828 8585 6837 8619
rect 6837 8585 6871 8619
rect 6871 8585 6880 8619
rect 6828 8576 6880 8585
rect 8484 8619 8536 8628
rect 8484 8585 8493 8619
rect 8493 8585 8527 8619
rect 8527 8585 8536 8619
rect 8484 8576 8536 8585
rect 10324 8576 10376 8628
rect 4344 8372 4396 8424
rect 7840 8440 7892 8492
rect 9680 8508 9732 8560
rect 8576 8440 8628 8492
rect 10416 8483 10468 8492
rect 8668 8415 8720 8424
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 11336 8440 11388 8492
rect 13176 8372 13228 8424
rect 13912 8415 13964 8424
rect 13912 8381 13921 8415
rect 13921 8381 13955 8415
rect 13955 8381 13964 8415
rect 13912 8372 13964 8381
rect 16488 8415 16540 8424
rect 16488 8381 16497 8415
rect 16497 8381 16531 8415
rect 16531 8381 16540 8415
rect 16488 8372 16540 8381
rect 10232 8304 10284 8356
rect 13820 8236 13872 8288
rect 16304 8279 16356 8288
rect 16304 8245 16313 8279
rect 16313 8245 16347 8279
rect 16347 8245 16356 8279
rect 16304 8236 16356 8245
rect 6226 8134 6278 8186
rect 6290 8134 6342 8186
rect 6354 8134 6406 8186
rect 6418 8134 6470 8186
rect 11470 8134 11522 8186
rect 11534 8134 11586 8186
rect 11598 8134 11650 8186
rect 11662 8134 11714 8186
rect 3148 8032 3200 8084
rect 11336 8032 11388 8084
rect 12348 8032 12400 8084
rect 13084 8032 13136 8084
rect 13728 8032 13780 8084
rect 13912 8032 13964 8084
rect 11244 7964 11296 8016
rect 13452 7964 13504 8016
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 2320 7939 2372 7948
rect 2320 7905 2329 7939
rect 2329 7905 2363 7939
rect 2363 7905 2372 7939
rect 2320 7896 2372 7905
rect 2964 7939 3016 7948
rect 2964 7905 2973 7939
rect 2973 7905 3007 7939
rect 3007 7905 3016 7939
rect 2964 7896 3016 7905
rect 4160 7896 4212 7948
rect 6092 7896 6144 7948
rect 6736 7896 6788 7948
rect 8668 7896 8720 7948
rect 11888 7939 11940 7948
rect 11888 7905 11897 7939
rect 11897 7905 11931 7939
rect 11931 7905 11940 7939
rect 11888 7896 11940 7905
rect 12624 7896 12676 7948
rect 12532 7828 12584 7880
rect 12256 7760 12308 7812
rect 13728 7896 13780 7948
rect 14556 7896 14608 7948
rect 15016 7896 15068 7948
rect 15660 7939 15712 7948
rect 15660 7905 15669 7939
rect 15669 7905 15703 7939
rect 15703 7905 15712 7939
rect 15660 7896 15712 7905
rect 14832 7828 14884 7880
rect 2412 7692 2464 7744
rect 2688 7692 2740 7744
rect 6828 7735 6880 7744
rect 6828 7701 6837 7735
rect 6837 7701 6871 7735
rect 6871 7701 6880 7735
rect 6828 7692 6880 7701
rect 9220 7692 9272 7744
rect 12348 7692 12400 7744
rect 16396 7760 16448 7812
rect 14556 7692 14608 7744
rect 14832 7692 14884 7744
rect 15108 7692 15160 7744
rect 15936 7692 15988 7744
rect 3604 7590 3656 7642
rect 3668 7590 3720 7642
rect 3732 7590 3784 7642
rect 3796 7590 3848 7642
rect 8848 7590 8900 7642
rect 8912 7590 8964 7642
rect 8976 7590 9028 7642
rect 9040 7590 9092 7642
rect 14092 7590 14144 7642
rect 14156 7590 14208 7642
rect 14220 7590 14272 7642
rect 14284 7590 14336 7642
rect 3424 7488 3476 7540
rect 4436 7488 4488 7540
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 11980 7488 12032 7540
rect 12532 7531 12584 7540
rect 2688 7352 2740 7404
rect 2964 7352 3016 7404
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 3424 7327 3476 7336
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 4068 7327 4120 7336
rect 4068 7293 4077 7327
rect 4077 7293 4111 7327
rect 4111 7293 4120 7327
rect 4068 7284 4120 7293
rect 2412 7216 2464 7268
rect 3516 7259 3568 7268
rect 3516 7225 3525 7259
rect 3525 7225 3559 7259
rect 3559 7225 3568 7259
rect 3516 7216 3568 7225
rect 4436 7327 4488 7336
rect 4436 7293 4445 7327
rect 4445 7293 4479 7327
rect 4479 7293 4488 7327
rect 4436 7284 4488 7293
rect 7932 7420 7984 7472
rect 9772 7352 9824 7404
rect 6092 7284 6144 7336
rect 3240 7191 3292 7200
rect 3240 7157 3249 7191
rect 3249 7157 3283 7191
rect 3283 7157 3292 7191
rect 5724 7216 5776 7268
rect 3240 7148 3292 7157
rect 4344 7148 4396 7200
rect 4712 7191 4764 7200
rect 4712 7157 4721 7191
rect 4721 7157 4755 7191
rect 4755 7157 4764 7191
rect 4712 7148 4764 7157
rect 5264 7148 5316 7200
rect 10232 7284 10284 7336
rect 10784 7327 10836 7336
rect 10784 7293 10793 7327
rect 10793 7293 10827 7327
rect 10827 7293 10836 7327
rect 10784 7284 10836 7293
rect 10968 7327 11020 7336
rect 10968 7293 10977 7327
rect 10977 7293 11011 7327
rect 11011 7293 11020 7327
rect 10968 7284 11020 7293
rect 11244 7327 11296 7336
rect 11244 7293 11253 7327
rect 11253 7293 11287 7327
rect 11287 7293 11296 7327
rect 11244 7284 11296 7293
rect 12256 7352 12308 7404
rect 12532 7497 12541 7531
rect 12541 7497 12575 7531
rect 12575 7497 12584 7531
rect 12532 7488 12584 7497
rect 13452 7488 13504 7540
rect 14648 7488 14700 7540
rect 16396 7531 16448 7540
rect 16396 7497 16405 7531
rect 16405 7497 16439 7531
rect 16439 7497 16448 7531
rect 16396 7488 16448 7497
rect 12348 7284 12400 7336
rect 13820 7352 13872 7404
rect 13912 7352 13964 7404
rect 12624 7327 12676 7336
rect 12624 7293 12633 7327
rect 12633 7293 12667 7327
rect 12667 7293 12676 7327
rect 13544 7327 13596 7336
rect 12624 7284 12676 7293
rect 13544 7293 13553 7327
rect 13553 7293 13587 7327
rect 13587 7293 13596 7327
rect 13544 7284 13596 7293
rect 6736 7259 6788 7268
rect 6736 7225 6745 7259
rect 6745 7225 6779 7259
rect 6779 7225 6788 7259
rect 6736 7216 6788 7225
rect 6828 7216 6880 7268
rect 9220 7216 9272 7268
rect 9864 7259 9916 7268
rect 9864 7225 9873 7259
rect 9873 7225 9907 7259
rect 9907 7225 9916 7259
rect 9864 7216 9916 7225
rect 10324 7259 10376 7268
rect 10324 7225 10333 7259
rect 10333 7225 10367 7259
rect 10367 7225 10376 7259
rect 10324 7216 10376 7225
rect 11980 7216 12032 7268
rect 7104 7148 7156 7200
rect 7472 7148 7524 7200
rect 8208 7148 8260 7200
rect 14372 7284 14424 7336
rect 14924 7352 14976 7404
rect 12440 7148 12492 7200
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 15936 7216 15988 7268
rect 15016 7148 15068 7200
rect 6226 7046 6278 7098
rect 6290 7046 6342 7098
rect 6354 7046 6406 7098
rect 6418 7046 6470 7098
rect 11470 7046 11522 7098
rect 11534 7046 11586 7098
rect 11598 7046 11650 7098
rect 11662 7046 11714 7098
rect 3516 6944 3568 6996
rect 5724 6987 5776 6996
rect 5724 6953 5733 6987
rect 5733 6953 5767 6987
rect 5767 6953 5776 6987
rect 5724 6944 5776 6953
rect 2504 6876 2556 6928
rect 5264 6876 5316 6928
rect 6644 6876 6696 6928
rect 7932 6919 7984 6928
rect 7932 6885 7941 6919
rect 7941 6885 7975 6919
rect 7975 6885 7984 6919
rect 7932 6876 7984 6885
rect 8208 6944 8260 6996
rect 1400 6740 1452 6792
rect 3240 6740 3292 6792
rect 2780 6672 2832 6724
rect 1492 6604 1544 6656
rect 4344 6740 4396 6792
rect 4712 6740 4764 6792
rect 5264 6740 5316 6792
rect 6920 6808 6972 6860
rect 6736 6672 6788 6724
rect 7196 6672 7248 6724
rect 10324 6808 10376 6860
rect 13544 6944 13596 6996
rect 12440 6876 12492 6928
rect 11888 6808 11940 6860
rect 12900 6808 12952 6860
rect 13360 6808 13412 6860
rect 9864 6672 9916 6724
rect 7472 6604 7524 6656
rect 12532 6740 12584 6792
rect 13452 6740 13504 6792
rect 15292 6808 15344 6860
rect 11520 6604 11572 6656
rect 11888 6672 11940 6724
rect 14648 6740 14700 6792
rect 12256 6604 12308 6656
rect 13820 6604 13872 6656
rect 3604 6502 3656 6554
rect 3668 6502 3720 6554
rect 3732 6502 3784 6554
rect 3796 6502 3848 6554
rect 8848 6502 8900 6554
rect 8912 6502 8964 6554
rect 8976 6502 9028 6554
rect 9040 6502 9092 6554
rect 14092 6502 14144 6554
rect 14156 6502 14208 6554
rect 14220 6502 14272 6554
rect 14284 6502 14336 6554
rect 2504 6443 2556 6452
rect 2504 6409 2513 6443
rect 2513 6409 2547 6443
rect 2547 6409 2556 6443
rect 2504 6400 2556 6409
rect 10784 6400 10836 6452
rect 8208 6332 8260 6384
rect 2596 6196 2648 6248
rect 3424 6196 3476 6248
rect 4068 6196 4120 6248
rect 7012 6196 7064 6248
rect 7840 6196 7892 6248
rect 8208 6239 8260 6248
rect 8208 6205 8217 6239
rect 8217 6205 8251 6239
rect 8251 6205 8260 6239
rect 8208 6196 8260 6205
rect 12532 6400 12584 6452
rect 13360 6443 13412 6452
rect 13360 6409 13369 6443
rect 13369 6409 13403 6443
rect 13403 6409 13412 6443
rect 13360 6400 13412 6409
rect 15292 6443 15344 6452
rect 15292 6409 15301 6443
rect 15301 6409 15335 6443
rect 15335 6409 15344 6443
rect 15292 6400 15344 6409
rect 15752 6400 15804 6452
rect 13452 6332 13504 6384
rect 11980 6307 12032 6316
rect 11980 6273 11989 6307
rect 11989 6273 12023 6307
rect 12023 6273 12032 6307
rect 11980 6264 12032 6273
rect 12900 6264 12952 6316
rect 13820 6307 13872 6316
rect 13820 6273 13829 6307
rect 13829 6273 13863 6307
rect 13863 6273 13872 6307
rect 13820 6264 13872 6273
rect 14464 6264 14516 6316
rect 15660 6264 15712 6316
rect 7196 6128 7248 6180
rect 8392 6171 8444 6180
rect 8392 6137 8401 6171
rect 8401 6137 8435 6171
rect 8435 6137 8444 6171
rect 9772 6196 9824 6248
rect 10324 6239 10376 6248
rect 8392 6128 8444 6137
rect 5264 6103 5316 6112
rect 5264 6069 5273 6103
rect 5273 6069 5307 6103
rect 5307 6069 5316 6103
rect 5264 6060 5316 6069
rect 6644 6060 6696 6112
rect 7564 6060 7616 6112
rect 8484 6060 8536 6112
rect 8852 6103 8904 6112
rect 8852 6069 8861 6103
rect 8861 6069 8895 6103
rect 8895 6069 8904 6103
rect 8852 6060 8904 6069
rect 10324 6205 10333 6239
rect 10333 6205 10367 6239
rect 10367 6205 10376 6239
rect 10324 6196 10376 6205
rect 10508 6239 10560 6248
rect 10508 6205 10517 6239
rect 10517 6205 10551 6239
rect 10551 6205 10560 6239
rect 10508 6196 10560 6205
rect 10968 6239 11020 6248
rect 10968 6205 10977 6239
rect 10977 6205 11011 6239
rect 11011 6205 11020 6239
rect 10968 6196 11020 6205
rect 12164 6196 12216 6248
rect 13452 6239 13504 6248
rect 13452 6205 13461 6239
rect 13461 6205 13495 6239
rect 13495 6205 13504 6239
rect 13452 6196 13504 6205
rect 16488 6239 16540 6248
rect 12348 6060 12400 6112
rect 16488 6205 16497 6239
rect 16497 6205 16531 6239
rect 16531 6205 16540 6239
rect 16488 6196 16540 6205
rect 14556 6128 14608 6180
rect 13820 6060 13872 6112
rect 14832 6060 14884 6112
rect 15936 6103 15988 6112
rect 15936 6069 15945 6103
rect 15945 6069 15979 6103
rect 15979 6069 15988 6103
rect 15936 6060 15988 6069
rect 6226 5958 6278 6010
rect 6290 5958 6342 6010
rect 6354 5958 6406 6010
rect 6418 5958 6470 6010
rect 11470 5958 11522 6010
rect 11534 5958 11586 6010
rect 11598 5958 11650 6010
rect 11662 5958 11714 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 4160 5856 4212 5908
rect 5264 5856 5316 5908
rect 7472 5856 7524 5908
rect 10232 5856 10284 5908
rect 12900 5856 12952 5908
rect 14556 5856 14608 5908
rect 14832 5856 14884 5908
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 6368 5788 6420 5840
rect 3424 5652 3476 5704
rect 4252 5720 4304 5772
rect 7380 5763 7432 5772
rect 7380 5729 7389 5763
rect 7389 5729 7423 5763
rect 7423 5729 7432 5763
rect 10508 5788 10560 5840
rect 12256 5831 12308 5840
rect 12256 5797 12265 5831
rect 12265 5797 12299 5831
rect 12299 5797 12308 5831
rect 12256 5788 12308 5797
rect 13268 5788 13320 5840
rect 15936 5788 15988 5840
rect 16304 5788 16356 5840
rect 7380 5720 7432 5729
rect 8852 5720 8904 5772
rect 10140 5763 10192 5772
rect 4620 5652 4672 5704
rect 7104 5695 7156 5704
rect 7104 5661 7113 5695
rect 7113 5661 7147 5695
rect 7147 5661 7156 5695
rect 7104 5652 7156 5661
rect 7564 5652 7616 5704
rect 8392 5652 8444 5704
rect 9220 5584 9272 5636
rect 10140 5729 10149 5763
rect 10149 5729 10183 5763
rect 10183 5729 10192 5763
rect 10140 5720 10192 5729
rect 14464 5763 14516 5772
rect 14464 5729 14473 5763
rect 14473 5729 14507 5763
rect 14507 5729 14516 5763
rect 14464 5720 14516 5729
rect 9956 5695 10008 5704
rect 9956 5661 9965 5695
rect 9965 5661 9999 5695
rect 9999 5661 10008 5695
rect 9956 5652 10008 5661
rect 10232 5652 10284 5704
rect 13820 5652 13872 5704
rect 3148 5559 3200 5568
rect 3148 5525 3157 5559
rect 3157 5525 3191 5559
rect 3191 5525 3200 5559
rect 3148 5516 3200 5525
rect 4160 5559 4212 5568
rect 4160 5525 4169 5559
rect 4169 5525 4203 5559
rect 4203 5525 4212 5559
rect 4160 5516 4212 5525
rect 5448 5516 5500 5568
rect 14832 5516 14884 5568
rect 3604 5414 3656 5466
rect 3668 5414 3720 5466
rect 3732 5414 3784 5466
rect 3796 5414 3848 5466
rect 8848 5414 8900 5466
rect 8912 5414 8964 5466
rect 8976 5414 9028 5466
rect 9040 5414 9092 5466
rect 14092 5414 14144 5466
rect 14156 5414 14208 5466
rect 14220 5414 14272 5466
rect 14284 5414 14336 5466
rect 6368 5312 6420 5364
rect 7104 5312 7156 5364
rect 10140 5312 10192 5364
rect 13268 5312 13320 5364
rect 4344 5244 4396 5296
rect 1492 5176 1544 5228
rect 3148 5176 3200 5228
rect 4160 5176 4212 5228
rect 6920 5219 6972 5228
rect 4620 5108 4672 5160
rect 6920 5185 6929 5219
rect 6929 5185 6963 5219
rect 6963 5185 6972 5219
rect 6920 5176 6972 5185
rect 6092 5151 6144 5160
rect 2596 5040 2648 5092
rect 6092 5117 6101 5151
rect 6101 5117 6135 5151
rect 6135 5117 6144 5151
rect 6092 5108 6144 5117
rect 7012 5151 7064 5160
rect 5448 5040 5500 5092
rect 7012 5117 7021 5151
rect 7021 5117 7055 5151
rect 7055 5117 7064 5151
rect 7012 5108 7064 5117
rect 7196 5151 7248 5160
rect 7196 5117 7205 5151
rect 7205 5117 7239 5151
rect 7239 5117 7248 5151
rect 7196 5108 7248 5117
rect 7288 5151 7340 5160
rect 7288 5117 7297 5151
rect 7297 5117 7331 5151
rect 7331 5117 7340 5151
rect 7288 5108 7340 5117
rect 8484 5176 8536 5228
rect 9220 5176 9272 5228
rect 9680 5151 9732 5160
rect 4252 5015 4304 5024
rect 4252 4981 4261 5015
rect 4261 4981 4295 5015
rect 4295 4981 4304 5015
rect 4252 4972 4304 4981
rect 4528 5015 4580 5024
rect 4528 4981 4537 5015
rect 4537 4981 4571 5015
rect 4571 4981 4580 5015
rect 4528 4972 4580 4981
rect 4712 4972 4764 5024
rect 7104 5040 7156 5092
rect 9680 5117 9689 5151
rect 9689 5117 9723 5151
rect 9723 5117 9732 5151
rect 9680 5108 9732 5117
rect 9864 5151 9916 5160
rect 9864 5117 9873 5151
rect 9873 5117 9907 5151
rect 9907 5117 9916 5151
rect 9864 5108 9916 5117
rect 10232 5151 10284 5160
rect 10232 5117 10241 5151
rect 10241 5117 10275 5151
rect 10275 5117 10284 5151
rect 10232 5108 10284 5117
rect 10508 5151 10560 5160
rect 10508 5117 10517 5151
rect 10517 5117 10551 5151
rect 10551 5117 10560 5151
rect 10508 5108 10560 5117
rect 11336 5108 11388 5160
rect 11888 5151 11940 5160
rect 11888 5117 11897 5151
rect 11897 5117 11931 5151
rect 11931 5117 11940 5151
rect 11888 5108 11940 5117
rect 12992 5151 13044 5160
rect 10968 5040 11020 5092
rect 11244 5083 11296 5092
rect 11244 5049 11253 5083
rect 11253 5049 11287 5083
rect 11287 5049 11296 5083
rect 11244 5040 11296 5049
rect 12072 5040 12124 5092
rect 12992 5117 13001 5151
rect 13001 5117 13035 5151
rect 13035 5117 13044 5151
rect 12992 5108 13044 5117
rect 6920 4972 6972 5024
rect 7288 4972 7340 5024
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 12716 4972 12768 5024
rect 6226 4870 6278 4922
rect 6290 4870 6342 4922
rect 6354 4870 6406 4922
rect 6418 4870 6470 4922
rect 11470 4870 11522 4922
rect 11534 4870 11586 4922
rect 11598 4870 11650 4922
rect 11662 4870 11714 4922
rect 5540 4768 5592 4820
rect 9864 4768 9916 4820
rect 11244 4768 11296 4820
rect 4344 4675 4396 4684
rect 4344 4641 4353 4675
rect 4353 4641 4387 4675
rect 4387 4641 4396 4675
rect 4344 4632 4396 4641
rect 4528 4632 4580 4684
rect 5724 4632 5776 4684
rect 6000 4675 6052 4684
rect 6000 4641 6009 4675
rect 6009 4641 6043 4675
rect 6043 4641 6052 4675
rect 6000 4632 6052 4641
rect 6184 4675 6236 4684
rect 6184 4641 6193 4675
rect 6193 4641 6227 4675
rect 6227 4641 6236 4675
rect 6184 4632 6236 4641
rect 9220 4675 9272 4684
rect 9220 4641 9229 4675
rect 9229 4641 9263 4675
rect 9263 4641 9272 4675
rect 9220 4632 9272 4641
rect 9404 4675 9456 4684
rect 9404 4641 9413 4675
rect 9413 4641 9447 4675
rect 9447 4641 9456 4675
rect 9404 4632 9456 4641
rect 10324 4700 10376 4752
rect 10232 4632 10284 4684
rect 5724 4496 5776 4548
rect 10508 4632 10560 4684
rect 11244 4675 11296 4684
rect 11244 4641 11253 4675
rect 11253 4641 11287 4675
rect 11287 4641 11296 4675
rect 11244 4632 11296 4641
rect 11796 4675 11848 4684
rect 11796 4641 11805 4675
rect 11805 4641 11839 4675
rect 11839 4641 11848 4675
rect 11796 4632 11848 4641
rect 12072 4632 12124 4684
rect 14740 4700 14792 4752
rect 12716 4675 12768 4684
rect 11336 4564 11388 4616
rect 12440 4607 12492 4616
rect 12440 4573 12449 4607
rect 12449 4573 12483 4607
rect 12483 4573 12492 4607
rect 12440 4564 12492 4573
rect 11888 4496 11940 4548
rect 12716 4641 12725 4675
rect 12725 4641 12759 4675
rect 12759 4641 12768 4675
rect 12716 4632 12768 4641
rect 12992 4632 13044 4684
rect 14464 4632 14516 4684
rect 16488 4675 16540 4684
rect 16488 4641 16497 4675
rect 16497 4641 16531 4675
rect 16531 4641 16540 4675
rect 16488 4632 16540 4641
rect 5080 4428 5132 4480
rect 6000 4428 6052 4480
rect 9404 4428 9456 4480
rect 9956 4428 10008 4480
rect 15200 4496 15252 4548
rect 13820 4471 13872 4480
rect 13820 4437 13829 4471
rect 13829 4437 13863 4471
rect 13863 4437 13872 4471
rect 13820 4428 13872 4437
rect 15568 4428 15620 4480
rect 3604 4326 3656 4378
rect 3668 4326 3720 4378
rect 3732 4326 3784 4378
rect 3796 4326 3848 4378
rect 8848 4326 8900 4378
rect 8912 4326 8964 4378
rect 8976 4326 9028 4378
rect 9040 4326 9092 4378
rect 14092 4326 14144 4378
rect 14156 4326 14208 4378
rect 14220 4326 14272 4378
rect 14284 4326 14336 4378
rect 6184 4224 6236 4276
rect 4896 4088 4948 4140
rect 5632 4156 5684 4208
rect 5724 4199 5776 4208
rect 5724 4165 5733 4199
rect 5733 4165 5767 4199
rect 5767 4165 5776 4199
rect 9680 4224 9732 4276
rect 10140 4224 10192 4276
rect 12992 4224 13044 4276
rect 14832 4267 14884 4276
rect 14832 4233 14862 4267
rect 14862 4233 14884 4267
rect 14832 4224 14884 4233
rect 5724 4156 5776 4165
rect 12440 4156 12492 4208
rect 5080 4063 5132 4072
rect 5080 4029 5089 4063
rect 5089 4029 5123 4063
rect 5123 4029 5132 4063
rect 5080 4020 5132 4029
rect 7012 4088 7064 4140
rect 5632 4063 5684 4072
rect 1584 3952 1636 4004
rect 5632 4029 5641 4063
rect 5641 4029 5675 4063
rect 5675 4029 5684 4063
rect 5632 4020 5684 4029
rect 6644 4063 6696 4072
rect 6644 4029 6653 4063
rect 6653 4029 6687 4063
rect 6687 4029 6696 4063
rect 6644 4020 6696 4029
rect 6736 4063 6788 4072
rect 6736 4029 6745 4063
rect 6745 4029 6779 4063
rect 6779 4029 6788 4063
rect 13728 4088 13780 4140
rect 14556 4131 14608 4140
rect 14556 4097 14565 4131
rect 14565 4097 14599 4131
rect 14599 4097 14608 4131
rect 14556 4088 14608 4097
rect 6736 4020 6788 4029
rect 7380 4063 7432 4072
rect 7380 4029 7389 4063
rect 7389 4029 7423 4063
rect 7423 4029 7432 4063
rect 7380 4020 7432 4029
rect 11244 4063 11296 4072
rect 11244 4029 11253 4063
rect 11253 4029 11287 4063
rect 11287 4029 11296 4063
rect 11244 4020 11296 4029
rect 12072 4063 12124 4072
rect 12072 4029 12081 4063
rect 12081 4029 12115 4063
rect 12115 4029 12124 4063
rect 12072 4020 12124 4029
rect 6828 3952 6880 4004
rect 4436 3884 4488 3936
rect 5264 3884 5316 3936
rect 6644 3884 6696 3936
rect 7104 3884 7156 3936
rect 8668 3952 8720 4004
rect 10048 3884 10100 3936
rect 12440 4063 12492 4072
rect 12440 4029 12449 4063
rect 12449 4029 12483 4063
rect 12483 4029 12492 4063
rect 12440 4020 12492 4029
rect 12348 3995 12400 4004
rect 12348 3961 12357 3995
rect 12357 3961 12391 3995
rect 12391 3961 12400 3995
rect 12348 3952 12400 3961
rect 15568 3952 15620 4004
rect 13820 3884 13872 3936
rect 14464 3927 14516 3936
rect 14464 3893 14473 3927
rect 14473 3893 14507 3927
rect 14507 3893 14516 3927
rect 14464 3884 14516 3893
rect 16396 3884 16448 3936
rect 6226 3782 6278 3834
rect 6290 3782 6342 3834
rect 6354 3782 6406 3834
rect 6418 3782 6470 3834
rect 11470 3782 11522 3834
rect 11534 3782 11586 3834
rect 11598 3782 11650 3834
rect 11662 3782 11714 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 4344 3680 4396 3732
rect 5172 3680 5224 3732
rect 7012 3680 7064 3732
rect 8668 3680 8720 3732
rect 11888 3680 11940 3732
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 2596 3544 2648 3596
rect 6092 3612 6144 3664
rect 3424 3544 3476 3596
rect 4620 3544 4672 3596
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 6920 3587 6972 3596
rect 4988 3476 5040 3528
rect 4620 3408 4672 3460
rect 6920 3553 6929 3587
rect 6929 3553 6963 3587
rect 6963 3553 6972 3587
rect 6920 3544 6972 3553
rect 7104 3587 7156 3596
rect 7104 3553 7113 3587
rect 7113 3553 7147 3587
rect 7147 3553 7156 3587
rect 7104 3544 7156 3553
rect 7196 3544 7248 3596
rect 10140 3544 10192 3596
rect 12348 3612 12400 3664
rect 11152 3544 11204 3596
rect 6644 3476 6696 3528
rect 7288 3408 7340 3460
rect 9404 3408 9456 3460
rect 11244 3408 11296 3460
rect 14464 3544 14516 3596
rect 15568 3587 15620 3596
rect 15568 3553 15577 3587
rect 15577 3553 15611 3587
rect 15611 3553 15620 3587
rect 15568 3544 15620 3553
rect 16304 3587 16356 3596
rect 16304 3553 16313 3587
rect 16313 3553 16347 3587
rect 16347 3553 16356 3587
rect 16304 3544 16356 3553
rect 16396 3519 16448 3528
rect 16396 3485 16405 3519
rect 16405 3485 16439 3519
rect 16439 3485 16448 3519
rect 16396 3476 16448 3485
rect 12164 3408 12216 3460
rect 15568 3408 15620 3460
rect 2412 3340 2464 3392
rect 4252 3340 4304 3392
rect 6184 3340 6236 3392
rect 8392 3340 8444 3392
rect 12440 3340 12492 3392
rect 3604 3238 3656 3290
rect 3668 3238 3720 3290
rect 3732 3238 3784 3290
rect 3796 3238 3848 3290
rect 8848 3238 8900 3290
rect 8912 3238 8964 3290
rect 8976 3238 9028 3290
rect 9040 3238 9092 3290
rect 14092 3238 14144 3290
rect 14156 3238 14208 3290
rect 14220 3238 14272 3290
rect 14284 3238 14336 3290
rect 1492 3136 1544 3188
rect 5632 3136 5684 3188
rect 6184 3179 6236 3188
rect 6184 3145 6193 3179
rect 6193 3145 6227 3179
rect 6227 3145 6236 3179
rect 6184 3136 6236 3145
rect 7104 3136 7156 3188
rect 10600 3179 10652 3188
rect 10600 3145 10609 3179
rect 10609 3145 10643 3179
rect 10643 3145 10652 3179
rect 10600 3136 10652 3145
rect 11336 3179 11388 3188
rect 11336 3145 11345 3179
rect 11345 3145 11379 3179
rect 11379 3145 11388 3179
rect 11336 3136 11388 3145
rect 13176 3136 13228 3188
rect 16304 3136 16356 3188
rect 4804 3068 4856 3120
rect 5172 3068 5224 3120
rect 3424 2975 3476 2984
rect 3424 2941 3433 2975
rect 3433 2941 3467 2975
rect 3467 2941 3476 2975
rect 3424 2932 3476 2941
rect 2412 2864 2464 2916
rect 3792 2907 3844 2916
rect 3792 2873 3801 2907
rect 3801 2873 3835 2907
rect 3835 2873 3844 2907
rect 3792 2864 3844 2873
rect 4252 2864 4304 2916
rect 5632 2975 5684 2984
rect 5632 2941 5641 2975
rect 5641 2941 5675 2975
rect 5675 2941 5684 2975
rect 5632 2932 5684 2941
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 7196 2975 7248 2984
rect 7196 2941 7205 2975
rect 7205 2941 7239 2975
rect 7239 2941 7248 2975
rect 8760 3068 8812 3120
rect 11152 3068 11204 3120
rect 12440 3068 12492 3120
rect 7196 2932 7248 2941
rect 8392 2975 8444 2984
rect 8392 2941 8401 2975
rect 8401 2941 8435 2975
rect 8435 2941 8444 2975
rect 8392 2932 8444 2941
rect 8576 2975 8628 2984
rect 8576 2941 8585 2975
rect 8585 2941 8619 2975
rect 8619 2941 8628 2975
rect 8576 2932 8628 2941
rect 6828 2864 6880 2916
rect 7104 2864 7156 2916
rect 8760 2975 8812 2984
rect 8760 2941 8769 2975
rect 8769 2941 8803 2975
rect 8803 2941 8812 2975
rect 8944 2975 8996 2984
rect 8760 2932 8812 2941
rect 8944 2941 8953 2975
rect 8953 2941 8987 2975
rect 8987 2941 8996 2975
rect 8944 2932 8996 2941
rect 9404 2975 9456 2984
rect 9404 2941 9413 2975
rect 9413 2941 9447 2975
rect 9447 2941 9456 2975
rect 9404 2932 9456 2941
rect 10048 2975 10100 2984
rect 10048 2941 10057 2975
rect 10057 2941 10091 2975
rect 10091 2941 10100 2975
rect 10048 2932 10100 2941
rect 10140 2975 10192 2984
rect 10140 2941 10149 2975
rect 10149 2941 10183 2975
rect 10183 2941 10192 2975
rect 10140 2932 10192 2941
rect 10324 2932 10376 2984
rect 11796 2932 11848 2984
rect 11888 2975 11940 2984
rect 11888 2941 11897 2975
rect 11897 2941 11931 2975
rect 11931 2941 11940 2975
rect 11888 2932 11940 2941
rect 12164 2932 12216 2984
rect 14096 3068 14148 3120
rect 14556 3000 14608 3052
rect 15568 3000 15620 3052
rect 13360 2932 13412 2984
rect 9588 2839 9640 2848
rect 9588 2805 9597 2839
rect 9597 2805 9631 2839
rect 9631 2805 9640 2839
rect 9588 2796 9640 2805
rect 10232 2796 10284 2848
rect 11980 2907 12032 2916
rect 11980 2873 11989 2907
rect 11989 2873 12023 2907
rect 12023 2873 12032 2907
rect 11980 2864 12032 2873
rect 12716 2907 12768 2916
rect 12716 2873 12725 2907
rect 12725 2873 12759 2907
rect 12759 2873 12768 2907
rect 12716 2864 12768 2873
rect 15752 2864 15804 2916
rect 6226 2694 6278 2746
rect 6290 2694 6342 2746
rect 6354 2694 6406 2746
rect 6418 2694 6470 2746
rect 11470 2694 11522 2746
rect 11534 2694 11586 2746
rect 11598 2694 11650 2746
rect 11662 2694 11714 2746
rect 3424 2592 3476 2644
rect 3792 2592 3844 2644
rect 5724 2592 5776 2644
rect 4988 2567 5040 2576
rect 4988 2533 4997 2567
rect 4997 2533 5031 2567
rect 5031 2533 5040 2567
rect 4988 2524 5040 2533
rect 7104 2592 7156 2644
rect 7380 2592 7432 2644
rect 7840 2592 7892 2644
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 6828 2524 6880 2576
rect 480 2456 532 2508
rect 1860 2499 1912 2508
rect 1860 2465 1869 2499
rect 1869 2465 1903 2499
rect 1903 2465 1912 2499
rect 1860 2456 1912 2465
rect 3424 2456 3476 2508
rect 4068 2499 4120 2508
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4068 2456 4120 2465
rect 4436 2499 4488 2508
rect 4436 2465 4445 2499
rect 4445 2465 4479 2499
rect 4479 2465 4488 2499
rect 4436 2456 4488 2465
rect 4712 2499 4764 2508
rect 4712 2465 4721 2499
rect 4721 2465 4755 2499
rect 4755 2465 4764 2499
rect 4712 2456 4764 2465
rect 4620 2388 4672 2440
rect 5080 2499 5132 2508
rect 5080 2465 5089 2499
rect 5089 2465 5123 2499
rect 5123 2465 5132 2499
rect 5080 2456 5132 2465
rect 4896 2320 4948 2372
rect 5632 2320 5684 2372
rect 6920 2363 6972 2372
rect 6920 2329 6929 2363
rect 6929 2329 6963 2363
rect 6963 2329 6972 2363
rect 6920 2320 6972 2329
rect 7012 2320 7064 2372
rect 8300 2456 8352 2508
rect 8576 2456 8628 2508
rect 8944 2524 8996 2576
rect 9588 2524 9640 2576
rect 10232 2524 10284 2576
rect 11796 2592 11848 2644
rect 11520 2456 11572 2508
rect 11980 2499 12032 2508
rect 11980 2465 12022 2499
rect 12022 2465 12032 2499
rect 11980 2456 12032 2465
rect 12716 2592 12768 2644
rect 15200 2635 15252 2644
rect 15200 2601 15209 2635
rect 15209 2601 15243 2635
rect 15243 2601 15252 2635
rect 15200 2592 15252 2601
rect 15752 2635 15804 2644
rect 15752 2601 15761 2635
rect 15761 2601 15795 2635
rect 15795 2601 15804 2635
rect 15752 2592 15804 2601
rect 16028 2635 16080 2644
rect 16028 2601 16037 2635
rect 16037 2601 16071 2635
rect 16071 2601 16080 2635
rect 16028 2592 16080 2601
rect 14556 2456 14608 2508
rect 14648 2456 14700 2508
rect 15200 2456 15252 2508
rect 16488 2499 16540 2508
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 16488 2465 16497 2499
rect 16497 2465 16531 2499
rect 16531 2465 16540 2499
rect 16488 2456 16540 2465
rect 16580 2388 16632 2440
rect 3976 2252 4028 2304
rect 7196 2252 7248 2304
rect 8024 2320 8076 2372
rect 7840 2252 7892 2304
rect 15844 2320 15896 2372
rect 3604 2150 3656 2202
rect 3668 2150 3720 2202
rect 3732 2150 3784 2202
rect 3796 2150 3848 2202
rect 8848 2150 8900 2202
rect 8912 2150 8964 2202
rect 8976 2150 9028 2202
rect 9040 2150 9092 2202
rect 14092 2150 14144 2202
rect 14156 2150 14208 2202
rect 14220 2150 14272 2202
rect 14284 2150 14336 2202
rect 3976 2048 4028 2100
rect 7748 2048 7800 2100
<< metal2 >>
rect 478 19371 534 20171
rect 2318 19371 2374 20171
rect 3698 19371 3754 20171
rect 5538 19371 5594 20171
rect 6918 19371 6974 20171
rect 8758 19371 8814 20171
rect 10138 19371 10194 20171
rect 11978 19371 12034 20171
rect 13818 19371 13874 20171
rect 15198 19371 15254 20171
rect 17038 19371 17094 20171
rect 492 17746 520 19371
rect 2332 17746 2360 19371
rect 3712 17746 3740 19371
rect 5080 17876 5132 17882
rect 5080 17818 5132 17824
rect 480 17740 532 17746
rect 480 17682 532 17688
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 3700 17740 3752 17746
rect 3700 17682 3752 17688
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4252 17604 4304 17610
rect 4252 17546 4304 17552
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 1400 17128 1452 17134
rect 1398 17096 1400 17105
rect 1452 17096 1454 17105
rect 1398 17031 1454 17040
rect 1596 16114 1624 17478
rect 3578 17436 3874 17456
rect 3634 17434 3658 17436
rect 3714 17434 3738 17436
rect 3794 17434 3818 17436
rect 3656 17382 3658 17434
rect 3720 17382 3732 17434
rect 3794 17382 3796 17434
rect 3634 17380 3658 17382
rect 3714 17380 3738 17382
rect 3794 17380 3818 17382
rect 3578 17360 3874 17380
rect 2688 17264 2740 17270
rect 2688 17206 2740 17212
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 15570 1808 15846
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1768 15564 1820 15570
rect 1768 15506 1820 15512
rect 2320 15564 2372 15570
rect 2320 15506 2372 15512
rect 1412 15065 1440 15506
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 1492 14952 1544 14958
rect 1492 14894 1544 14900
rect 1504 14414 1532 14894
rect 2332 14890 2360 15506
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 2320 14884 2372 14890
rect 2320 14826 2372 14832
rect 2424 14414 2452 14962
rect 2516 14958 2544 15642
rect 2504 14952 2556 14958
rect 2504 14894 2556 14900
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2608 14482 2636 14758
rect 2596 14476 2648 14482
rect 2596 14418 2648 14424
rect 1492 14408 1544 14414
rect 1492 14350 1544 14356
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2228 12708 2280 12714
rect 2228 12650 2280 12656
rect 2136 12368 2188 12374
rect 1398 12336 1454 12345
rect 2136 12310 2188 12316
rect 1398 12271 1400 12280
rect 1452 12271 1454 12280
rect 1400 12242 1452 12248
rect 1582 12200 1638 12209
rect 1582 12135 1584 12144
rect 1636 12135 1638 12144
rect 1584 12106 1636 12112
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1780 11694 1808 12038
rect 1768 11688 1820 11694
rect 1768 11630 1820 11636
rect 1584 11212 1636 11218
rect 1584 11154 1636 11160
rect 1398 10296 1454 10305
rect 1398 10231 1454 10240
rect 1412 10130 1440 10231
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1412 7585 1440 7890
rect 1398 7576 1454 7585
rect 1398 7511 1454 7520
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1412 6798 1440 7278
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1412 5545 1440 5714
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 1504 5234 1532 6598
rect 1596 5914 1624 11154
rect 2148 11082 2176 12310
rect 2240 11626 2268 12650
rect 2228 11620 2280 11626
rect 2228 11562 2280 11568
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 2148 10606 2176 11018
rect 2136 10600 2188 10606
rect 2136 10542 2188 10548
rect 2148 10130 2176 10542
rect 2240 10538 2268 11562
rect 2332 11082 2360 14350
rect 2424 13394 2452 14350
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 2424 11694 2452 13330
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2700 11218 2728 17206
rect 3988 17202 4016 17478
rect 4264 17270 4292 17546
rect 4344 17536 4396 17542
rect 4344 17478 4396 17484
rect 4252 17264 4304 17270
rect 4252 17206 4304 17212
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 3578 16348 3874 16368
rect 3634 16346 3658 16348
rect 3714 16346 3738 16348
rect 3794 16346 3818 16348
rect 3656 16294 3658 16346
rect 3720 16294 3732 16346
rect 3794 16294 3796 16346
rect 3634 16292 3658 16294
rect 3714 16292 3738 16294
rect 3794 16292 3818 16294
rect 3578 16272 3874 16292
rect 4080 16250 4108 17070
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3252 15638 3280 15846
rect 3240 15632 3292 15638
rect 3240 15574 3292 15580
rect 3578 15260 3874 15280
rect 3634 15258 3658 15260
rect 3714 15258 3738 15260
rect 3794 15258 3818 15260
rect 3656 15206 3658 15258
rect 3720 15206 3732 15258
rect 3794 15206 3796 15258
rect 3634 15204 3658 15206
rect 3714 15204 3738 15206
rect 3794 15204 3818 15206
rect 3578 15184 3874 15204
rect 3988 15162 4016 15982
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 4080 15094 4108 16186
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 4356 14618 4384 17478
rect 4448 17338 4476 17614
rect 4896 17604 4948 17610
rect 4896 17546 4948 17552
rect 4436 17332 4488 17338
rect 4436 17274 4488 17280
rect 4908 16794 4936 17546
rect 5092 17338 5120 17818
rect 5552 17746 5580 19371
rect 6200 17980 6496 18000
rect 6256 17978 6280 17980
rect 6336 17978 6360 17980
rect 6416 17978 6440 17980
rect 6278 17926 6280 17978
rect 6342 17926 6354 17978
rect 6416 17926 6418 17978
rect 6256 17924 6280 17926
rect 6336 17924 6360 17926
rect 6416 17924 6440 17926
rect 6200 17904 6496 17924
rect 6932 17814 6960 19371
rect 6920 17808 6972 17814
rect 6920 17750 6972 17756
rect 8772 17746 8800 19371
rect 10152 17746 10180 19371
rect 11444 17980 11740 18000
rect 11500 17978 11524 17980
rect 11580 17978 11604 17980
rect 11660 17978 11684 17980
rect 11522 17926 11524 17978
rect 11586 17926 11598 17978
rect 11660 17926 11662 17978
rect 11500 17924 11524 17926
rect 11580 17924 11604 17926
rect 11660 17924 11684 17926
rect 11444 17904 11740 17924
rect 11992 17746 12020 19371
rect 13832 17746 13860 19371
rect 15212 17746 15240 19371
rect 16118 18456 16174 18465
rect 16118 18391 16174 18400
rect 16132 17746 16160 18391
rect 17052 17814 17080 19371
rect 17040 17808 17092 17814
rect 17040 17750 17092 17756
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 8760 17740 8812 17746
rect 8760 17682 8812 17688
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 5724 17536 5776 17542
rect 5724 17478 5776 17484
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5092 16794 5120 17274
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5080 16652 5132 16658
rect 5184 16640 5212 17070
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5132 16612 5212 16640
rect 5080 16594 5132 16600
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4724 16182 4752 16390
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 5092 16046 5120 16594
rect 5644 16250 5672 16934
rect 5632 16244 5684 16250
rect 5632 16186 5684 16192
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 4436 15360 4488 15366
rect 4436 15302 4488 15308
rect 4448 15026 4476 15302
rect 4436 15020 4488 15026
rect 4436 14962 4488 14968
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4540 14414 4568 14962
rect 5540 14884 5592 14890
rect 5540 14826 5592 14832
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 3148 14272 3200 14278
rect 3148 14214 3200 14220
rect 3160 12850 3188 14214
rect 3578 14172 3874 14192
rect 3634 14170 3658 14172
rect 3714 14170 3738 14172
rect 3794 14170 3818 14172
rect 3656 14118 3658 14170
rect 3720 14118 3732 14170
rect 3794 14118 3796 14170
rect 3634 14116 3658 14118
rect 3714 14116 3738 14118
rect 3794 14116 3818 14118
rect 3578 14096 3874 14116
rect 4252 13728 4304 13734
rect 4252 13670 4304 13676
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4264 13462 4292 13670
rect 4252 13456 4304 13462
rect 3882 13424 3938 13433
rect 4252 13398 4304 13404
rect 3938 13368 4016 13376
rect 3882 13359 3884 13368
rect 3936 13348 4016 13368
rect 3884 13330 3936 13336
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 2780 12844 2832 12850
rect 2780 12786 2832 12792
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 2792 12306 2820 12786
rect 3252 12782 3280 13126
rect 3578 13084 3874 13104
rect 3634 13082 3658 13084
rect 3714 13082 3738 13084
rect 3794 13082 3818 13084
rect 3656 13030 3658 13082
rect 3720 13030 3732 13082
rect 3794 13030 3796 13082
rect 3634 13028 3658 13030
rect 3714 13028 3738 13030
rect 3794 13028 3818 13030
rect 3578 13008 3874 13028
rect 3988 12782 4016 13348
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4448 12850 4476 13126
rect 4816 12918 4844 13670
rect 5170 13424 5226 13433
rect 5170 13359 5172 13368
rect 5224 13359 5226 13368
rect 5172 13330 5224 13336
rect 4804 12912 4856 12918
rect 4804 12854 4856 12860
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 3578 11996 3874 12016
rect 3634 11994 3658 11996
rect 3714 11994 3738 11996
rect 3794 11994 3818 11996
rect 3656 11942 3658 11994
rect 3720 11942 3732 11994
rect 3794 11942 3796 11994
rect 3634 11940 3658 11942
rect 3714 11940 3738 11942
rect 3794 11940 3818 11942
rect 3578 11920 3874 11940
rect 5000 11694 5028 12582
rect 5368 12306 5396 14758
rect 5552 14550 5580 14826
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 3332 11280 3384 11286
rect 3332 11222 3384 11228
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 2320 11076 2372 11082
rect 2320 11018 2372 11024
rect 3160 10674 3188 11086
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2228 10532 2280 10538
rect 2228 10474 2280 10480
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2240 9518 2268 10474
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 2056 9042 2084 9318
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 2332 7954 2360 9998
rect 2792 9586 2820 10542
rect 3160 10130 3188 10610
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3252 10266 3280 10406
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 3160 9110 3188 10066
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2332 7018 2360 7890
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 7274 2452 7686
rect 2608 7290 2636 8774
rect 3160 8090 3188 8910
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2700 7410 2728 7686
rect 2976 7410 3004 7890
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2412 7268 2464 7274
rect 2608 7262 2728 7290
rect 2412 7210 2464 7216
rect 2332 6990 2636 7018
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2516 6458 2544 6870
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2608 6254 2636 6990
rect 2700 6712 2728 7262
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3252 6798 3280 7142
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 2780 6724 2832 6730
rect 2700 6684 2780 6712
rect 2780 6666 2832 6672
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1412 2825 1440 3538
rect 1504 3194 1532 5170
rect 2608 5098 2636 6190
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3160 5234 3188 5510
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 2596 5092 2648 5098
rect 2596 5034 2648 5040
rect 1584 4004 1636 4010
rect 1584 3946 1636 3952
rect 1596 3738 1624 3946
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 2608 3602 2636 5034
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2412 3392 2464 3398
rect 2412 3334 2464 3340
rect 1492 3188 1544 3194
rect 1492 3130 1544 3136
rect 2424 2922 2452 3334
rect 2412 2916 2464 2922
rect 2412 2858 2464 2864
rect 1398 2816 1454 2825
rect 1398 2751 1454 2760
rect 3344 2774 3372 11222
rect 4356 11218 4384 11494
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 3578 10908 3874 10928
rect 3634 10906 3658 10908
rect 3714 10906 3738 10908
rect 3794 10906 3818 10908
rect 3656 10854 3658 10906
rect 3720 10854 3732 10906
rect 3794 10854 3796 10906
rect 3634 10852 3658 10854
rect 3714 10852 3738 10854
rect 3794 10852 3818 10854
rect 3578 10832 3874 10852
rect 4356 10606 4384 11154
rect 4804 10736 4856 10742
rect 4804 10678 4856 10684
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4816 10470 4844 10678
rect 5092 10606 5120 11290
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5552 10470 5580 14486
rect 5644 14414 5672 15982
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 3578 9820 3874 9840
rect 3634 9818 3658 9820
rect 3714 9818 3738 9820
rect 3794 9818 3818 9820
rect 3656 9766 3658 9818
rect 3720 9766 3732 9818
rect 3794 9766 3796 9818
rect 3634 9764 3658 9766
rect 3714 9764 3738 9766
rect 3794 9764 3818 9766
rect 3578 9744 3874 9764
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3620 9178 3648 9454
rect 3896 9178 3924 9454
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 4356 9110 4384 9318
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 3578 8732 3874 8752
rect 3634 8730 3658 8732
rect 3714 8730 3738 8732
rect 3794 8730 3818 8732
rect 3656 8678 3658 8730
rect 3720 8678 3732 8730
rect 3794 8678 3796 8730
rect 3634 8676 3658 8678
rect 3714 8676 3738 8678
rect 3794 8676 3818 8678
rect 3578 8656 3874 8676
rect 4356 8430 4384 9046
rect 4724 9042 4752 9522
rect 4816 9450 4844 10406
rect 5644 9654 5672 13806
rect 5736 13530 5764 17478
rect 6564 17338 6592 17682
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 6000 17060 6052 17066
rect 6000 17002 6052 17008
rect 6012 16794 6040 17002
rect 6200 16892 6496 16912
rect 6256 16890 6280 16892
rect 6336 16890 6360 16892
rect 6416 16890 6440 16892
rect 6278 16838 6280 16890
rect 6342 16838 6354 16890
rect 6416 16838 6418 16890
rect 6256 16836 6280 16838
rect 6336 16836 6360 16838
rect 6416 16836 6440 16838
rect 6200 16816 6496 16836
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 7208 16658 7236 17070
rect 8404 16726 8432 17070
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 5920 15094 5948 16594
rect 5908 15088 5960 15094
rect 5908 15030 5960 15036
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 4804 9444 4856 9450
rect 4804 9386 4856 9392
rect 5552 9178 5580 9454
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5552 9042 5580 9114
rect 5644 9110 5672 9590
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4908 8634 4936 8910
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 3578 7644 3874 7664
rect 3634 7642 3658 7644
rect 3714 7642 3738 7644
rect 3794 7642 3818 7644
rect 3656 7590 3658 7642
rect 3720 7590 3732 7642
rect 3794 7590 3796 7642
rect 3634 7588 3658 7590
rect 3714 7588 3738 7590
rect 3794 7588 3818 7590
rect 3578 7568 3874 7588
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3436 7342 3464 7482
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 4068 7336 4120 7342
rect 4172 7324 4200 7890
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4448 7342 4476 7482
rect 4120 7296 4200 7324
rect 4068 7278 4120 7284
rect 3436 6254 3464 7278
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3528 7002 3556 7210
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 3578 6556 3874 6576
rect 3634 6554 3658 6556
rect 3714 6554 3738 6556
rect 3794 6554 3818 6556
rect 3656 6502 3658 6554
rect 3720 6502 3732 6554
rect 3794 6502 3796 6554
rect 3634 6500 3658 6502
rect 3714 6500 3738 6502
rect 3794 6500 3818 6502
rect 3578 6480 3874 6500
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 3436 5710 3464 6190
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3578 5468 3874 5488
rect 3634 5466 3658 5468
rect 3714 5466 3738 5468
rect 3794 5466 3818 5468
rect 3656 5414 3658 5466
rect 3720 5414 3732 5466
rect 3794 5414 3796 5466
rect 3634 5412 3658 5414
rect 3714 5412 3738 5414
rect 3794 5412 3818 5414
rect 3578 5392 3874 5412
rect 3578 4380 3874 4400
rect 3634 4378 3658 4380
rect 3714 4378 3738 4380
rect 3794 4378 3818 4380
rect 3656 4326 3658 4378
rect 3720 4326 3732 4378
rect 3794 4326 3796 4378
rect 3634 4324 3658 4326
rect 3714 4324 3738 4326
rect 3794 4324 3818 4326
rect 3578 4304 3874 4324
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3436 2990 3464 3538
rect 3578 3292 3874 3312
rect 3634 3290 3658 3292
rect 3714 3290 3738 3292
rect 3794 3290 3818 3292
rect 3656 3238 3658 3290
rect 3720 3238 3732 3290
rect 3794 3238 3796 3290
rect 3634 3236 3658 3238
rect 3714 3236 3738 3238
rect 3794 3236 3818 3238
rect 3578 3216 3874 3236
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3792 2916 3844 2922
rect 3792 2858 3844 2864
rect 3344 2746 3464 2774
rect 3436 2650 3464 2746
rect 3804 2650 3832 2858
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 4080 2514 4108 6190
rect 4172 5914 4200 7296
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 5724 7268 5776 7274
rect 5724 7210 5776 7216
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 4356 6798 4384 7142
rect 4724 6798 4752 7142
rect 5276 6934 5304 7142
rect 5736 7002 5764 7210
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5276 6118 5304 6734
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5276 5914 5304 6054
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4172 5234 4200 5510
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4264 5030 4292 5714
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4344 5296 4396 5302
rect 4344 5238 4396 5244
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4356 4690 4384 5238
rect 4632 5166 4660 5646
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4528 5024 4580 5030
rect 4632 5012 4660 5102
rect 4712 5024 4764 5030
rect 4632 4984 4712 5012
rect 4528 4966 4580 4972
rect 4712 4966 4764 4972
rect 4540 4690 4568 4966
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 4356 3738 4384 4626
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4264 2922 4292 3334
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4448 2514 4476 3878
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4632 3466 4660 3538
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 480 2508 532 2514
rect 480 2450 532 2456
rect 1860 2508 1912 2514
rect 1860 2450 1912 2456
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 492 800 520 2450
rect 1872 800 1900 2450
rect 3436 1306 3464 2450
rect 4632 2446 4660 3402
rect 4804 3120 4856 3126
rect 4724 3080 4804 3108
rect 4724 2514 4752 3080
rect 4804 3062 4856 3068
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4908 2378 4936 4082
rect 5092 4078 5120 4422
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 5276 3942 5304 5850
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5460 5098 5488 5510
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5552 4060 5580 4762
rect 5724 4684 5776 4690
rect 5644 4644 5724 4672
rect 5644 4214 5672 4644
rect 5724 4626 5776 4632
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5736 4214 5764 4490
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 5724 4208 5776 4214
rect 5724 4150 5776 4156
rect 5632 4072 5684 4078
rect 5552 4032 5632 4060
rect 5632 4014 5684 4020
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5184 3602 5212 3674
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 5000 2582 5028 3470
rect 5184 3126 5212 3538
rect 5644 3194 5672 4014
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 4988 2576 5040 2582
rect 4988 2518 5040 2524
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 4896 2372 4948 2378
rect 4896 2314 4948 2320
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3578 2204 3874 2224
rect 3634 2202 3658 2204
rect 3714 2202 3738 2204
rect 3794 2202 3818 2204
rect 3656 2150 3658 2202
rect 3720 2150 3732 2202
rect 3794 2150 3796 2202
rect 3634 2148 3658 2150
rect 3714 2148 3738 2150
rect 3794 2148 3818 2150
rect 3578 2128 3874 2148
rect 3988 2106 4016 2246
rect 3976 2100 4028 2106
rect 3976 2042 4028 2048
rect 3436 1278 3740 1306
rect 3712 800 3740 1278
rect 5092 800 5120 2450
rect 5644 2378 5672 2926
rect 5828 2774 5856 14962
rect 6000 14884 6052 14890
rect 5920 14844 6000 14872
rect 5920 14278 5948 14844
rect 6000 14826 6052 14832
rect 6104 14618 6132 16594
rect 8128 16250 8156 16594
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6200 15804 6496 15824
rect 6256 15802 6280 15804
rect 6336 15802 6360 15804
rect 6416 15802 6440 15804
rect 6278 15750 6280 15802
rect 6342 15750 6354 15802
rect 6416 15750 6418 15802
rect 6256 15748 6280 15750
rect 6336 15748 6360 15750
rect 6416 15748 6440 15750
rect 6200 15728 6496 15748
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 6200 14716 6496 14736
rect 6256 14714 6280 14716
rect 6336 14714 6360 14716
rect 6416 14714 6440 14716
rect 6278 14662 6280 14714
rect 6342 14662 6354 14714
rect 6416 14662 6418 14714
rect 6256 14660 6280 14662
rect 6336 14660 6360 14662
rect 6416 14660 6440 14662
rect 6200 14640 6496 14660
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 6182 14512 6238 14521
rect 6182 14447 6184 14456
rect 6236 14447 6238 14456
rect 6184 14418 6236 14424
rect 5998 14376 6054 14385
rect 6054 14320 6132 14328
rect 5998 14311 6000 14320
rect 6052 14300 6132 14320
rect 6000 14282 6052 14288
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5920 12850 5948 14214
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 6012 10742 6040 13262
rect 6104 12714 6132 14300
rect 6200 13628 6496 13648
rect 6256 13626 6280 13628
rect 6336 13626 6360 13628
rect 6416 13626 6440 13628
rect 6278 13574 6280 13626
rect 6342 13574 6354 13626
rect 6416 13574 6418 13626
rect 6256 13572 6280 13574
rect 6336 13572 6360 13574
rect 6416 13572 6440 13574
rect 6200 13552 6496 13572
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6472 12986 6500 13330
rect 6564 13326 6592 14962
rect 6644 14408 6696 14414
rect 6642 14376 6644 14385
rect 6696 14376 6698 14385
rect 6642 14311 6698 14320
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6840 12986 6868 16050
rect 8128 15910 8156 16186
rect 8588 16046 8616 17002
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8588 15706 8616 15982
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6932 14822 6960 14894
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6932 14521 6960 14758
rect 8588 14618 8616 15506
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 6918 14512 6974 14521
rect 6918 14447 6920 14456
rect 6972 14447 6974 14456
rect 7564 14476 7616 14482
rect 6920 14418 6972 14424
rect 7564 14418 7616 14424
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 6932 14387 6960 14418
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6092 12708 6144 12714
rect 6092 12650 6144 12656
rect 6104 12288 6132 12650
rect 6200 12540 6496 12560
rect 6256 12538 6280 12540
rect 6336 12538 6360 12540
rect 6416 12538 6440 12540
rect 6278 12486 6280 12538
rect 6342 12486 6354 12538
rect 6416 12486 6418 12538
rect 6256 12484 6280 12486
rect 6336 12484 6360 12486
rect 6416 12484 6440 12486
rect 6200 12464 6496 12484
rect 6104 12260 6224 12288
rect 6196 12102 6224 12260
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 6104 10588 6132 12038
rect 6564 11694 6592 12922
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6656 11830 6684 12786
rect 6932 12782 6960 14282
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6748 12306 6776 12718
rect 6932 12646 6960 12718
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6644 11824 6696 11830
rect 6644 11766 6696 11772
rect 6748 11694 6776 12242
rect 6932 12238 6960 12582
rect 7116 12306 7144 12786
rect 7208 12442 7236 12922
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6200 11452 6496 11472
rect 6256 11450 6280 11452
rect 6336 11450 6360 11452
rect 6416 11450 6440 11452
rect 6278 11398 6280 11450
rect 6342 11398 6354 11450
rect 6416 11398 6418 11450
rect 6256 11396 6280 11398
rect 6336 11396 6360 11398
rect 6416 11396 6440 11398
rect 6200 11376 6496 11396
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6472 10810 6500 10950
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6184 10600 6236 10606
rect 6104 10560 6184 10588
rect 6012 10266 6040 10542
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6104 9178 6132 10560
rect 6184 10542 6236 10548
rect 6200 10364 6496 10384
rect 6256 10362 6280 10364
rect 6336 10362 6360 10364
rect 6416 10362 6440 10364
rect 6278 10310 6280 10362
rect 6342 10310 6354 10362
rect 6416 10310 6418 10362
rect 6256 10308 6280 10310
rect 6336 10308 6360 10310
rect 6416 10308 6440 10310
rect 6200 10288 6496 10308
rect 6564 10130 6592 10610
rect 6656 10470 6684 10746
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6656 10198 6684 10406
rect 6748 10266 6776 11630
rect 6932 10810 6960 12174
rect 7208 11694 7236 12174
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7208 10606 7236 11630
rect 7300 10810 7328 13806
rect 7576 12986 7604 14418
rect 8036 13870 8064 14418
rect 8208 14000 8260 14006
rect 8312 13954 8340 14418
rect 8260 13948 8340 13954
rect 8208 13942 8340 13948
rect 8220 13926 8340 13942
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 8312 13734 8340 13926
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8680 13530 8708 17478
rect 8822 17436 9118 17456
rect 8878 17434 8902 17436
rect 8958 17434 8982 17436
rect 9038 17434 9062 17436
rect 8900 17382 8902 17434
rect 8964 17382 8976 17434
rect 9038 17382 9040 17434
rect 8878 17380 8902 17382
rect 8958 17380 8982 17382
rect 9038 17380 9062 17382
rect 8822 17360 9118 17380
rect 10796 17202 11100 17218
rect 10784 17196 11100 17202
rect 10836 17190 11100 17196
rect 10784 17138 10836 17144
rect 10968 17128 11020 17134
rect 10888 17076 10968 17082
rect 10888 17070 11020 17076
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10888 17054 11008 17070
rect 11072 17066 11100 17190
rect 11060 17060 11112 17066
rect 8822 16348 9118 16368
rect 8878 16346 8902 16348
rect 8958 16346 8982 16348
rect 9038 16346 9062 16348
rect 8900 16294 8902 16346
rect 8964 16294 8976 16346
rect 9038 16294 9040 16346
rect 8878 16292 8902 16294
rect 8958 16292 8982 16294
rect 9038 16292 9062 16294
rect 8822 16272 9118 16292
rect 9496 16176 9548 16182
rect 9496 16118 9548 16124
rect 9508 16046 9536 16118
rect 9876 16046 9904 17002
rect 10796 16794 10824 17002
rect 10888 16998 10916 17054
rect 11060 17002 11112 17008
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 11444 16892 11740 16912
rect 11500 16890 11524 16892
rect 11580 16890 11604 16892
rect 11660 16890 11684 16892
rect 11522 16838 11524 16890
rect 11586 16838 11598 16890
rect 11660 16838 11662 16890
rect 11500 16836 11524 16838
rect 11580 16836 11604 16838
rect 11660 16836 11684 16838
rect 11444 16816 11740 16836
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10704 16182 10732 16390
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 9496 16040 9548 16046
rect 9496 15982 9548 15988
rect 9864 16040 9916 16046
rect 9864 15982 9916 15988
rect 8822 15260 9118 15280
rect 8878 15258 8902 15260
rect 8958 15258 8982 15260
rect 9038 15258 9062 15260
rect 8900 15206 8902 15258
rect 8964 15206 8976 15258
rect 9038 15206 9040 15258
rect 8878 15204 8902 15206
rect 8958 15204 8982 15206
rect 9038 15204 9062 15206
rect 8822 15184 9118 15204
rect 9508 15162 9536 15982
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10520 15638 10548 15846
rect 11444 15804 11740 15824
rect 11500 15802 11524 15804
rect 11580 15802 11604 15804
rect 11660 15802 11684 15804
rect 11522 15750 11524 15802
rect 11586 15750 11598 15802
rect 11660 15750 11662 15802
rect 11500 15748 11524 15750
rect 11580 15748 11604 15750
rect 11660 15748 11684 15750
rect 11444 15728 11740 15748
rect 10508 15632 10560 15638
rect 10508 15574 10560 15580
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 10060 14482 10088 15030
rect 11336 14884 11388 14890
rect 11336 14826 11388 14832
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10428 14482 10456 14758
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10416 14476 10468 14482
rect 10416 14418 10468 14424
rect 8822 14172 9118 14192
rect 8878 14170 8902 14172
rect 8958 14170 8982 14172
rect 9038 14170 9062 14172
rect 8900 14118 8902 14170
rect 8964 14118 8976 14170
rect 9038 14118 9040 14170
rect 8878 14116 8902 14118
rect 8958 14116 8982 14118
rect 9038 14116 9062 14118
rect 8822 14096 9118 14116
rect 9232 14074 9260 14418
rect 11348 14414 11376 14826
rect 11444 14716 11740 14736
rect 11500 14714 11524 14716
rect 11580 14714 11604 14716
rect 11660 14714 11684 14716
rect 11522 14662 11524 14714
rect 11586 14662 11598 14714
rect 11660 14662 11662 14714
rect 11500 14660 11524 14662
rect 11580 14660 11604 14662
rect 11660 14660 11684 14662
rect 11444 14640 11740 14660
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 10612 13870 10640 14214
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11444 13628 11740 13648
rect 11500 13626 11524 13628
rect 11580 13626 11604 13628
rect 11660 13626 11684 13628
rect 11522 13574 11524 13626
rect 11586 13574 11598 13626
rect 11660 13574 11662 13626
rect 11500 13572 11524 13574
rect 11580 13572 11604 13574
rect 11660 13572 11684 13574
rect 11444 13552 11740 13572
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 10508 13456 10560 13462
rect 10508 13398 10560 13404
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 8588 12986 8616 13330
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 7392 11064 7420 12650
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 7852 12306 7880 12582
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7668 11626 7696 12038
rect 7944 11898 7972 12038
rect 7932 11892 7984 11898
rect 7852 11852 7932 11880
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7852 11354 7880 11852
rect 7932 11834 7984 11840
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7472 11076 7524 11082
rect 7392 11036 7472 11064
rect 7472 11018 7524 11024
rect 7760 10810 7788 11154
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7012 10600 7064 10606
rect 7196 10600 7248 10606
rect 7012 10542 7064 10548
rect 7194 10568 7196 10577
rect 7248 10568 7250 10577
rect 7024 10266 7052 10542
rect 7194 10503 7250 10512
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6200 9276 6496 9296
rect 6256 9274 6280 9276
rect 6336 9274 6360 9276
rect 6416 9274 6440 9276
rect 6278 9222 6280 9274
rect 6342 9222 6354 9274
rect 6416 9222 6418 9274
rect 6256 9220 6280 9222
rect 6336 9220 6360 9222
rect 6416 9220 6440 9222
rect 6200 9200 6496 9220
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6564 8974 6592 10066
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 6828 9444 6880 9450
rect 6828 9386 6880 9392
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6200 8188 6496 8208
rect 6256 8186 6280 8188
rect 6336 8186 6360 8188
rect 6416 8186 6440 8188
rect 6278 8134 6280 8186
rect 6342 8134 6354 8186
rect 6416 8134 6418 8186
rect 6256 8132 6280 8134
rect 6336 8132 6360 8134
rect 6416 8132 6440 8134
rect 6200 8112 6496 8132
rect 6748 7954 6776 8978
rect 6840 8634 6868 9386
rect 7024 9178 7052 9386
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 7116 8974 7144 9522
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6104 7342 6132 7890
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6104 5166 6132 7278
rect 6840 7274 6868 7686
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6828 7268 6880 7274
rect 6828 7210 6880 7216
rect 6200 7100 6496 7120
rect 6256 7098 6280 7100
rect 6336 7098 6360 7100
rect 6416 7098 6440 7100
rect 6278 7046 6280 7098
rect 6342 7046 6354 7098
rect 6416 7046 6418 7098
rect 6256 7044 6280 7046
rect 6336 7044 6360 7046
rect 6416 7044 6440 7046
rect 6200 7024 6496 7044
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 6656 6118 6684 6870
rect 6748 6730 6776 7210
rect 7116 7206 7144 8910
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6200 6012 6496 6032
rect 6256 6010 6280 6012
rect 6336 6010 6360 6012
rect 6416 6010 6440 6012
rect 6278 5958 6280 6010
rect 6342 5958 6354 6010
rect 6416 5958 6418 6010
rect 6256 5956 6280 5958
rect 6336 5956 6360 5958
rect 6416 5956 6440 5958
rect 6200 5936 6496 5956
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6380 5370 6408 5782
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6932 5234 6960 6802
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 7024 5166 7052 6190
rect 7208 6186 7236 6666
rect 7484 6662 7512 7142
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7116 5370 7144 5646
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 7208 5166 7236 6122
rect 7484 5914 7512 6598
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6012 4486 6040 4626
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 6104 3670 6132 5102
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6200 4924 6496 4944
rect 6256 4922 6280 4924
rect 6336 4922 6360 4924
rect 6416 4922 6440 4924
rect 6278 4870 6280 4922
rect 6342 4870 6354 4922
rect 6416 4870 6418 4922
rect 6256 4868 6280 4870
rect 6336 4868 6360 4870
rect 6416 4868 6440 4870
rect 6200 4848 6496 4868
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6196 4282 6224 4626
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6736 4072 6788 4078
rect 6932 4026 6960 4966
rect 7024 4146 7052 5102
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 6736 4014 6788 4020
rect 6656 3942 6684 4014
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6200 3836 6496 3856
rect 6256 3834 6280 3836
rect 6336 3834 6360 3836
rect 6416 3834 6440 3836
rect 6278 3782 6280 3834
rect 6342 3782 6354 3834
rect 6416 3782 6418 3834
rect 6256 3780 6280 3782
rect 6336 3780 6360 3782
rect 6416 3780 6440 3782
rect 6200 3760 6496 3780
rect 6092 3664 6144 3670
rect 6092 3606 6144 3612
rect 6656 3534 6684 3878
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 6196 3194 6224 3334
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6748 3074 6776 4014
rect 6840 4010 6960 4026
rect 6828 4004 6960 4010
rect 6880 3998 6960 4004
rect 6828 3946 6880 3952
rect 6932 3602 6960 3998
rect 7024 3738 7052 4082
rect 7116 3942 7144 5034
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7116 3602 7144 3878
rect 7208 3602 7236 5102
rect 7300 5030 7328 5102
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7392 4078 7420 5714
rect 7576 5710 7604 6054
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7116 3194 7144 3538
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 6748 3046 7052 3074
rect 7024 2961 7052 3046
rect 7208 2990 7236 3538
rect 7288 3460 7340 3466
rect 7288 3402 7340 3408
rect 7300 3058 7328 3402
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7196 2984 7248 2990
rect 7010 2952 7066 2961
rect 6828 2916 6880 2922
rect 7196 2926 7248 2932
rect 7010 2887 7066 2896
rect 7104 2916 7156 2922
rect 6828 2858 6880 2864
rect 5736 2746 5856 2774
rect 6200 2748 6496 2768
rect 6256 2746 6280 2748
rect 6336 2746 6360 2748
rect 6416 2746 6440 2748
rect 5736 2650 5764 2746
rect 6278 2694 6280 2746
rect 6342 2694 6354 2746
rect 6416 2694 6418 2746
rect 6256 2692 6280 2694
rect 6336 2692 6360 2694
rect 6416 2692 6440 2694
rect 6200 2672 6496 2692
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 6840 2582 6868 2858
rect 6828 2576 6880 2582
rect 6828 2518 6880 2524
rect 7024 2378 7052 2887
rect 7104 2858 7156 2864
rect 7116 2650 7144 2858
rect 7392 2650 7420 4014
rect 7104 2644 7156 2650
rect 7380 2644 7432 2650
rect 7104 2586 7156 2592
rect 7208 2604 7380 2632
rect 5632 2372 5684 2378
rect 5632 2314 5684 2320
rect 6920 2372 6972 2378
rect 6920 2314 6972 2320
rect 7012 2372 7064 2378
rect 7012 2314 7064 2320
rect 6932 800 6960 2314
rect 7208 2310 7236 2604
rect 7380 2586 7432 2592
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 7760 2106 7788 10406
rect 7852 9654 7880 11290
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 7944 10674 7972 11086
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7840 9648 7892 9654
rect 7840 9590 7892 9596
rect 7852 8498 7880 9590
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7932 7472 7984 7478
rect 7932 7414 7984 7420
rect 7944 6934 7972 7414
rect 7932 6928 7984 6934
rect 7932 6870 7984 6876
rect 7840 6248 7892 6254
rect 7944 6236 7972 6870
rect 7892 6208 7972 6236
rect 7840 6190 7892 6196
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7852 2310 7880 2586
rect 8036 2378 8064 12582
rect 8220 12102 8248 12718
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8312 12238 8340 12650
rect 8496 12374 8524 12854
rect 8680 12850 8708 13262
rect 8822 13084 9118 13104
rect 8878 13082 8902 13084
rect 8958 13082 8982 13084
rect 9038 13082 9062 13084
rect 8900 13030 8902 13082
rect 8964 13030 8976 13082
rect 9038 13030 9040 13082
rect 8878 13028 8902 13030
rect 8958 13028 8982 13030
rect 9038 13028 9062 13030
rect 8822 13008 9118 13028
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8300 12232 8352 12238
rect 8392 12232 8444 12238
rect 8300 12174 8352 12180
rect 8390 12200 8392 12209
rect 8444 12200 8446 12209
rect 8390 12135 8446 12144
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8496 11778 8524 12310
rect 9692 12238 9720 13262
rect 9876 12442 9904 13330
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 10152 12850 10180 13126
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9416 12073 9444 12106
rect 9402 12064 9458 12073
rect 8822 11996 9118 12016
rect 9402 11999 9458 12008
rect 8878 11994 8902 11996
rect 8958 11994 8982 11996
rect 9038 11994 9062 11996
rect 8900 11942 8902 11994
rect 8964 11942 8976 11994
rect 9038 11942 9040 11994
rect 8878 11940 8902 11942
rect 8958 11940 8982 11942
rect 9038 11940 9062 11942
rect 8822 11920 9118 11940
rect 8852 11824 8904 11830
rect 8496 11762 8616 11778
rect 8852 11766 8904 11772
rect 8944 11824 8996 11830
rect 8944 11766 8996 11772
rect 8496 11756 8628 11762
rect 8496 11750 8576 11756
rect 8576 11698 8628 11704
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8220 10606 8248 10950
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8220 7002 8248 7142
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8220 6390 8248 6938
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 8220 6254 8248 6326
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8312 2650 8340 11154
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8404 10674 8432 11018
rect 8496 11014 8524 11630
rect 8864 11529 8892 11766
rect 8850 11520 8906 11529
rect 8850 11455 8906 11464
rect 8956 11218 8984 11766
rect 9220 11552 9272 11558
rect 9272 11512 9352 11540
rect 9220 11494 9272 11500
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9036 11280 9088 11286
rect 9232 11234 9260 11290
rect 9088 11228 9260 11234
rect 9036 11222 9260 11228
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8944 11212 8996 11218
rect 9048 11206 9260 11222
rect 8944 11154 8996 11160
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8496 10538 8524 10950
rect 8680 10742 8708 11154
rect 8822 10908 9118 10928
rect 8878 10906 8902 10908
rect 8958 10906 8982 10908
rect 9038 10906 9062 10908
rect 8900 10854 8902 10906
rect 8964 10854 8976 10906
rect 9038 10854 9040 10906
rect 8878 10852 8902 10854
rect 8958 10852 8982 10854
rect 9038 10852 9062 10854
rect 8822 10832 9118 10852
rect 9232 10810 9260 11206
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 8668 10736 8720 10742
rect 9232 10690 9260 10746
rect 8668 10678 8720 10684
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 9048 10662 9260 10690
rect 8576 10600 8628 10606
rect 8864 10577 8892 10610
rect 9048 10606 9076 10662
rect 9036 10600 9088 10606
rect 8576 10542 8628 10548
rect 8850 10568 8906 10577
rect 8484 10532 8536 10538
rect 8484 10474 8536 10480
rect 8588 10441 8616 10542
rect 9036 10542 9088 10548
rect 9220 10600 9272 10606
rect 9324 10588 9352 11512
rect 9508 11268 9536 12106
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9680 11620 9732 11626
rect 9784 11608 9812 11834
rect 9876 11830 9904 12378
rect 10232 12368 10284 12374
rect 10232 12310 10284 12316
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 9732 11580 9812 11608
rect 9680 11562 9732 11568
rect 9588 11280 9640 11286
rect 9508 11240 9588 11268
rect 9588 11222 9640 11228
rect 9600 10742 9628 11222
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9956 11212 10008 11218
rect 10060 11200 10088 12242
rect 10244 12170 10272 12310
rect 10336 12306 10364 12582
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 10232 12164 10284 12170
rect 10232 12106 10284 12112
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10008 11172 10088 11200
rect 9956 11154 10008 11160
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 9272 10560 9352 10588
rect 9220 10542 9272 10548
rect 8850 10503 8906 10512
rect 8574 10432 8630 10441
rect 8574 10367 8630 10376
rect 8822 9820 9118 9840
rect 8878 9818 8902 9820
rect 8958 9818 8982 9820
rect 9038 9818 9062 9820
rect 8900 9766 8902 9818
rect 8964 9766 8976 9818
rect 9038 9766 9040 9818
rect 8878 9764 8902 9766
rect 8958 9764 8982 9766
rect 9038 9764 9062 9766
rect 8822 9744 9118 9764
rect 9232 9178 9260 10542
rect 9496 10532 9548 10538
rect 9496 10474 9548 10480
rect 9508 10441 9536 10474
rect 9494 10432 9550 10441
rect 9494 10367 9550 10376
rect 9600 9450 9628 10678
rect 9692 10606 9720 11154
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9784 10588 9812 11018
rect 10152 10810 10180 11834
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10232 10736 10284 10742
rect 10230 10704 10232 10713
rect 10284 10704 10286 10713
rect 10428 10674 10456 11154
rect 10230 10639 10286 10648
rect 10416 10668 10468 10674
rect 9864 10600 9916 10606
rect 9784 10560 9864 10588
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9600 9178 9628 9386
rect 9784 9382 9812 10560
rect 9864 10542 9916 10548
rect 10244 10266 10272 10639
rect 10416 10610 10468 10616
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8496 8634 8524 8978
rect 9784 8906 9812 9318
rect 10060 9042 10088 9454
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8588 8498 8616 8774
rect 8822 8732 9118 8752
rect 8878 8730 8902 8732
rect 8958 8730 8982 8732
rect 9038 8730 9062 8732
rect 8900 8678 8902 8730
rect 8964 8678 8976 8730
rect 9038 8678 9040 8730
rect 8878 8676 8902 8678
rect 8958 8676 8982 8678
rect 9038 8676 9062 8678
rect 8822 8656 9118 8676
rect 9692 8566 9720 8774
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8680 7954 8708 8366
rect 10244 8362 10272 8842
rect 10336 8634 10364 8978
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10428 8498 10456 9318
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 8822 7644 9118 7664
rect 8878 7642 8902 7644
rect 8958 7642 8982 7644
rect 9038 7642 9062 7644
rect 8900 7590 8902 7642
rect 8964 7590 8976 7642
rect 9038 7590 9040 7642
rect 8878 7588 8902 7590
rect 8958 7588 8982 7590
rect 9038 7588 9062 7590
rect 8822 7568 9118 7588
rect 9232 7274 9260 7686
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 8822 6556 9118 6576
rect 8878 6554 8902 6556
rect 8958 6554 8982 6556
rect 9038 6554 9062 6556
rect 8900 6502 8902 6554
rect 8964 6502 8976 6554
rect 9038 6502 9040 6554
rect 8878 6500 8902 6502
rect 8958 6500 8982 6502
rect 9038 6500 9062 6502
rect 8822 6480 9118 6500
rect 9784 6254 9812 7346
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9876 6730 9904 7210
rect 9864 6724 9916 6730
rect 9864 6666 9916 6672
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8404 5710 8432 6122
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8496 5234 8524 6054
rect 8864 5778 8892 6054
rect 10244 5914 10272 7278
rect 10324 7268 10376 7274
rect 10324 7210 10376 7216
rect 10336 6866 10364 7210
rect 10520 7154 10548 13398
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10612 12442 10640 13330
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10796 12782 10824 13194
rect 11808 12986 11836 13806
rect 11900 13530 11928 14418
rect 12084 13870 12112 16934
rect 12176 15026 12204 17478
rect 12452 17202 12480 17614
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 15200 17536 15252 17542
rect 15200 17478 15252 17484
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 14066 17436 14362 17456
rect 14122 17434 14146 17436
rect 14202 17434 14226 17436
rect 14282 17434 14306 17436
rect 14144 17382 14146 17434
rect 14208 17382 14220 17434
rect 14282 17382 14284 17434
rect 14122 17380 14146 17382
rect 14202 17380 14226 17382
rect 14282 17380 14306 17382
rect 14066 17360 14362 17380
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12544 16658 12572 17002
rect 12636 16726 12664 17206
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 12900 17060 12952 17066
rect 12900 17002 12952 17008
rect 12624 16720 12676 16726
rect 12624 16662 12676 16668
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12452 15026 12480 15438
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 12072 13864 12124 13870
rect 11992 13812 12072 13818
rect 11992 13806 12124 13812
rect 11992 13790 12112 13806
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11336 12844 11388 12850
rect 11256 12804 11336 12832
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10888 12374 10916 12718
rect 11256 12646 11284 12804
rect 11336 12786 11388 12792
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 11152 12300 11204 12306
rect 11256 12288 11284 12582
rect 11348 12442 11376 12650
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11444 12540 11740 12560
rect 11500 12538 11524 12540
rect 11580 12538 11604 12540
rect 11660 12538 11684 12540
rect 11522 12486 11524 12538
rect 11586 12486 11598 12538
rect 11660 12486 11662 12538
rect 11500 12484 11524 12486
rect 11580 12484 11604 12486
rect 11660 12484 11684 12486
rect 11444 12464 11740 12484
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11808 12306 11836 12582
rect 11992 12442 12020 13790
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 12084 13530 12112 13670
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 12084 12306 12112 12378
rect 11204 12260 11284 12288
rect 11796 12300 11848 12306
rect 11152 12242 11204 12248
rect 11796 12242 11848 12248
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10704 10538 10732 11630
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10796 10198 10824 12242
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10888 11354 10916 12174
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 11164 11762 11192 12106
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10888 10674 10916 11290
rect 11164 11218 11192 11698
rect 11444 11452 11740 11472
rect 11500 11450 11524 11452
rect 11580 11450 11604 11452
rect 11660 11450 11684 11452
rect 11522 11398 11524 11450
rect 11586 11398 11598 11450
rect 11660 11398 11662 11450
rect 11500 11396 11524 11398
rect 11580 11396 11604 11398
rect 11660 11396 11684 11398
rect 11444 11376 11740 11396
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11164 10810 11192 11154
rect 11440 11082 11468 11154
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 10876 10668 10928 10674
rect 10928 10628 11008 10656
rect 10876 10610 10928 10616
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10980 9586 11008 10628
rect 11164 10606 11192 10746
rect 11440 10606 11468 11018
rect 11532 10742 11560 11086
rect 11808 11082 11836 12242
rect 11992 12170 12020 12242
rect 11980 12164 12032 12170
rect 11980 12106 12032 12112
rect 11992 11762 12020 12106
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 12084 11694 12112 12242
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11624 10810 11652 10950
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11520 10736 11572 10742
rect 11520 10678 11572 10684
rect 11704 10736 11756 10742
rect 11756 10696 11836 10724
rect 11704 10678 11756 10684
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10876 9512 10928 9518
rect 10874 9480 10876 9489
rect 10928 9480 10930 9489
rect 11072 9450 11100 9930
rect 10874 9415 10930 9424
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 10782 9072 10838 9081
rect 10782 9007 10784 9016
rect 10836 9007 10838 9016
rect 10784 8978 10836 8984
rect 11164 8294 11192 10406
rect 11348 10198 11376 10406
rect 11444 10364 11740 10384
rect 11500 10362 11524 10364
rect 11580 10362 11604 10364
rect 11660 10362 11684 10364
rect 11522 10310 11524 10362
rect 11586 10310 11598 10362
rect 11660 10310 11662 10362
rect 11500 10308 11524 10310
rect 11580 10308 11604 10310
rect 11660 10308 11684 10310
rect 11444 10288 11740 10308
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11256 9110 11284 9590
rect 11808 9518 11836 10696
rect 11796 9512 11848 9518
rect 11888 9512 11940 9518
rect 11796 9454 11848 9460
rect 11886 9480 11888 9489
rect 11940 9480 11942 9489
rect 11886 9415 11942 9424
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11244 9104 11296 9110
rect 11244 9046 11296 9052
rect 11348 9042 11376 9318
rect 11444 9276 11740 9296
rect 11500 9274 11524 9276
rect 11580 9274 11604 9276
rect 11660 9274 11684 9276
rect 11522 9222 11524 9274
rect 11586 9222 11598 9274
rect 11660 9222 11662 9274
rect 11500 9220 11524 9222
rect 11580 9220 11604 9222
rect 11660 9220 11684 9222
rect 11444 9200 11740 9220
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11808 9081 11836 9114
rect 11794 9072 11850 9081
rect 11336 9036 11388 9042
rect 11794 9007 11850 9016
rect 11336 8978 11388 8984
rect 11348 8498 11376 8978
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11164 8266 11284 8294
rect 11256 8022 11284 8266
rect 11348 8090 11376 8434
rect 11444 8188 11740 8208
rect 11500 8186 11524 8188
rect 11580 8186 11604 8188
rect 11660 8186 11684 8188
rect 11522 8134 11524 8186
rect 11586 8134 11598 8186
rect 11660 8134 11662 8186
rect 11500 8132 11524 8134
rect 11580 8132 11604 8134
rect 11660 8132 11684 8134
rect 11444 8112 11740 8132
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 11256 7342 11284 7958
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11900 7546 11928 7890
rect 11992 7546 12020 11018
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 12084 9110 12112 9386
rect 12072 9104 12124 9110
rect 12072 9046 12124 9052
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 10784 7336 10836 7342
rect 10968 7336 11020 7342
rect 10784 7278 10836 7284
rect 10966 7304 10968 7313
rect 11244 7336 11296 7342
rect 11020 7304 11022 7313
rect 10520 7126 10640 7154
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 9220 5636 9272 5642
rect 9220 5578 9272 5584
rect 8822 5468 9118 5488
rect 8878 5466 8902 5468
rect 8958 5466 8982 5468
rect 9038 5466 9062 5468
rect 8900 5414 8902 5466
rect 8964 5414 8976 5466
rect 9038 5414 9040 5466
rect 8878 5412 8902 5414
rect 8958 5412 8982 5414
rect 9038 5412 9062 5414
rect 8822 5392 9118 5412
rect 9232 5234 9260 5578
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9232 4690 9260 5170
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 9416 4486 9444 4626
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 8822 4380 9118 4400
rect 8878 4378 8902 4380
rect 8958 4378 8982 4380
rect 9038 4378 9062 4380
rect 8900 4326 8902 4378
rect 8964 4326 8976 4378
rect 9038 4326 9040 4378
rect 8878 4324 8902 4326
rect 8958 4324 8982 4326
rect 9038 4324 9062 4326
rect 8822 4304 9118 4324
rect 9692 4282 9720 5102
rect 9876 4826 9904 5102
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9968 4486 9996 5646
rect 10152 5370 10180 5714
rect 10244 5710 10272 5850
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10244 4690 10272 5102
rect 10336 4758 10364 6190
rect 10520 5846 10548 6190
rect 10508 5840 10560 5846
rect 10508 5782 10560 5788
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 10520 4690 10548 5102
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 8668 4004 8720 4010
rect 8668 3946 8720 3952
rect 8680 3738 8708 3946
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 9404 3460 9456 3466
rect 9404 3402 9456 3408
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8404 2990 8432 3334
rect 8822 3292 9118 3312
rect 8878 3290 8902 3292
rect 8958 3290 8982 3292
rect 9038 3290 9062 3292
rect 8900 3238 8902 3290
rect 8964 3238 8976 3290
rect 9038 3238 9040 3290
rect 8878 3236 8902 3238
rect 8958 3236 8982 3238
rect 9038 3236 9062 3238
rect 8822 3216 9118 3236
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8772 2990 8800 3062
rect 9416 2990 9444 3402
rect 10060 2990 10088 3878
rect 10152 3602 10180 4218
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10152 2990 10180 3538
rect 10612 3194 10640 7126
rect 10796 6458 10824 7278
rect 11244 7278 11296 7284
rect 10966 7239 11022 7248
rect 11444 7100 11740 7120
rect 11500 7098 11524 7100
rect 11580 7098 11604 7100
rect 11660 7098 11684 7100
rect 11522 7046 11524 7098
rect 11586 7046 11598 7098
rect 11660 7046 11662 7098
rect 11500 7044 11524 7046
rect 11580 7044 11604 7046
rect 11660 7044 11684 7046
rect 11444 7024 11740 7044
rect 11900 6866 11928 7482
rect 11980 7268 12032 7274
rect 11980 7210 12032 7216
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11532 6730 11928 6746
rect 11532 6724 11940 6730
rect 11532 6718 11888 6724
rect 11532 6662 11560 6718
rect 11888 6666 11940 6672
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 11992 6322 12020 7210
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 12176 6254 12204 12854
rect 12360 12442 12388 14758
rect 12452 13326 12480 14962
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12820 12306 12848 12786
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12714 12064 12770 12073
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12268 11694 12296 11834
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12268 10674 12296 11630
rect 12360 11150 12388 12038
rect 12714 11999 12770 12008
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12452 11694 12480 11766
rect 12728 11694 12756 11999
rect 12820 11762 12848 12242
rect 12912 11898 12940 17002
rect 13188 15502 13216 17138
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13372 16114 13400 16594
rect 13820 16584 13872 16590
rect 15028 16574 15056 17478
rect 15212 17338 15240 17478
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15948 17134 15976 17478
rect 15936 17128 15988 17134
rect 15936 17070 15988 17076
rect 13820 16526 13872 16532
rect 14752 16546 15056 16574
rect 13832 16250 13860 16526
rect 14066 16348 14362 16368
rect 14122 16346 14146 16348
rect 14202 16346 14226 16348
rect 14282 16346 14306 16348
rect 14144 16294 14146 16346
rect 14208 16294 14220 16346
rect 14282 16294 14284 16346
rect 14122 16292 14146 16294
rect 14202 16292 14226 16294
rect 14282 16292 14306 16294
rect 14066 16272 14362 16292
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13464 15570 13492 15982
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13740 15706 13768 15846
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13924 15570 13952 15982
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13176 12368 13228 12374
rect 13176 12310 13228 12316
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 13084 11824 13136 11830
rect 13084 11766 13136 11772
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12360 10996 12388 11086
rect 12360 10968 12480 10996
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12360 10130 12388 10746
rect 12452 10606 12480 10968
rect 12622 10704 12678 10713
rect 12622 10639 12678 10648
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12636 10588 12664 10639
rect 13096 10606 13124 11766
rect 13188 11218 13216 12310
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13280 11898 13308 12174
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13280 11286 13308 11630
rect 13372 11354 13400 15506
rect 13636 15428 13688 15434
rect 13636 15370 13688 15376
rect 13648 14958 13676 15370
rect 13924 15162 13952 15506
rect 14066 15260 14362 15280
rect 14122 15258 14146 15260
rect 14202 15258 14226 15260
rect 14282 15258 14306 15260
rect 14144 15206 14146 15258
rect 14208 15206 14220 15258
rect 14282 15206 14284 15258
rect 14122 15204 14146 15206
rect 14202 15204 14226 15206
rect 14282 15204 14306 15206
rect 14066 15184 14362 15204
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13648 14090 13676 14894
rect 13912 14884 13964 14890
rect 13912 14826 13964 14832
rect 13648 14062 13768 14090
rect 13924 14074 13952 14826
rect 14066 14172 14362 14192
rect 14122 14170 14146 14172
rect 14202 14170 14226 14172
rect 14282 14170 14306 14172
rect 14144 14118 14146 14170
rect 14208 14118 14220 14170
rect 14282 14118 14284 14170
rect 14122 14116 14146 14118
rect 14202 14116 14226 14118
rect 14282 14116 14306 14118
rect 14066 14096 14362 14116
rect 13740 14006 13768 14062
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 13728 14000 13780 14006
rect 13728 13942 13780 13948
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 13740 11898 13768 13806
rect 14108 13530 14136 13806
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13924 12986 13952 13330
rect 14066 13084 14362 13104
rect 14122 13082 14146 13084
rect 14202 13082 14226 13084
rect 14282 13082 14306 13084
rect 14144 13030 14146 13082
rect 14208 13030 14220 13082
rect 14282 13030 14284 13082
rect 14122 13028 14146 13030
rect 14202 13028 14226 13030
rect 14282 13028 14306 13030
rect 14066 13008 14362 13028
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 14004 12776 14056 12782
rect 14280 12776 14332 12782
rect 14056 12724 14280 12730
rect 14004 12718 14332 12724
rect 14016 12702 14320 12718
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13268 11280 13320 11286
rect 13268 11222 13320 11228
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13280 11098 13308 11222
rect 13832 11218 13860 12038
rect 14066 11996 14362 12016
rect 14122 11994 14146 11996
rect 14202 11994 14226 11996
rect 14282 11994 14306 11996
rect 14144 11942 14146 11994
rect 14208 11942 14220 11994
rect 14282 11942 14284 11994
rect 14122 11940 14146 11942
rect 14202 11940 14226 11942
rect 14282 11940 14306 11942
rect 14066 11920 14362 11940
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 14292 11558 14320 11698
rect 14568 11626 14596 12106
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14004 11552 14056 11558
rect 14096 11552 14148 11558
rect 14056 11512 14096 11540
rect 14004 11494 14056 11500
rect 14096 11494 14148 11500
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14568 11218 14596 11562
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 13280 11070 13400 11098
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 12716 10600 12768 10606
rect 12636 10560 12716 10588
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 12268 9500 12296 9930
rect 12360 9654 12388 10066
rect 12636 10033 12664 10560
rect 12716 10542 12768 10548
rect 13084 10600 13136 10606
rect 13084 10542 13136 10548
rect 12716 10056 12768 10062
rect 12622 10024 12678 10033
rect 12716 9998 12768 10004
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 12622 9959 12678 9968
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12544 9722 12572 9862
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12348 9512 12400 9518
rect 12268 9472 12348 9500
rect 12268 7818 12296 9472
rect 12348 9454 12400 9460
rect 12636 9110 12664 9959
rect 12728 9722 12756 9998
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12624 9104 12676 9110
rect 12728 9092 12756 9658
rect 13096 9654 13124 9998
rect 13084 9648 13136 9654
rect 13084 9590 13136 9596
rect 13096 9518 13124 9590
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 12808 9104 12860 9110
rect 12728 9064 12808 9092
rect 12624 9046 12676 9052
rect 12808 9046 12860 9052
rect 13096 8090 13124 9454
rect 13188 9042 13216 9522
rect 13280 9518 13308 10950
rect 13372 10606 13400 11070
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 13372 10130 13400 10542
rect 13832 10130 13860 11154
rect 14066 10908 14362 10928
rect 14122 10906 14146 10908
rect 14202 10906 14226 10908
rect 14282 10906 14306 10908
rect 14144 10854 14146 10906
rect 14208 10854 14220 10906
rect 14282 10854 14284 10906
rect 14122 10852 14146 10854
rect 14202 10852 14226 10854
rect 14282 10852 14306 10854
rect 14066 10832 14362 10852
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13832 9654 13860 9862
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13924 9518 13952 9930
rect 14066 9820 14362 9840
rect 14122 9818 14146 9820
rect 14202 9818 14226 9820
rect 14282 9818 14306 9820
rect 14144 9766 14146 9818
rect 14208 9766 14220 9818
rect 14282 9766 14284 9818
rect 14122 9764 14146 9766
rect 14202 9764 14226 9766
rect 14282 9764 14306 9766
rect 14066 9744 14362 9764
rect 14476 9722 14504 10610
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14568 9602 14596 10066
rect 14476 9574 14596 9602
rect 14476 9518 14504 9574
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13372 9042 13400 9386
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13648 8906 13676 9454
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12268 7410 12296 7754
rect 12360 7750 12388 8026
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12360 7342 12388 7686
rect 12544 7546 12572 7822
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 10980 5098 11008 6190
rect 11444 6012 11740 6032
rect 11500 6010 11524 6012
rect 11580 6010 11604 6012
rect 11660 6010 11684 6012
rect 11522 5958 11524 6010
rect 11586 5958 11598 6010
rect 11660 5958 11662 6010
rect 11500 5956 11524 5958
rect 11580 5956 11604 5958
rect 11660 5956 11684 5958
rect 11444 5936 11740 5956
rect 12268 5846 12296 6598
rect 12360 6118 12388 7278
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12452 6934 12480 7142
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12544 6798 12572 7482
rect 12636 7342 12664 7890
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12898 7304 12954 7313
rect 12898 7239 12954 7248
rect 12912 7206 12940 7239
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12544 6458 12572 6734
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12912 6322 12940 6802
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12912 5914 12940 6258
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 12256 5840 12308 5846
rect 12256 5782 12308 5788
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 11256 4826 11284 5034
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11256 4078 11284 4626
rect 11348 4622 11376 5102
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11444 4924 11740 4944
rect 11500 4922 11524 4924
rect 11580 4922 11604 4924
rect 11660 4922 11684 4924
rect 11522 4870 11524 4922
rect 11586 4870 11598 4922
rect 11660 4870 11662 4922
rect 11500 4868 11524 4870
rect 11580 4868 11604 4870
rect 11660 4868 11684 4870
rect 11444 4848 11740 4868
rect 11808 4690 11836 4966
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 11164 3126 11192 3538
rect 11256 3466 11284 4014
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 11348 3194 11376 4558
rect 11900 4554 11928 5102
rect 12072 5092 12124 5098
rect 12072 5034 12124 5040
rect 12084 4690 12112 5034
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12728 4690 12756 4966
rect 13004 4690 13032 5102
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 12452 4214 12480 4558
rect 13004 4282 13032 4626
rect 12992 4276 13044 4282
rect 12992 4218 13044 4224
rect 12440 4208 12492 4214
rect 12440 4150 12492 4156
rect 12072 4072 12124 4078
rect 12440 4072 12492 4078
rect 12124 4032 12204 4060
rect 12072 4014 12124 4020
rect 11444 3836 11740 3856
rect 11500 3834 11524 3836
rect 11580 3834 11604 3836
rect 11660 3834 11684 3836
rect 11522 3782 11524 3834
rect 11586 3782 11598 3834
rect 11660 3782 11662 3834
rect 11500 3780 11524 3782
rect 11580 3780 11604 3782
rect 11660 3780 11684 3782
rect 11444 3760 11740 3780
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 11900 2990 11928 3674
rect 12176 3466 12204 4032
rect 12440 4014 12492 4020
rect 12348 4004 12400 4010
rect 12348 3946 12400 3952
rect 12360 3670 12388 3946
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 12176 2990 12204 3402
rect 12452 3398 12480 4014
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12452 3126 12480 3334
rect 13188 3194 13216 8366
rect 13452 8016 13504 8022
rect 13452 7958 13504 7964
rect 13464 7546 13492 7958
rect 13648 7732 13676 8842
rect 14066 8732 14362 8752
rect 14122 8730 14146 8732
rect 14202 8730 14226 8732
rect 14282 8730 14306 8732
rect 14144 8678 14146 8730
rect 14208 8678 14220 8730
rect 14282 8678 14284 8730
rect 14122 8676 14146 8678
rect 14202 8676 14226 8678
rect 14282 8676 14306 8678
rect 14066 8656 14362 8676
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13740 7954 13768 8026
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13556 7704 13676 7732
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13556 7342 13584 7704
rect 13832 7410 13860 8230
rect 13924 8090 13952 8366
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13924 7410 13952 8026
rect 14568 7954 14596 9318
rect 14660 9178 14688 10542
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14066 7644 14362 7664
rect 14122 7642 14146 7644
rect 14202 7642 14226 7644
rect 14282 7642 14306 7644
rect 14144 7590 14146 7642
rect 14208 7590 14220 7642
rect 14282 7590 14284 7642
rect 14122 7588 14146 7590
rect 14202 7588 14226 7590
rect 14282 7588 14306 7590
rect 14066 7568 14362 7588
rect 14568 7426 14596 7686
rect 14660 7546 14688 9114
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 14384 7398 14596 7426
rect 14384 7342 14412 7398
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 13556 7002 13584 7278
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13372 6458 13400 6802
rect 14660 6798 14688 7482
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13464 6390 13492 6734
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13452 6384 13504 6390
rect 13452 6326 13504 6332
rect 13464 6254 13492 6326
rect 13832 6322 13860 6598
rect 14066 6556 14362 6576
rect 14122 6554 14146 6556
rect 14202 6554 14226 6556
rect 14282 6554 14306 6556
rect 14144 6502 14146 6554
rect 14208 6502 14220 6554
rect 14282 6502 14284 6554
rect 14122 6500 14146 6502
rect 14202 6500 14226 6502
rect 14282 6500 14306 6502
rect 14066 6480 14362 6500
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 13452 6248 13504 6254
rect 13452 6190 13504 6196
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13268 5840 13320 5846
rect 13268 5782 13320 5788
rect 13280 5370 13308 5782
rect 13832 5710 13860 6054
rect 14476 5778 14504 6258
rect 14556 6180 14608 6186
rect 14556 6122 14608 6128
rect 14568 5914 14596 6122
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 13832 4570 13860 5646
rect 14066 5468 14362 5488
rect 14122 5466 14146 5468
rect 14202 5466 14226 5468
rect 14282 5466 14306 5468
rect 14144 5414 14146 5466
rect 14208 5414 14220 5466
rect 14282 5414 14284 5466
rect 14122 5412 14146 5414
rect 14202 5412 14226 5414
rect 14282 5412 14306 5414
rect 14066 5392 14362 5412
rect 14476 4690 14504 5714
rect 14752 4758 14780 16546
rect 14924 16176 14976 16182
rect 14924 16118 14976 16124
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14844 13802 14872 14010
rect 14832 13796 14884 13802
rect 14832 13738 14884 13744
rect 14844 12782 14872 13738
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 14844 11694 14872 12310
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14844 7886 14872 11630
rect 14936 11082 14964 16118
rect 16486 15736 16542 15745
rect 16486 15671 16542 15680
rect 16500 15570 16528 15671
rect 15752 15564 15804 15570
rect 15752 15506 15804 15512
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 15764 15162 15792 15506
rect 15844 15360 15896 15366
rect 15844 15302 15896 15308
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15120 12850 15148 13262
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 15120 11762 15148 12786
rect 15212 11898 15240 14894
rect 15764 14822 15792 15098
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15856 14006 15884 15302
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15396 12986 15424 13806
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15764 12442 15792 12582
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15120 11218 15148 11698
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14924 10464 14976 10470
rect 14924 10406 14976 10412
rect 14936 10198 14964 10406
rect 14924 10192 14976 10198
rect 14924 10134 14976 10140
rect 14924 10056 14976 10062
rect 15580 10033 15608 12242
rect 15752 11688 15804 11694
rect 15750 11656 15752 11665
rect 15804 11656 15806 11665
rect 15750 11591 15806 11600
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 14924 9998 14976 10004
rect 15566 10024 15622 10033
rect 14936 8974 14964 9998
rect 15566 9959 15622 9968
rect 15568 9512 15620 9518
rect 15672 9500 15700 10542
rect 15620 9472 15700 9500
rect 15568 9454 15620 9460
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14936 8242 14964 8910
rect 14936 8214 15148 8242
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14844 7426 14872 7686
rect 14844 7410 14964 7426
rect 14844 7404 14976 7410
rect 14844 7398 14924 7404
rect 14844 6118 14872 7398
rect 14924 7346 14976 7352
rect 15028 7206 15056 7890
rect 15120 7750 15148 8214
rect 15580 7936 15608 9454
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15672 9110 15700 9318
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15660 7948 15712 7954
rect 15580 7908 15660 7936
rect 15660 7890 15712 7896
rect 15108 7744 15160 7750
rect 15108 7686 15160 7692
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15304 6458 15332 6802
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15672 6322 15700 7890
rect 15764 6458 15792 11494
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14844 5914 14872 6054
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 14740 4752 14792 4758
rect 14740 4694 14792 4700
rect 14464 4684 14516 4690
rect 14516 4644 14688 4672
rect 14464 4626 14516 4632
rect 13740 4542 13860 4570
rect 13740 4146 13768 4542
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13832 3942 13860 4422
rect 14066 4380 14362 4400
rect 14122 4378 14146 4380
rect 14202 4378 14226 4380
rect 14282 4378 14306 4380
rect 14144 4326 14146 4378
rect 14208 4326 14220 4378
rect 14282 4326 14284 4378
rect 14122 4324 14146 4326
rect 14202 4324 14226 4326
rect 14282 4324 14306 4326
rect 14066 4304 14362 4324
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14476 3602 14504 3878
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14066 3292 14362 3312
rect 14122 3290 14146 3292
rect 14202 3290 14226 3292
rect 14282 3290 14306 3292
rect 14144 3238 14146 3290
rect 14208 3238 14220 3290
rect 14282 3238 14284 3290
rect 14122 3236 14146 3238
rect 14202 3236 14226 3238
rect 14282 3236 14306 3238
rect 14066 3216 14362 3236
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8576 2984 8628 2990
rect 8760 2984 8812 2990
rect 8576 2926 8628 2932
rect 8758 2952 8760 2961
rect 8944 2984 8996 2990
rect 8812 2952 8814 2961
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8588 2514 8616 2926
rect 8944 2926 8996 2932
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10324 2984 10376 2990
rect 10324 2926 10376 2932
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 8758 2887 8814 2896
rect 8956 2582 8984 2926
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 9600 2582 9628 2790
rect 10244 2582 10272 2790
rect 8944 2576 8996 2582
rect 8944 2518 8996 2524
rect 9588 2576 9640 2582
rect 9588 2518 9640 2524
rect 10232 2576 10284 2582
rect 10232 2518 10284 2524
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8024 2372 8076 2378
rect 8024 2314 8076 2320
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 7748 2100 7800 2106
rect 7748 2042 7800 2048
rect 8312 800 8340 2450
rect 8822 2204 9118 2224
rect 8878 2202 8902 2204
rect 8958 2202 8982 2204
rect 9038 2202 9062 2204
rect 8900 2150 8902 2202
rect 8964 2150 8976 2202
rect 9038 2150 9040 2202
rect 8878 2148 8902 2150
rect 8958 2148 8982 2150
rect 9038 2148 9062 2150
rect 8822 2128 9118 2148
rect 10336 1578 10364 2926
rect 11444 2748 11740 2768
rect 11500 2746 11524 2748
rect 11580 2746 11604 2748
rect 11660 2746 11684 2748
rect 11522 2694 11524 2746
rect 11586 2694 11598 2746
rect 11660 2694 11662 2746
rect 11500 2692 11524 2694
rect 11580 2692 11604 2694
rect 11660 2692 11684 2694
rect 11444 2672 11740 2692
rect 11808 2650 11836 2926
rect 11980 2916 12032 2922
rect 11980 2858 12032 2864
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 11992 2514 12020 2858
rect 12728 2650 12756 2858
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 10152 1550 10364 1578
rect 10152 800 10180 1550
rect 11532 800 11560 2450
rect 13372 800 13400 2926
rect 14108 2446 14136 3062
rect 14568 3058 14596 4082
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14568 2514 14596 2994
rect 14660 2514 14688 4644
rect 14844 4282 14872 5510
rect 15200 4548 15252 4554
rect 15200 4490 15252 4496
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 15212 2650 15240 4490
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15580 4010 15608 4422
rect 15568 4004 15620 4010
rect 15568 3946 15620 3952
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 15580 3466 15608 3538
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 15580 3058 15608 3402
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 15764 2650 15792 2858
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14066 2204 14362 2224
rect 14122 2202 14146 2204
rect 14202 2202 14226 2204
rect 14282 2202 14306 2204
rect 14144 2150 14146 2202
rect 14208 2150 14220 2202
rect 14282 2150 14284 2202
rect 14122 2148 14146 2150
rect 14202 2148 14226 2150
rect 14282 2148 14306 2150
rect 14066 2128 14362 2148
rect 15212 800 15240 2450
rect 15856 2378 15884 11222
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15948 10198 15976 10406
rect 15936 10192 15988 10198
rect 15936 10134 15988 10140
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 15948 7274 15976 7686
rect 15936 7268 15988 7274
rect 15936 7210 15988 7216
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15948 5846 15976 6054
rect 15936 5840 15988 5846
rect 15936 5782 15988 5788
rect 16040 2650 16068 11494
rect 16224 11354 16252 13398
rect 16316 12782 16344 14214
rect 16500 13705 16528 14418
rect 16486 13696 16542 13705
rect 16486 13631 16542 13640
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16500 10985 16528 11154
rect 16486 10976 16542 10985
rect 16486 10911 16542 10920
rect 16302 10024 16358 10033
rect 16302 9959 16358 9968
rect 16316 9178 16344 9959
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16304 8288 16356 8294
rect 16500 8265 16528 8366
rect 16304 8230 16356 8236
rect 16486 8256 16542 8265
rect 16316 5846 16344 8230
rect 16486 8191 16542 8200
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 16408 7546 16436 7754
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16488 6248 16540 6254
rect 16486 6216 16488 6225
rect 16540 6216 16542 6225
rect 16486 6151 16542 6160
rect 16304 5840 16356 5846
rect 16304 5782 16356 5788
rect 16488 4684 16540 4690
rect 16488 4626 16540 4632
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16316 3194 16344 3538
rect 16408 3534 16436 3878
rect 16396 3528 16448 3534
rect 16500 3505 16528 4626
rect 16396 3470 16448 3476
rect 16486 3496 16542 3505
rect 16486 3431 16542 3440
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16028 2644 16080 2650
rect 16028 2586 16080 2592
rect 16488 2508 16540 2514
rect 16488 2450 16540 2456
rect 15844 2372 15896 2378
rect 15844 2314 15896 2320
rect 16500 1465 16528 2450
rect 16580 2440 16632 2446
rect 16580 2382 16632 2388
rect 16486 1456 16542 1465
rect 16486 1391 16542 1400
rect 16592 800 16620 2382
rect 478 0 534 800
rect 1858 0 1914 800
rect 3698 0 3754 800
rect 5078 0 5134 800
rect 6918 0 6974 800
rect 8298 0 8354 800
rect 10138 0 10194 800
rect 11518 0 11574 800
rect 13358 0 13414 800
rect 15198 0 15254 800
rect 16578 0 16634 800
<< via2 >>
rect 1398 17076 1400 17096
rect 1400 17076 1452 17096
rect 1452 17076 1454 17096
rect 1398 17040 1454 17076
rect 3578 17434 3634 17436
rect 3658 17434 3714 17436
rect 3738 17434 3794 17436
rect 3818 17434 3874 17436
rect 3578 17382 3604 17434
rect 3604 17382 3634 17434
rect 3658 17382 3668 17434
rect 3668 17382 3714 17434
rect 3738 17382 3784 17434
rect 3784 17382 3794 17434
rect 3818 17382 3848 17434
rect 3848 17382 3874 17434
rect 3578 17380 3634 17382
rect 3658 17380 3714 17382
rect 3738 17380 3794 17382
rect 3818 17380 3874 17382
rect 1398 15000 1454 15056
rect 1398 12300 1454 12336
rect 1398 12280 1400 12300
rect 1400 12280 1452 12300
rect 1452 12280 1454 12300
rect 1582 12164 1638 12200
rect 1582 12144 1584 12164
rect 1584 12144 1636 12164
rect 1636 12144 1638 12164
rect 1398 10240 1454 10296
rect 1398 7520 1454 7576
rect 1398 5480 1454 5536
rect 3578 16346 3634 16348
rect 3658 16346 3714 16348
rect 3738 16346 3794 16348
rect 3818 16346 3874 16348
rect 3578 16294 3604 16346
rect 3604 16294 3634 16346
rect 3658 16294 3668 16346
rect 3668 16294 3714 16346
rect 3738 16294 3784 16346
rect 3784 16294 3794 16346
rect 3818 16294 3848 16346
rect 3848 16294 3874 16346
rect 3578 16292 3634 16294
rect 3658 16292 3714 16294
rect 3738 16292 3794 16294
rect 3818 16292 3874 16294
rect 3578 15258 3634 15260
rect 3658 15258 3714 15260
rect 3738 15258 3794 15260
rect 3818 15258 3874 15260
rect 3578 15206 3604 15258
rect 3604 15206 3634 15258
rect 3658 15206 3668 15258
rect 3668 15206 3714 15258
rect 3738 15206 3784 15258
rect 3784 15206 3794 15258
rect 3818 15206 3848 15258
rect 3848 15206 3874 15258
rect 3578 15204 3634 15206
rect 3658 15204 3714 15206
rect 3738 15204 3794 15206
rect 3818 15204 3874 15206
rect 6200 17978 6256 17980
rect 6280 17978 6336 17980
rect 6360 17978 6416 17980
rect 6440 17978 6496 17980
rect 6200 17926 6226 17978
rect 6226 17926 6256 17978
rect 6280 17926 6290 17978
rect 6290 17926 6336 17978
rect 6360 17926 6406 17978
rect 6406 17926 6416 17978
rect 6440 17926 6470 17978
rect 6470 17926 6496 17978
rect 6200 17924 6256 17926
rect 6280 17924 6336 17926
rect 6360 17924 6416 17926
rect 6440 17924 6496 17926
rect 11444 17978 11500 17980
rect 11524 17978 11580 17980
rect 11604 17978 11660 17980
rect 11684 17978 11740 17980
rect 11444 17926 11470 17978
rect 11470 17926 11500 17978
rect 11524 17926 11534 17978
rect 11534 17926 11580 17978
rect 11604 17926 11650 17978
rect 11650 17926 11660 17978
rect 11684 17926 11714 17978
rect 11714 17926 11740 17978
rect 11444 17924 11500 17926
rect 11524 17924 11580 17926
rect 11604 17924 11660 17926
rect 11684 17924 11740 17926
rect 16118 18400 16174 18456
rect 3578 14170 3634 14172
rect 3658 14170 3714 14172
rect 3738 14170 3794 14172
rect 3818 14170 3874 14172
rect 3578 14118 3604 14170
rect 3604 14118 3634 14170
rect 3658 14118 3668 14170
rect 3668 14118 3714 14170
rect 3738 14118 3784 14170
rect 3784 14118 3794 14170
rect 3818 14118 3848 14170
rect 3848 14118 3874 14170
rect 3578 14116 3634 14118
rect 3658 14116 3714 14118
rect 3738 14116 3794 14118
rect 3818 14116 3874 14118
rect 3882 13388 3938 13424
rect 3882 13368 3884 13388
rect 3884 13368 3936 13388
rect 3936 13368 3938 13388
rect 3578 13082 3634 13084
rect 3658 13082 3714 13084
rect 3738 13082 3794 13084
rect 3818 13082 3874 13084
rect 3578 13030 3604 13082
rect 3604 13030 3634 13082
rect 3658 13030 3668 13082
rect 3668 13030 3714 13082
rect 3738 13030 3784 13082
rect 3784 13030 3794 13082
rect 3818 13030 3848 13082
rect 3848 13030 3874 13082
rect 3578 13028 3634 13030
rect 3658 13028 3714 13030
rect 3738 13028 3794 13030
rect 3818 13028 3874 13030
rect 5170 13388 5226 13424
rect 5170 13368 5172 13388
rect 5172 13368 5224 13388
rect 5224 13368 5226 13388
rect 3578 11994 3634 11996
rect 3658 11994 3714 11996
rect 3738 11994 3794 11996
rect 3818 11994 3874 11996
rect 3578 11942 3604 11994
rect 3604 11942 3634 11994
rect 3658 11942 3668 11994
rect 3668 11942 3714 11994
rect 3738 11942 3784 11994
rect 3784 11942 3794 11994
rect 3818 11942 3848 11994
rect 3848 11942 3874 11994
rect 3578 11940 3634 11942
rect 3658 11940 3714 11942
rect 3738 11940 3794 11942
rect 3818 11940 3874 11942
rect 1398 2760 1454 2816
rect 3578 10906 3634 10908
rect 3658 10906 3714 10908
rect 3738 10906 3794 10908
rect 3818 10906 3874 10908
rect 3578 10854 3604 10906
rect 3604 10854 3634 10906
rect 3658 10854 3668 10906
rect 3668 10854 3714 10906
rect 3738 10854 3784 10906
rect 3784 10854 3794 10906
rect 3818 10854 3848 10906
rect 3848 10854 3874 10906
rect 3578 10852 3634 10854
rect 3658 10852 3714 10854
rect 3738 10852 3794 10854
rect 3818 10852 3874 10854
rect 3578 9818 3634 9820
rect 3658 9818 3714 9820
rect 3738 9818 3794 9820
rect 3818 9818 3874 9820
rect 3578 9766 3604 9818
rect 3604 9766 3634 9818
rect 3658 9766 3668 9818
rect 3668 9766 3714 9818
rect 3738 9766 3784 9818
rect 3784 9766 3794 9818
rect 3818 9766 3848 9818
rect 3848 9766 3874 9818
rect 3578 9764 3634 9766
rect 3658 9764 3714 9766
rect 3738 9764 3794 9766
rect 3818 9764 3874 9766
rect 3578 8730 3634 8732
rect 3658 8730 3714 8732
rect 3738 8730 3794 8732
rect 3818 8730 3874 8732
rect 3578 8678 3604 8730
rect 3604 8678 3634 8730
rect 3658 8678 3668 8730
rect 3668 8678 3714 8730
rect 3738 8678 3784 8730
rect 3784 8678 3794 8730
rect 3818 8678 3848 8730
rect 3848 8678 3874 8730
rect 3578 8676 3634 8678
rect 3658 8676 3714 8678
rect 3738 8676 3794 8678
rect 3818 8676 3874 8678
rect 6200 16890 6256 16892
rect 6280 16890 6336 16892
rect 6360 16890 6416 16892
rect 6440 16890 6496 16892
rect 6200 16838 6226 16890
rect 6226 16838 6256 16890
rect 6280 16838 6290 16890
rect 6290 16838 6336 16890
rect 6360 16838 6406 16890
rect 6406 16838 6416 16890
rect 6440 16838 6470 16890
rect 6470 16838 6496 16890
rect 6200 16836 6256 16838
rect 6280 16836 6336 16838
rect 6360 16836 6416 16838
rect 6440 16836 6496 16838
rect 3578 7642 3634 7644
rect 3658 7642 3714 7644
rect 3738 7642 3794 7644
rect 3818 7642 3874 7644
rect 3578 7590 3604 7642
rect 3604 7590 3634 7642
rect 3658 7590 3668 7642
rect 3668 7590 3714 7642
rect 3738 7590 3784 7642
rect 3784 7590 3794 7642
rect 3818 7590 3848 7642
rect 3848 7590 3874 7642
rect 3578 7588 3634 7590
rect 3658 7588 3714 7590
rect 3738 7588 3794 7590
rect 3818 7588 3874 7590
rect 3578 6554 3634 6556
rect 3658 6554 3714 6556
rect 3738 6554 3794 6556
rect 3818 6554 3874 6556
rect 3578 6502 3604 6554
rect 3604 6502 3634 6554
rect 3658 6502 3668 6554
rect 3668 6502 3714 6554
rect 3738 6502 3784 6554
rect 3784 6502 3794 6554
rect 3818 6502 3848 6554
rect 3848 6502 3874 6554
rect 3578 6500 3634 6502
rect 3658 6500 3714 6502
rect 3738 6500 3794 6502
rect 3818 6500 3874 6502
rect 3578 5466 3634 5468
rect 3658 5466 3714 5468
rect 3738 5466 3794 5468
rect 3818 5466 3874 5468
rect 3578 5414 3604 5466
rect 3604 5414 3634 5466
rect 3658 5414 3668 5466
rect 3668 5414 3714 5466
rect 3738 5414 3784 5466
rect 3784 5414 3794 5466
rect 3818 5414 3848 5466
rect 3848 5414 3874 5466
rect 3578 5412 3634 5414
rect 3658 5412 3714 5414
rect 3738 5412 3794 5414
rect 3818 5412 3874 5414
rect 3578 4378 3634 4380
rect 3658 4378 3714 4380
rect 3738 4378 3794 4380
rect 3818 4378 3874 4380
rect 3578 4326 3604 4378
rect 3604 4326 3634 4378
rect 3658 4326 3668 4378
rect 3668 4326 3714 4378
rect 3738 4326 3784 4378
rect 3784 4326 3794 4378
rect 3818 4326 3848 4378
rect 3848 4326 3874 4378
rect 3578 4324 3634 4326
rect 3658 4324 3714 4326
rect 3738 4324 3794 4326
rect 3818 4324 3874 4326
rect 3578 3290 3634 3292
rect 3658 3290 3714 3292
rect 3738 3290 3794 3292
rect 3818 3290 3874 3292
rect 3578 3238 3604 3290
rect 3604 3238 3634 3290
rect 3658 3238 3668 3290
rect 3668 3238 3714 3290
rect 3738 3238 3784 3290
rect 3784 3238 3794 3290
rect 3818 3238 3848 3290
rect 3848 3238 3874 3290
rect 3578 3236 3634 3238
rect 3658 3236 3714 3238
rect 3738 3236 3794 3238
rect 3818 3236 3874 3238
rect 3578 2202 3634 2204
rect 3658 2202 3714 2204
rect 3738 2202 3794 2204
rect 3818 2202 3874 2204
rect 3578 2150 3604 2202
rect 3604 2150 3634 2202
rect 3658 2150 3668 2202
rect 3668 2150 3714 2202
rect 3738 2150 3784 2202
rect 3784 2150 3794 2202
rect 3818 2150 3848 2202
rect 3848 2150 3874 2202
rect 3578 2148 3634 2150
rect 3658 2148 3714 2150
rect 3738 2148 3794 2150
rect 3818 2148 3874 2150
rect 6200 15802 6256 15804
rect 6280 15802 6336 15804
rect 6360 15802 6416 15804
rect 6440 15802 6496 15804
rect 6200 15750 6226 15802
rect 6226 15750 6256 15802
rect 6280 15750 6290 15802
rect 6290 15750 6336 15802
rect 6360 15750 6406 15802
rect 6406 15750 6416 15802
rect 6440 15750 6470 15802
rect 6470 15750 6496 15802
rect 6200 15748 6256 15750
rect 6280 15748 6336 15750
rect 6360 15748 6416 15750
rect 6440 15748 6496 15750
rect 6200 14714 6256 14716
rect 6280 14714 6336 14716
rect 6360 14714 6416 14716
rect 6440 14714 6496 14716
rect 6200 14662 6226 14714
rect 6226 14662 6256 14714
rect 6280 14662 6290 14714
rect 6290 14662 6336 14714
rect 6360 14662 6406 14714
rect 6406 14662 6416 14714
rect 6440 14662 6470 14714
rect 6470 14662 6496 14714
rect 6200 14660 6256 14662
rect 6280 14660 6336 14662
rect 6360 14660 6416 14662
rect 6440 14660 6496 14662
rect 6182 14476 6238 14512
rect 6182 14456 6184 14476
rect 6184 14456 6236 14476
rect 6236 14456 6238 14476
rect 5998 14340 6054 14376
rect 5998 14320 6000 14340
rect 6000 14320 6052 14340
rect 6052 14320 6054 14340
rect 6200 13626 6256 13628
rect 6280 13626 6336 13628
rect 6360 13626 6416 13628
rect 6440 13626 6496 13628
rect 6200 13574 6226 13626
rect 6226 13574 6256 13626
rect 6280 13574 6290 13626
rect 6290 13574 6336 13626
rect 6360 13574 6406 13626
rect 6406 13574 6416 13626
rect 6440 13574 6470 13626
rect 6470 13574 6496 13626
rect 6200 13572 6256 13574
rect 6280 13572 6336 13574
rect 6360 13572 6416 13574
rect 6440 13572 6496 13574
rect 6642 14356 6644 14376
rect 6644 14356 6696 14376
rect 6696 14356 6698 14376
rect 6642 14320 6698 14356
rect 6918 14476 6974 14512
rect 6918 14456 6920 14476
rect 6920 14456 6972 14476
rect 6972 14456 6974 14476
rect 6200 12538 6256 12540
rect 6280 12538 6336 12540
rect 6360 12538 6416 12540
rect 6440 12538 6496 12540
rect 6200 12486 6226 12538
rect 6226 12486 6256 12538
rect 6280 12486 6290 12538
rect 6290 12486 6336 12538
rect 6360 12486 6406 12538
rect 6406 12486 6416 12538
rect 6440 12486 6470 12538
rect 6470 12486 6496 12538
rect 6200 12484 6256 12486
rect 6280 12484 6336 12486
rect 6360 12484 6416 12486
rect 6440 12484 6496 12486
rect 6200 11450 6256 11452
rect 6280 11450 6336 11452
rect 6360 11450 6416 11452
rect 6440 11450 6496 11452
rect 6200 11398 6226 11450
rect 6226 11398 6256 11450
rect 6280 11398 6290 11450
rect 6290 11398 6336 11450
rect 6360 11398 6406 11450
rect 6406 11398 6416 11450
rect 6440 11398 6470 11450
rect 6470 11398 6496 11450
rect 6200 11396 6256 11398
rect 6280 11396 6336 11398
rect 6360 11396 6416 11398
rect 6440 11396 6496 11398
rect 6200 10362 6256 10364
rect 6280 10362 6336 10364
rect 6360 10362 6416 10364
rect 6440 10362 6496 10364
rect 6200 10310 6226 10362
rect 6226 10310 6256 10362
rect 6280 10310 6290 10362
rect 6290 10310 6336 10362
rect 6360 10310 6406 10362
rect 6406 10310 6416 10362
rect 6440 10310 6470 10362
rect 6470 10310 6496 10362
rect 6200 10308 6256 10310
rect 6280 10308 6336 10310
rect 6360 10308 6416 10310
rect 6440 10308 6496 10310
rect 8822 17434 8878 17436
rect 8902 17434 8958 17436
rect 8982 17434 9038 17436
rect 9062 17434 9118 17436
rect 8822 17382 8848 17434
rect 8848 17382 8878 17434
rect 8902 17382 8912 17434
rect 8912 17382 8958 17434
rect 8982 17382 9028 17434
rect 9028 17382 9038 17434
rect 9062 17382 9092 17434
rect 9092 17382 9118 17434
rect 8822 17380 8878 17382
rect 8902 17380 8958 17382
rect 8982 17380 9038 17382
rect 9062 17380 9118 17382
rect 8822 16346 8878 16348
rect 8902 16346 8958 16348
rect 8982 16346 9038 16348
rect 9062 16346 9118 16348
rect 8822 16294 8848 16346
rect 8848 16294 8878 16346
rect 8902 16294 8912 16346
rect 8912 16294 8958 16346
rect 8982 16294 9028 16346
rect 9028 16294 9038 16346
rect 9062 16294 9092 16346
rect 9092 16294 9118 16346
rect 8822 16292 8878 16294
rect 8902 16292 8958 16294
rect 8982 16292 9038 16294
rect 9062 16292 9118 16294
rect 11444 16890 11500 16892
rect 11524 16890 11580 16892
rect 11604 16890 11660 16892
rect 11684 16890 11740 16892
rect 11444 16838 11470 16890
rect 11470 16838 11500 16890
rect 11524 16838 11534 16890
rect 11534 16838 11580 16890
rect 11604 16838 11650 16890
rect 11650 16838 11660 16890
rect 11684 16838 11714 16890
rect 11714 16838 11740 16890
rect 11444 16836 11500 16838
rect 11524 16836 11580 16838
rect 11604 16836 11660 16838
rect 11684 16836 11740 16838
rect 8822 15258 8878 15260
rect 8902 15258 8958 15260
rect 8982 15258 9038 15260
rect 9062 15258 9118 15260
rect 8822 15206 8848 15258
rect 8848 15206 8878 15258
rect 8902 15206 8912 15258
rect 8912 15206 8958 15258
rect 8982 15206 9028 15258
rect 9028 15206 9038 15258
rect 9062 15206 9092 15258
rect 9092 15206 9118 15258
rect 8822 15204 8878 15206
rect 8902 15204 8958 15206
rect 8982 15204 9038 15206
rect 9062 15204 9118 15206
rect 11444 15802 11500 15804
rect 11524 15802 11580 15804
rect 11604 15802 11660 15804
rect 11684 15802 11740 15804
rect 11444 15750 11470 15802
rect 11470 15750 11500 15802
rect 11524 15750 11534 15802
rect 11534 15750 11580 15802
rect 11604 15750 11650 15802
rect 11650 15750 11660 15802
rect 11684 15750 11714 15802
rect 11714 15750 11740 15802
rect 11444 15748 11500 15750
rect 11524 15748 11580 15750
rect 11604 15748 11660 15750
rect 11684 15748 11740 15750
rect 8822 14170 8878 14172
rect 8902 14170 8958 14172
rect 8982 14170 9038 14172
rect 9062 14170 9118 14172
rect 8822 14118 8848 14170
rect 8848 14118 8878 14170
rect 8902 14118 8912 14170
rect 8912 14118 8958 14170
rect 8982 14118 9028 14170
rect 9028 14118 9038 14170
rect 9062 14118 9092 14170
rect 9092 14118 9118 14170
rect 8822 14116 8878 14118
rect 8902 14116 8958 14118
rect 8982 14116 9038 14118
rect 9062 14116 9118 14118
rect 11444 14714 11500 14716
rect 11524 14714 11580 14716
rect 11604 14714 11660 14716
rect 11684 14714 11740 14716
rect 11444 14662 11470 14714
rect 11470 14662 11500 14714
rect 11524 14662 11534 14714
rect 11534 14662 11580 14714
rect 11604 14662 11650 14714
rect 11650 14662 11660 14714
rect 11684 14662 11714 14714
rect 11714 14662 11740 14714
rect 11444 14660 11500 14662
rect 11524 14660 11580 14662
rect 11604 14660 11660 14662
rect 11684 14660 11740 14662
rect 11444 13626 11500 13628
rect 11524 13626 11580 13628
rect 11604 13626 11660 13628
rect 11684 13626 11740 13628
rect 11444 13574 11470 13626
rect 11470 13574 11500 13626
rect 11524 13574 11534 13626
rect 11534 13574 11580 13626
rect 11604 13574 11650 13626
rect 11650 13574 11660 13626
rect 11684 13574 11714 13626
rect 11714 13574 11740 13626
rect 11444 13572 11500 13574
rect 11524 13572 11580 13574
rect 11604 13572 11660 13574
rect 11684 13572 11740 13574
rect 7194 10548 7196 10568
rect 7196 10548 7248 10568
rect 7248 10548 7250 10568
rect 7194 10512 7250 10548
rect 6200 9274 6256 9276
rect 6280 9274 6336 9276
rect 6360 9274 6416 9276
rect 6440 9274 6496 9276
rect 6200 9222 6226 9274
rect 6226 9222 6256 9274
rect 6280 9222 6290 9274
rect 6290 9222 6336 9274
rect 6360 9222 6406 9274
rect 6406 9222 6416 9274
rect 6440 9222 6470 9274
rect 6470 9222 6496 9274
rect 6200 9220 6256 9222
rect 6280 9220 6336 9222
rect 6360 9220 6416 9222
rect 6440 9220 6496 9222
rect 6200 8186 6256 8188
rect 6280 8186 6336 8188
rect 6360 8186 6416 8188
rect 6440 8186 6496 8188
rect 6200 8134 6226 8186
rect 6226 8134 6256 8186
rect 6280 8134 6290 8186
rect 6290 8134 6336 8186
rect 6360 8134 6406 8186
rect 6406 8134 6416 8186
rect 6440 8134 6470 8186
rect 6470 8134 6496 8186
rect 6200 8132 6256 8134
rect 6280 8132 6336 8134
rect 6360 8132 6416 8134
rect 6440 8132 6496 8134
rect 6200 7098 6256 7100
rect 6280 7098 6336 7100
rect 6360 7098 6416 7100
rect 6440 7098 6496 7100
rect 6200 7046 6226 7098
rect 6226 7046 6256 7098
rect 6280 7046 6290 7098
rect 6290 7046 6336 7098
rect 6360 7046 6406 7098
rect 6406 7046 6416 7098
rect 6440 7046 6470 7098
rect 6470 7046 6496 7098
rect 6200 7044 6256 7046
rect 6280 7044 6336 7046
rect 6360 7044 6416 7046
rect 6440 7044 6496 7046
rect 6200 6010 6256 6012
rect 6280 6010 6336 6012
rect 6360 6010 6416 6012
rect 6440 6010 6496 6012
rect 6200 5958 6226 6010
rect 6226 5958 6256 6010
rect 6280 5958 6290 6010
rect 6290 5958 6336 6010
rect 6360 5958 6406 6010
rect 6406 5958 6416 6010
rect 6440 5958 6470 6010
rect 6470 5958 6496 6010
rect 6200 5956 6256 5958
rect 6280 5956 6336 5958
rect 6360 5956 6416 5958
rect 6440 5956 6496 5958
rect 6200 4922 6256 4924
rect 6280 4922 6336 4924
rect 6360 4922 6416 4924
rect 6440 4922 6496 4924
rect 6200 4870 6226 4922
rect 6226 4870 6256 4922
rect 6280 4870 6290 4922
rect 6290 4870 6336 4922
rect 6360 4870 6406 4922
rect 6406 4870 6416 4922
rect 6440 4870 6470 4922
rect 6470 4870 6496 4922
rect 6200 4868 6256 4870
rect 6280 4868 6336 4870
rect 6360 4868 6416 4870
rect 6440 4868 6496 4870
rect 6200 3834 6256 3836
rect 6280 3834 6336 3836
rect 6360 3834 6416 3836
rect 6440 3834 6496 3836
rect 6200 3782 6226 3834
rect 6226 3782 6256 3834
rect 6280 3782 6290 3834
rect 6290 3782 6336 3834
rect 6360 3782 6406 3834
rect 6406 3782 6416 3834
rect 6440 3782 6470 3834
rect 6470 3782 6496 3834
rect 6200 3780 6256 3782
rect 6280 3780 6336 3782
rect 6360 3780 6416 3782
rect 6440 3780 6496 3782
rect 7010 2896 7066 2952
rect 6200 2746 6256 2748
rect 6280 2746 6336 2748
rect 6360 2746 6416 2748
rect 6440 2746 6496 2748
rect 6200 2694 6226 2746
rect 6226 2694 6256 2746
rect 6280 2694 6290 2746
rect 6290 2694 6336 2746
rect 6360 2694 6406 2746
rect 6406 2694 6416 2746
rect 6440 2694 6470 2746
rect 6470 2694 6496 2746
rect 6200 2692 6256 2694
rect 6280 2692 6336 2694
rect 6360 2692 6416 2694
rect 6440 2692 6496 2694
rect 8822 13082 8878 13084
rect 8902 13082 8958 13084
rect 8982 13082 9038 13084
rect 9062 13082 9118 13084
rect 8822 13030 8848 13082
rect 8848 13030 8878 13082
rect 8902 13030 8912 13082
rect 8912 13030 8958 13082
rect 8982 13030 9028 13082
rect 9028 13030 9038 13082
rect 9062 13030 9092 13082
rect 9092 13030 9118 13082
rect 8822 13028 8878 13030
rect 8902 13028 8958 13030
rect 8982 13028 9038 13030
rect 9062 13028 9118 13030
rect 8390 12180 8392 12200
rect 8392 12180 8444 12200
rect 8444 12180 8446 12200
rect 8390 12144 8446 12180
rect 9402 12008 9458 12064
rect 8822 11994 8878 11996
rect 8902 11994 8958 11996
rect 8982 11994 9038 11996
rect 9062 11994 9118 11996
rect 8822 11942 8848 11994
rect 8848 11942 8878 11994
rect 8902 11942 8912 11994
rect 8912 11942 8958 11994
rect 8982 11942 9028 11994
rect 9028 11942 9038 11994
rect 9062 11942 9092 11994
rect 9092 11942 9118 11994
rect 8822 11940 8878 11942
rect 8902 11940 8958 11942
rect 8982 11940 9038 11942
rect 9062 11940 9118 11942
rect 8850 11464 8906 11520
rect 8822 10906 8878 10908
rect 8902 10906 8958 10908
rect 8982 10906 9038 10908
rect 9062 10906 9118 10908
rect 8822 10854 8848 10906
rect 8848 10854 8878 10906
rect 8902 10854 8912 10906
rect 8912 10854 8958 10906
rect 8982 10854 9028 10906
rect 9028 10854 9038 10906
rect 9062 10854 9092 10906
rect 9092 10854 9118 10906
rect 8822 10852 8878 10854
rect 8902 10852 8958 10854
rect 8982 10852 9038 10854
rect 9062 10852 9118 10854
rect 8850 10512 8906 10568
rect 8574 10376 8630 10432
rect 8822 9818 8878 9820
rect 8902 9818 8958 9820
rect 8982 9818 9038 9820
rect 9062 9818 9118 9820
rect 8822 9766 8848 9818
rect 8848 9766 8878 9818
rect 8902 9766 8912 9818
rect 8912 9766 8958 9818
rect 8982 9766 9028 9818
rect 9028 9766 9038 9818
rect 9062 9766 9092 9818
rect 9092 9766 9118 9818
rect 8822 9764 8878 9766
rect 8902 9764 8958 9766
rect 8982 9764 9038 9766
rect 9062 9764 9118 9766
rect 9494 10376 9550 10432
rect 10230 10684 10232 10704
rect 10232 10684 10284 10704
rect 10284 10684 10286 10704
rect 10230 10648 10286 10684
rect 8822 8730 8878 8732
rect 8902 8730 8958 8732
rect 8982 8730 9038 8732
rect 9062 8730 9118 8732
rect 8822 8678 8848 8730
rect 8848 8678 8878 8730
rect 8902 8678 8912 8730
rect 8912 8678 8958 8730
rect 8982 8678 9028 8730
rect 9028 8678 9038 8730
rect 9062 8678 9092 8730
rect 9092 8678 9118 8730
rect 8822 8676 8878 8678
rect 8902 8676 8958 8678
rect 8982 8676 9038 8678
rect 9062 8676 9118 8678
rect 8822 7642 8878 7644
rect 8902 7642 8958 7644
rect 8982 7642 9038 7644
rect 9062 7642 9118 7644
rect 8822 7590 8848 7642
rect 8848 7590 8878 7642
rect 8902 7590 8912 7642
rect 8912 7590 8958 7642
rect 8982 7590 9028 7642
rect 9028 7590 9038 7642
rect 9062 7590 9092 7642
rect 9092 7590 9118 7642
rect 8822 7588 8878 7590
rect 8902 7588 8958 7590
rect 8982 7588 9038 7590
rect 9062 7588 9118 7590
rect 8822 6554 8878 6556
rect 8902 6554 8958 6556
rect 8982 6554 9038 6556
rect 9062 6554 9118 6556
rect 8822 6502 8848 6554
rect 8848 6502 8878 6554
rect 8902 6502 8912 6554
rect 8912 6502 8958 6554
rect 8982 6502 9028 6554
rect 9028 6502 9038 6554
rect 9062 6502 9092 6554
rect 9092 6502 9118 6554
rect 8822 6500 8878 6502
rect 8902 6500 8958 6502
rect 8982 6500 9038 6502
rect 9062 6500 9118 6502
rect 14066 17434 14122 17436
rect 14146 17434 14202 17436
rect 14226 17434 14282 17436
rect 14306 17434 14362 17436
rect 14066 17382 14092 17434
rect 14092 17382 14122 17434
rect 14146 17382 14156 17434
rect 14156 17382 14202 17434
rect 14226 17382 14272 17434
rect 14272 17382 14282 17434
rect 14306 17382 14336 17434
rect 14336 17382 14362 17434
rect 14066 17380 14122 17382
rect 14146 17380 14202 17382
rect 14226 17380 14282 17382
rect 14306 17380 14362 17382
rect 11444 12538 11500 12540
rect 11524 12538 11580 12540
rect 11604 12538 11660 12540
rect 11684 12538 11740 12540
rect 11444 12486 11470 12538
rect 11470 12486 11500 12538
rect 11524 12486 11534 12538
rect 11534 12486 11580 12538
rect 11604 12486 11650 12538
rect 11650 12486 11660 12538
rect 11684 12486 11714 12538
rect 11714 12486 11740 12538
rect 11444 12484 11500 12486
rect 11524 12484 11580 12486
rect 11604 12484 11660 12486
rect 11684 12484 11740 12486
rect 11444 11450 11500 11452
rect 11524 11450 11580 11452
rect 11604 11450 11660 11452
rect 11684 11450 11740 11452
rect 11444 11398 11470 11450
rect 11470 11398 11500 11450
rect 11524 11398 11534 11450
rect 11534 11398 11580 11450
rect 11604 11398 11650 11450
rect 11650 11398 11660 11450
rect 11684 11398 11714 11450
rect 11714 11398 11740 11450
rect 11444 11396 11500 11398
rect 11524 11396 11580 11398
rect 11604 11396 11660 11398
rect 11684 11396 11740 11398
rect 10874 9460 10876 9480
rect 10876 9460 10928 9480
rect 10928 9460 10930 9480
rect 10874 9424 10930 9460
rect 10782 9036 10838 9072
rect 10782 9016 10784 9036
rect 10784 9016 10836 9036
rect 10836 9016 10838 9036
rect 11444 10362 11500 10364
rect 11524 10362 11580 10364
rect 11604 10362 11660 10364
rect 11684 10362 11740 10364
rect 11444 10310 11470 10362
rect 11470 10310 11500 10362
rect 11524 10310 11534 10362
rect 11534 10310 11580 10362
rect 11604 10310 11650 10362
rect 11650 10310 11660 10362
rect 11684 10310 11714 10362
rect 11714 10310 11740 10362
rect 11444 10308 11500 10310
rect 11524 10308 11580 10310
rect 11604 10308 11660 10310
rect 11684 10308 11740 10310
rect 11886 9460 11888 9480
rect 11888 9460 11940 9480
rect 11940 9460 11942 9480
rect 11886 9424 11942 9460
rect 11444 9274 11500 9276
rect 11524 9274 11580 9276
rect 11604 9274 11660 9276
rect 11684 9274 11740 9276
rect 11444 9222 11470 9274
rect 11470 9222 11500 9274
rect 11524 9222 11534 9274
rect 11534 9222 11580 9274
rect 11604 9222 11650 9274
rect 11650 9222 11660 9274
rect 11684 9222 11714 9274
rect 11714 9222 11740 9274
rect 11444 9220 11500 9222
rect 11524 9220 11580 9222
rect 11604 9220 11660 9222
rect 11684 9220 11740 9222
rect 11794 9016 11850 9072
rect 11444 8186 11500 8188
rect 11524 8186 11580 8188
rect 11604 8186 11660 8188
rect 11684 8186 11740 8188
rect 11444 8134 11470 8186
rect 11470 8134 11500 8186
rect 11524 8134 11534 8186
rect 11534 8134 11580 8186
rect 11604 8134 11650 8186
rect 11650 8134 11660 8186
rect 11684 8134 11714 8186
rect 11714 8134 11740 8186
rect 11444 8132 11500 8134
rect 11524 8132 11580 8134
rect 11604 8132 11660 8134
rect 11684 8132 11740 8134
rect 10966 7284 10968 7304
rect 10968 7284 11020 7304
rect 11020 7284 11022 7304
rect 8822 5466 8878 5468
rect 8902 5466 8958 5468
rect 8982 5466 9038 5468
rect 9062 5466 9118 5468
rect 8822 5414 8848 5466
rect 8848 5414 8878 5466
rect 8902 5414 8912 5466
rect 8912 5414 8958 5466
rect 8982 5414 9028 5466
rect 9028 5414 9038 5466
rect 9062 5414 9092 5466
rect 9092 5414 9118 5466
rect 8822 5412 8878 5414
rect 8902 5412 8958 5414
rect 8982 5412 9038 5414
rect 9062 5412 9118 5414
rect 8822 4378 8878 4380
rect 8902 4378 8958 4380
rect 8982 4378 9038 4380
rect 9062 4378 9118 4380
rect 8822 4326 8848 4378
rect 8848 4326 8878 4378
rect 8902 4326 8912 4378
rect 8912 4326 8958 4378
rect 8982 4326 9028 4378
rect 9028 4326 9038 4378
rect 9062 4326 9092 4378
rect 9092 4326 9118 4378
rect 8822 4324 8878 4326
rect 8902 4324 8958 4326
rect 8982 4324 9038 4326
rect 9062 4324 9118 4326
rect 8822 3290 8878 3292
rect 8902 3290 8958 3292
rect 8982 3290 9038 3292
rect 9062 3290 9118 3292
rect 8822 3238 8848 3290
rect 8848 3238 8878 3290
rect 8902 3238 8912 3290
rect 8912 3238 8958 3290
rect 8982 3238 9028 3290
rect 9028 3238 9038 3290
rect 9062 3238 9092 3290
rect 9092 3238 9118 3290
rect 8822 3236 8878 3238
rect 8902 3236 8958 3238
rect 8982 3236 9038 3238
rect 9062 3236 9118 3238
rect 10966 7248 11022 7284
rect 11444 7098 11500 7100
rect 11524 7098 11580 7100
rect 11604 7098 11660 7100
rect 11684 7098 11740 7100
rect 11444 7046 11470 7098
rect 11470 7046 11500 7098
rect 11524 7046 11534 7098
rect 11534 7046 11580 7098
rect 11604 7046 11650 7098
rect 11650 7046 11660 7098
rect 11684 7046 11714 7098
rect 11714 7046 11740 7098
rect 11444 7044 11500 7046
rect 11524 7044 11580 7046
rect 11604 7044 11660 7046
rect 11684 7044 11740 7046
rect 12714 12008 12770 12064
rect 14066 16346 14122 16348
rect 14146 16346 14202 16348
rect 14226 16346 14282 16348
rect 14306 16346 14362 16348
rect 14066 16294 14092 16346
rect 14092 16294 14122 16346
rect 14146 16294 14156 16346
rect 14156 16294 14202 16346
rect 14226 16294 14272 16346
rect 14272 16294 14282 16346
rect 14306 16294 14336 16346
rect 14336 16294 14362 16346
rect 14066 16292 14122 16294
rect 14146 16292 14202 16294
rect 14226 16292 14282 16294
rect 14306 16292 14362 16294
rect 12622 10648 12678 10704
rect 14066 15258 14122 15260
rect 14146 15258 14202 15260
rect 14226 15258 14282 15260
rect 14306 15258 14362 15260
rect 14066 15206 14092 15258
rect 14092 15206 14122 15258
rect 14146 15206 14156 15258
rect 14156 15206 14202 15258
rect 14226 15206 14272 15258
rect 14272 15206 14282 15258
rect 14306 15206 14336 15258
rect 14336 15206 14362 15258
rect 14066 15204 14122 15206
rect 14146 15204 14202 15206
rect 14226 15204 14282 15206
rect 14306 15204 14362 15206
rect 14066 14170 14122 14172
rect 14146 14170 14202 14172
rect 14226 14170 14282 14172
rect 14306 14170 14362 14172
rect 14066 14118 14092 14170
rect 14092 14118 14122 14170
rect 14146 14118 14156 14170
rect 14156 14118 14202 14170
rect 14226 14118 14272 14170
rect 14272 14118 14282 14170
rect 14306 14118 14336 14170
rect 14336 14118 14362 14170
rect 14066 14116 14122 14118
rect 14146 14116 14202 14118
rect 14226 14116 14282 14118
rect 14306 14116 14362 14118
rect 14066 13082 14122 13084
rect 14146 13082 14202 13084
rect 14226 13082 14282 13084
rect 14306 13082 14362 13084
rect 14066 13030 14092 13082
rect 14092 13030 14122 13082
rect 14146 13030 14156 13082
rect 14156 13030 14202 13082
rect 14226 13030 14272 13082
rect 14272 13030 14282 13082
rect 14306 13030 14336 13082
rect 14336 13030 14362 13082
rect 14066 13028 14122 13030
rect 14146 13028 14202 13030
rect 14226 13028 14282 13030
rect 14306 13028 14362 13030
rect 14066 11994 14122 11996
rect 14146 11994 14202 11996
rect 14226 11994 14282 11996
rect 14306 11994 14362 11996
rect 14066 11942 14092 11994
rect 14092 11942 14122 11994
rect 14146 11942 14156 11994
rect 14156 11942 14202 11994
rect 14226 11942 14272 11994
rect 14272 11942 14282 11994
rect 14306 11942 14336 11994
rect 14336 11942 14362 11994
rect 14066 11940 14122 11942
rect 14146 11940 14202 11942
rect 14226 11940 14282 11942
rect 14306 11940 14362 11942
rect 12622 9968 12678 10024
rect 14066 10906 14122 10908
rect 14146 10906 14202 10908
rect 14226 10906 14282 10908
rect 14306 10906 14362 10908
rect 14066 10854 14092 10906
rect 14092 10854 14122 10906
rect 14146 10854 14156 10906
rect 14156 10854 14202 10906
rect 14226 10854 14272 10906
rect 14272 10854 14282 10906
rect 14306 10854 14336 10906
rect 14336 10854 14362 10906
rect 14066 10852 14122 10854
rect 14146 10852 14202 10854
rect 14226 10852 14282 10854
rect 14306 10852 14362 10854
rect 14066 9818 14122 9820
rect 14146 9818 14202 9820
rect 14226 9818 14282 9820
rect 14306 9818 14362 9820
rect 14066 9766 14092 9818
rect 14092 9766 14122 9818
rect 14146 9766 14156 9818
rect 14156 9766 14202 9818
rect 14226 9766 14272 9818
rect 14272 9766 14282 9818
rect 14306 9766 14336 9818
rect 14336 9766 14362 9818
rect 14066 9764 14122 9766
rect 14146 9764 14202 9766
rect 14226 9764 14282 9766
rect 14306 9764 14362 9766
rect 11444 6010 11500 6012
rect 11524 6010 11580 6012
rect 11604 6010 11660 6012
rect 11684 6010 11740 6012
rect 11444 5958 11470 6010
rect 11470 5958 11500 6010
rect 11524 5958 11534 6010
rect 11534 5958 11580 6010
rect 11604 5958 11650 6010
rect 11650 5958 11660 6010
rect 11684 5958 11714 6010
rect 11714 5958 11740 6010
rect 11444 5956 11500 5958
rect 11524 5956 11580 5958
rect 11604 5956 11660 5958
rect 11684 5956 11740 5958
rect 12898 7248 12954 7304
rect 11444 4922 11500 4924
rect 11524 4922 11580 4924
rect 11604 4922 11660 4924
rect 11684 4922 11740 4924
rect 11444 4870 11470 4922
rect 11470 4870 11500 4922
rect 11524 4870 11534 4922
rect 11534 4870 11580 4922
rect 11604 4870 11650 4922
rect 11650 4870 11660 4922
rect 11684 4870 11714 4922
rect 11714 4870 11740 4922
rect 11444 4868 11500 4870
rect 11524 4868 11580 4870
rect 11604 4868 11660 4870
rect 11684 4868 11740 4870
rect 11444 3834 11500 3836
rect 11524 3834 11580 3836
rect 11604 3834 11660 3836
rect 11684 3834 11740 3836
rect 11444 3782 11470 3834
rect 11470 3782 11500 3834
rect 11524 3782 11534 3834
rect 11534 3782 11580 3834
rect 11604 3782 11650 3834
rect 11650 3782 11660 3834
rect 11684 3782 11714 3834
rect 11714 3782 11740 3834
rect 11444 3780 11500 3782
rect 11524 3780 11580 3782
rect 11604 3780 11660 3782
rect 11684 3780 11740 3782
rect 14066 8730 14122 8732
rect 14146 8730 14202 8732
rect 14226 8730 14282 8732
rect 14306 8730 14362 8732
rect 14066 8678 14092 8730
rect 14092 8678 14122 8730
rect 14146 8678 14156 8730
rect 14156 8678 14202 8730
rect 14226 8678 14272 8730
rect 14272 8678 14282 8730
rect 14306 8678 14336 8730
rect 14336 8678 14362 8730
rect 14066 8676 14122 8678
rect 14146 8676 14202 8678
rect 14226 8676 14282 8678
rect 14306 8676 14362 8678
rect 14066 7642 14122 7644
rect 14146 7642 14202 7644
rect 14226 7642 14282 7644
rect 14306 7642 14362 7644
rect 14066 7590 14092 7642
rect 14092 7590 14122 7642
rect 14146 7590 14156 7642
rect 14156 7590 14202 7642
rect 14226 7590 14272 7642
rect 14272 7590 14282 7642
rect 14306 7590 14336 7642
rect 14336 7590 14362 7642
rect 14066 7588 14122 7590
rect 14146 7588 14202 7590
rect 14226 7588 14282 7590
rect 14306 7588 14362 7590
rect 14066 6554 14122 6556
rect 14146 6554 14202 6556
rect 14226 6554 14282 6556
rect 14306 6554 14362 6556
rect 14066 6502 14092 6554
rect 14092 6502 14122 6554
rect 14146 6502 14156 6554
rect 14156 6502 14202 6554
rect 14226 6502 14272 6554
rect 14272 6502 14282 6554
rect 14306 6502 14336 6554
rect 14336 6502 14362 6554
rect 14066 6500 14122 6502
rect 14146 6500 14202 6502
rect 14226 6500 14282 6502
rect 14306 6500 14362 6502
rect 14066 5466 14122 5468
rect 14146 5466 14202 5468
rect 14226 5466 14282 5468
rect 14306 5466 14362 5468
rect 14066 5414 14092 5466
rect 14092 5414 14122 5466
rect 14146 5414 14156 5466
rect 14156 5414 14202 5466
rect 14226 5414 14272 5466
rect 14272 5414 14282 5466
rect 14306 5414 14336 5466
rect 14336 5414 14362 5466
rect 14066 5412 14122 5414
rect 14146 5412 14202 5414
rect 14226 5412 14282 5414
rect 14306 5412 14362 5414
rect 16486 15680 16542 15736
rect 15750 11636 15752 11656
rect 15752 11636 15804 11656
rect 15804 11636 15806 11656
rect 15750 11600 15806 11636
rect 15566 9968 15622 10024
rect 14066 4378 14122 4380
rect 14146 4378 14202 4380
rect 14226 4378 14282 4380
rect 14306 4378 14362 4380
rect 14066 4326 14092 4378
rect 14092 4326 14122 4378
rect 14146 4326 14156 4378
rect 14156 4326 14202 4378
rect 14226 4326 14272 4378
rect 14272 4326 14282 4378
rect 14306 4326 14336 4378
rect 14336 4326 14362 4378
rect 14066 4324 14122 4326
rect 14146 4324 14202 4326
rect 14226 4324 14282 4326
rect 14306 4324 14362 4326
rect 14066 3290 14122 3292
rect 14146 3290 14202 3292
rect 14226 3290 14282 3292
rect 14306 3290 14362 3292
rect 14066 3238 14092 3290
rect 14092 3238 14122 3290
rect 14146 3238 14156 3290
rect 14156 3238 14202 3290
rect 14226 3238 14272 3290
rect 14272 3238 14282 3290
rect 14306 3238 14336 3290
rect 14336 3238 14362 3290
rect 14066 3236 14122 3238
rect 14146 3236 14202 3238
rect 14226 3236 14282 3238
rect 14306 3236 14362 3238
rect 8758 2932 8760 2952
rect 8760 2932 8812 2952
rect 8812 2932 8814 2952
rect 8758 2896 8814 2932
rect 8822 2202 8878 2204
rect 8902 2202 8958 2204
rect 8982 2202 9038 2204
rect 9062 2202 9118 2204
rect 8822 2150 8848 2202
rect 8848 2150 8878 2202
rect 8902 2150 8912 2202
rect 8912 2150 8958 2202
rect 8982 2150 9028 2202
rect 9028 2150 9038 2202
rect 9062 2150 9092 2202
rect 9092 2150 9118 2202
rect 8822 2148 8878 2150
rect 8902 2148 8958 2150
rect 8982 2148 9038 2150
rect 9062 2148 9118 2150
rect 11444 2746 11500 2748
rect 11524 2746 11580 2748
rect 11604 2746 11660 2748
rect 11684 2746 11740 2748
rect 11444 2694 11470 2746
rect 11470 2694 11500 2746
rect 11524 2694 11534 2746
rect 11534 2694 11580 2746
rect 11604 2694 11650 2746
rect 11650 2694 11660 2746
rect 11684 2694 11714 2746
rect 11714 2694 11740 2746
rect 11444 2692 11500 2694
rect 11524 2692 11580 2694
rect 11604 2692 11660 2694
rect 11684 2692 11740 2694
rect 14066 2202 14122 2204
rect 14146 2202 14202 2204
rect 14226 2202 14282 2204
rect 14306 2202 14362 2204
rect 14066 2150 14092 2202
rect 14092 2150 14122 2202
rect 14146 2150 14156 2202
rect 14156 2150 14202 2202
rect 14226 2150 14272 2202
rect 14272 2150 14282 2202
rect 14306 2150 14336 2202
rect 14336 2150 14362 2202
rect 14066 2148 14122 2150
rect 14146 2148 14202 2150
rect 14226 2148 14282 2150
rect 14306 2148 14362 2150
rect 16486 13640 16542 13696
rect 16486 10920 16542 10976
rect 16302 9968 16358 10024
rect 16486 8200 16542 8256
rect 16486 6196 16488 6216
rect 16488 6196 16540 6216
rect 16540 6196 16542 6216
rect 16486 6160 16542 6196
rect 16486 3440 16542 3496
rect 16486 1400 16542 1456
<< metal3 >>
rect 16113 18458 16179 18461
rect 17227 18458 18027 18488
rect 16113 18456 18027 18458
rect 16113 18400 16118 18456
rect 16174 18400 18027 18456
rect 16113 18398 18027 18400
rect 16113 18395 16179 18398
rect 17227 18368 18027 18398
rect 6188 17984 6508 17985
rect 6188 17920 6196 17984
rect 6260 17920 6276 17984
rect 6340 17920 6356 17984
rect 6420 17920 6436 17984
rect 6500 17920 6508 17984
rect 6188 17919 6508 17920
rect 11432 17984 11752 17985
rect 11432 17920 11440 17984
rect 11504 17920 11520 17984
rect 11584 17920 11600 17984
rect 11664 17920 11680 17984
rect 11744 17920 11752 17984
rect 11432 17919 11752 17920
rect 3566 17440 3886 17441
rect 3566 17376 3574 17440
rect 3638 17376 3654 17440
rect 3718 17376 3734 17440
rect 3798 17376 3814 17440
rect 3878 17376 3886 17440
rect 3566 17375 3886 17376
rect 8810 17440 9130 17441
rect 8810 17376 8818 17440
rect 8882 17376 8898 17440
rect 8962 17376 8978 17440
rect 9042 17376 9058 17440
rect 9122 17376 9130 17440
rect 8810 17375 9130 17376
rect 14054 17440 14374 17441
rect 14054 17376 14062 17440
rect 14126 17376 14142 17440
rect 14206 17376 14222 17440
rect 14286 17376 14302 17440
rect 14366 17376 14374 17440
rect 14054 17375 14374 17376
rect 0 17098 800 17128
rect 1393 17098 1459 17101
rect 0 17096 1459 17098
rect 0 17040 1398 17096
rect 1454 17040 1459 17096
rect 0 17038 1459 17040
rect 0 17008 800 17038
rect 1393 17035 1459 17038
rect 6188 16896 6508 16897
rect 6188 16832 6196 16896
rect 6260 16832 6276 16896
rect 6340 16832 6356 16896
rect 6420 16832 6436 16896
rect 6500 16832 6508 16896
rect 6188 16831 6508 16832
rect 11432 16896 11752 16897
rect 11432 16832 11440 16896
rect 11504 16832 11520 16896
rect 11584 16832 11600 16896
rect 11664 16832 11680 16896
rect 11744 16832 11752 16896
rect 11432 16831 11752 16832
rect 3566 16352 3886 16353
rect 3566 16288 3574 16352
rect 3638 16288 3654 16352
rect 3718 16288 3734 16352
rect 3798 16288 3814 16352
rect 3878 16288 3886 16352
rect 3566 16287 3886 16288
rect 8810 16352 9130 16353
rect 8810 16288 8818 16352
rect 8882 16288 8898 16352
rect 8962 16288 8978 16352
rect 9042 16288 9058 16352
rect 9122 16288 9130 16352
rect 8810 16287 9130 16288
rect 14054 16352 14374 16353
rect 14054 16288 14062 16352
rect 14126 16288 14142 16352
rect 14206 16288 14222 16352
rect 14286 16288 14302 16352
rect 14366 16288 14374 16352
rect 14054 16287 14374 16288
rect 6188 15808 6508 15809
rect 6188 15744 6196 15808
rect 6260 15744 6276 15808
rect 6340 15744 6356 15808
rect 6420 15744 6436 15808
rect 6500 15744 6508 15808
rect 6188 15743 6508 15744
rect 11432 15808 11752 15809
rect 11432 15744 11440 15808
rect 11504 15744 11520 15808
rect 11584 15744 11600 15808
rect 11664 15744 11680 15808
rect 11744 15744 11752 15808
rect 11432 15743 11752 15744
rect 16481 15738 16547 15741
rect 17227 15738 18027 15768
rect 16481 15736 18027 15738
rect 16481 15680 16486 15736
rect 16542 15680 18027 15736
rect 16481 15678 18027 15680
rect 16481 15675 16547 15678
rect 17227 15648 18027 15678
rect 3566 15264 3886 15265
rect 3566 15200 3574 15264
rect 3638 15200 3654 15264
rect 3718 15200 3734 15264
rect 3798 15200 3814 15264
rect 3878 15200 3886 15264
rect 3566 15199 3886 15200
rect 8810 15264 9130 15265
rect 8810 15200 8818 15264
rect 8882 15200 8898 15264
rect 8962 15200 8978 15264
rect 9042 15200 9058 15264
rect 9122 15200 9130 15264
rect 8810 15199 9130 15200
rect 14054 15264 14374 15265
rect 14054 15200 14062 15264
rect 14126 15200 14142 15264
rect 14206 15200 14222 15264
rect 14286 15200 14302 15264
rect 14366 15200 14374 15264
rect 14054 15199 14374 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 6188 14720 6508 14721
rect 6188 14656 6196 14720
rect 6260 14656 6276 14720
rect 6340 14656 6356 14720
rect 6420 14656 6436 14720
rect 6500 14656 6508 14720
rect 6188 14655 6508 14656
rect 11432 14720 11752 14721
rect 11432 14656 11440 14720
rect 11504 14656 11520 14720
rect 11584 14656 11600 14720
rect 11664 14656 11680 14720
rect 11744 14656 11752 14720
rect 11432 14655 11752 14656
rect 6177 14514 6243 14517
rect 6913 14514 6979 14517
rect 6177 14512 6979 14514
rect 6177 14456 6182 14512
rect 6238 14456 6918 14512
rect 6974 14456 6979 14512
rect 6177 14454 6979 14456
rect 6177 14451 6243 14454
rect 6913 14451 6979 14454
rect 5993 14378 6059 14381
rect 6637 14378 6703 14381
rect 5993 14376 6703 14378
rect 5993 14320 5998 14376
rect 6054 14320 6642 14376
rect 6698 14320 6703 14376
rect 5993 14318 6703 14320
rect 5993 14315 6059 14318
rect 6637 14315 6703 14318
rect 3566 14176 3886 14177
rect 3566 14112 3574 14176
rect 3638 14112 3654 14176
rect 3718 14112 3734 14176
rect 3798 14112 3814 14176
rect 3878 14112 3886 14176
rect 3566 14111 3886 14112
rect 8810 14176 9130 14177
rect 8810 14112 8818 14176
rect 8882 14112 8898 14176
rect 8962 14112 8978 14176
rect 9042 14112 9058 14176
rect 9122 14112 9130 14176
rect 8810 14111 9130 14112
rect 14054 14176 14374 14177
rect 14054 14112 14062 14176
rect 14126 14112 14142 14176
rect 14206 14112 14222 14176
rect 14286 14112 14302 14176
rect 14366 14112 14374 14176
rect 14054 14111 14374 14112
rect 16481 13698 16547 13701
rect 17227 13698 18027 13728
rect 16481 13696 18027 13698
rect 16481 13640 16486 13696
rect 16542 13640 18027 13696
rect 16481 13638 18027 13640
rect 16481 13635 16547 13638
rect 6188 13632 6508 13633
rect 6188 13568 6196 13632
rect 6260 13568 6276 13632
rect 6340 13568 6356 13632
rect 6420 13568 6436 13632
rect 6500 13568 6508 13632
rect 6188 13567 6508 13568
rect 11432 13632 11752 13633
rect 11432 13568 11440 13632
rect 11504 13568 11520 13632
rect 11584 13568 11600 13632
rect 11664 13568 11680 13632
rect 11744 13568 11752 13632
rect 17227 13608 18027 13638
rect 11432 13567 11752 13568
rect 3877 13426 3943 13429
rect 5165 13426 5231 13429
rect 3877 13424 5231 13426
rect 3877 13368 3882 13424
rect 3938 13368 5170 13424
rect 5226 13368 5231 13424
rect 3877 13366 5231 13368
rect 3877 13363 3943 13366
rect 5165 13363 5231 13366
rect 3566 13088 3886 13089
rect 3566 13024 3574 13088
rect 3638 13024 3654 13088
rect 3718 13024 3734 13088
rect 3798 13024 3814 13088
rect 3878 13024 3886 13088
rect 3566 13023 3886 13024
rect 8810 13088 9130 13089
rect 8810 13024 8818 13088
rect 8882 13024 8898 13088
rect 8962 13024 8978 13088
rect 9042 13024 9058 13088
rect 9122 13024 9130 13088
rect 8810 13023 9130 13024
rect 14054 13088 14374 13089
rect 14054 13024 14062 13088
rect 14126 13024 14142 13088
rect 14206 13024 14222 13088
rect 14286 13024 14302 13088
rect 14366 13024 14374 13088
rect 14054 13023 14374 13024
rect 6188 12544 6508 12545
rect 6188 12480 6196 12544
rect 6260 12480 6276 12544
rect 6340 12480 6356 12544
rect 6420 12480 6436 12544
rect 6500 12480 6508 12544
rect 6188 12479 6508 12480
rect 11432 12544 11752 12545
rect 11432 12480 11440 12544
rect 11504 12480 11520 12544
rect 11584 12480 11600 12544
rect 11664 12480 11680 12544
rect 11744 12480 11752 12544
rect 11432 12479 11752 12480
rect 0 12338 800 12368
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 1577 12202 1643 12205
rect 8385 12202 8451 12205
rect 1577 12200 8451 12202
rect 1577 12144 1582 12200
rect 1638 12144 8390 12200
rect 8446 12144 8451 12200
rect 1577 12142 8451 12144
rect 1577 12139 1643 12142
rect 8385 12139 8451 12142
rect 9397 12066 9463 12069
rect 12709 12066 12775 12069
rect 9397 12064 12775 12066
rect 9397 12008 9402 12064
rect 9458 12008 12714 12064
rect 12770 12008 12775 12064
rect 9397 12006 12775 12008
rect 9397 12003 9463 12006
rect 12709 12003 12775 12006
rect 3566 12000 3886 12001
rect 3566 11936 3574 12000
rect 3638 11936 3654 12000
rect 3718 11936 3734 12000
rect 3798 11936 3814 12000
rect 3878 11936 3886 12000
rect 3566 11935 3886 11936
rect 8810 12000 9130 12001
rect 8810 11936 8818 12000
rect 8882 11936 8898 12000
rect 8962 11936 8978 12000
rect 9042 11936 9058 12000
rect 9122 11936 9130 12000
rect 8810 11935 9130 11936
rect 14054 12000 14374 12001
rect 14054 11936 14062 12000
rect 14126 11936 14142 12000
rect 14206 11936 14222 12000
rect 14286 11936 14302 12000
rect 14366 11936 14374 12000
rect 14054 11935 14374 11936
rect 15745 11658 15811 11661
rect 11286 11656 15811 11658
rect 11286 11600 15750 11656
rect 15806 11600 15811 11656
rect 11286 11598 15811 11600
rect 8845 11522 8911 11525
rect 11286 11522 11346 11598
rect 15745 11595 15811 11598
rect 8845 11520 11346 11522
rect 8845 11464 8850 11520
rect 8906 11464 11346 11520
rect 8845 11462 11346 11464
rect 8845 11459 8911 11462
rect 6188 11456 6508 11457
rect 6188 11392 6196 11456
rect 6260 11392 6276 11456
rect 6340 11392 6356 11456
rect 6420 11392 6436 11456
rect 6500 11392 6508 11456
rect 6188 11391 6508 11392
rect 11432 11456 11752 11457
rect 11432 11392 11440 11456
rect 11504 11392 11520 11456
rect 11584 11392 11600 11456
rect 11664 11392 11680 11456
rect 11744 11392 11752 11456
rect 11432 11391 11752 11392
rect 16481 10978 16547 10981
rect 17227 10978 18027 11008
rect 16481 10976 18027 10978
rect 16481 10920 16486 10976
rect 16542 10920 18027 10976
rect 16481 10918 18027 10920
rect 16481 10915 16547 10918
rect 3566 10912 3886 10913
rect 3566 10848 3574 10912
rect 3638 10848 3654 10912
rect 3718 10848 3734 10912
rect 3798 10848 3814 10912
rect 3878 10848 3886 10912
rect 3566 10847 3886 10848
rect 8810 10912 9130 10913
rect 8810 10848 8818 10912
rect 8882 10848 8898 10912
rect 8962 10848 8978 10912
rect 9042 10848 9058 10912
rect 9122 10848 9130 10912
rect 8810 10847 9130 10848
rect 14054 10912 14374 10913
rect 14054 10848 14062 10912
rect 14126 10848 14142 10912
rect 14206 10848 14222 10912
rect 14286 10848 14302 10912
rect 14366 10848 14374 10912
rect 17227 10888 18027 10918
rect 14054 10847 14374 10848
rect 10225 10706 10291 10709
rect 12617 10706 12683 10709
rect 10225 10704 12683 10706
rect 10225 10648 10230 10704
rect 10286 10648 12622 10704
rect 12678 10648 12683 10704
rect 10225 10646 12683 10648
rect 10225 10643 10291 10646
rect 12617 10643 12683 10646
rect 7189 10570 7255 10573
rect 8845 10570 8911 10573
rect 7189 10568 8911 10570
rect 7189 10512 7194 10568
rect 7250 10512 8850 10568
rect 8906 10512 8911 10568
rect 7189 10510 8911 10512
rect 7189 10507 7255 10510
rect 8845 10507 8911 10510
rect 8569 10434 8635 10437
rect 9489 10434 9555 10437
rect 8569 10432 9555 10434
rect 8569 10376 8574 10432
rect 8630 10376 9494 10432
rect 9550 10376 9555 10432
rect 8569 10374 9555 10376
rect 8569 10371 8635 10374
rect 9489 10371 9555 10374
rect 6188 10368 6508 10369
rect 0 10298 800 10328
rect 6188 10304 6196 10368
rect 6260 10304 6276 10368
rect 6340 10304 6356 10368
rect 6420 10304 6436 10368
rect 6500 10304 6508 10368
rect 6188 10303 6508 10304
rect 11432 10368 11752 10369
rect 11432 10304 11440 10368
rect 11504 10304 11520 10368
rect 11584 10304 11600 10368
rect 11664 10304 11680 10368
rect 11744 10304 11752 10368
rect 11432 10303 11752 10304
rect 1393 10298 1459 10301
rect 0 10296 1459 10298
rect 0 10240 1398 10296
rect 1454 10240 1459 10296
rect 0 10238 1459 10240
rect 0 10208 800 10238
rect 1393 10235 1459 10238
rect 12617 10026 12683 10029
rect 15561 10026 15627 10029
rect 16297 10026 16363 10029
rect 12617 10024 16363 10026
rect 12617 9968 12622 10024
rect 12678 9968 15566 10024
rect 15622 9968 16302 10024
rect 16358 9968 16363 10024
rect 12617 9966 16363 9968
rect 12617 9963 12683 9966
rect 15561 9963 15627 9966
rect 16297 9963 16363 9966
rect 3566 9824 3886 9825
rect 3566 9760 3574 9824
rect 3638 9760 3654 9824
rect 3718 9760 3734 9824
rect 3798 9760 3814 9824
rect 3878 9760 3886 9824
rect 3566 9759 3886 9760
rect 8810 9824 9130 9825
rect 8810 9760 8818 9824
rect 8882 9760 8898 9824
rect 8962 9760 8978 9824
rect 9042 9760 9058 9824
rect 9122 9760 9130 9824
rect 8810 9759 9130 9760
rect 14054 9824 14374 9825
rect 14054 9760 14062 9824
rect 14126 9760 14142 9824
rect 14206 9760 14222 9824
rect 14286 9760 14302 9824
rect 14366 9760 14374 9824
rect 14054 9759 14374 9760
rect 10869 9482 10935 9485
rect 11881 9482 11947 9485
rect 10869 9480 11947 9482
rect 10869 9424 10874 9480
rect 10930 9424 11886 9480
rect 11942 9424 11947 9480
rect 10869 9422 11947 9424
rect 10869 9419 10935 9422
rect 11881 9419 11947 9422
rect 6188 9280 6508 9281
rect 6188 9216 6196 9280
rect 6260 9216 6276 9280
rect 6340 9216 6356 9280
rect 6420 9216 6436 9280
rect 6500 9216 6508 9280
rect 6188 9215 6508 9216
rect 11432 9280 11752 9281
rect 11432 9216 11440 9280
rect 11504 9216 11520 9280
rect 11584 9216 11600 9280
rect 11664 9216 11680 9280
rect 11744 9216 11752 9280
rect 11432 9215 11752 9216
rect 10777 9074 10843 9077
rect 11789 9074 11855 9077
rect 10777 9072 11855 9074
rect 10777 9016 10782 9072
rect 10838 9016 11794 9072
rect 11850 9016 11855 9072
rect 10777 9014 11855 9016
rect 10777 9011 10843 9014
rect 11789 9011 11855 9014
rect 3566 8736 3886 8737
rect 3566 8672 3574 8736
rect 3638 8672 3654 8736
rect 3718 8672 3734 8736
rect 3798 8672 3814 8736
rect 3878 8672 3886 8736
rect 3566 8671 3886 8672
rect 8810 8736 9130 8737
rect 8810 8672 8818 8736
rect 8882 8672 8898 8736
rect 8962 8672 8978 8736
rect 9042 8672 9058 8736
rect 9122 8672 9130 8736
rect 8810 8671 9130 8672
rect 14054 8736 14374 8737
rect 14054 8672 14062 8736
rect 14126 8672 14142 8736
rect 14206 8672 14222 8736
rect 14286 8672 14302 8736
rect 14366 8672 14374 8736
rect 14054 8671 14374 8672
rect 16481 8258 16547 8261
rect 17227 8258 18027 8288
rect 16481 8256 18027 8258
rect 16481 8200 16486 8256
rect 16542 8200 18027 8256
rect 16481 8198 18027 8200
rect 16481 8195 16547 8198
rect 6188 8192 6508 8193
rect 6188 8128 6196 8192
rect 6260 8128 6276 8192
rect 6340 8128 6356 8192
rect 6420 8128 6436 8192
rect 6500 8128 6508 8192
rect 6188 8127 6508 8128
rect 11432 8192 11752 8193
rect 11432 8128 11440 8192
rect 11504 8128 11520 8192
rect 11584 8128 11600 8192
rect 11664 8128 11680 8192
rect 11744 8128 11752 8192
rect 17227 8168 18027 8198
rect 11432 8127 11752 8128
rect 3566 7648 3886 7649
rect 0 7578 800 7608
rect 3566 7584 3574 7648
rect 3638 7584 3654 7648
rect 3718 7584 3734 7648
rect 3798 7584 3814 7648
rect 3878 7584 3886 7648
rect 3566 7583 3886 7584
rect 8810 7648 9130 7649
rect 8810 7584 8818 7648
rect 8882 7584 8898 7648
rect 8962 7584 8978 7648
rect 9042 7584 9058 7648
rect 9122 7584 9130 7648
rect 8810 7583 9130 7584
rect 14054 7648 14374 7649
rect 14054 7584 14062 7648
rect 14126 7584 14142 7648
rect 14206 7584 14222 7648
rect 14286 7584 14302 7648
rect 14366 7584 14374 7648
rect 14054 7583 14374 7584
rect 1393 7578 1459 7581
rect 0 7576 1459 7578
rect 0 7520 1398 7576
rect 1454 7520 1459 7576
rect 0 7518 1459 7520
rect 0 7488 800 7518
rect 1393 7515 1459 7518
rect 10961 7306 11027 7309
rect 12893 7306 12959 7309
rect 10961 7304 12959 7306
rect 10961 7248 10966 7304
rect 11022 7248 12898 7304
rect 12954 7248 12959 7304
rect 10961 7246 12959 7248
rect 10961 7243 11027 7246
rect 12893 7243 12959 7246
rect 6188 7104 6508 7105
rect 6188 7040 6196 7104
rect 6260 7040 6276 7104
rect 6340 7040 6356 7104
rect 6420 7040 6436 7104
rect 6500 7040 6508 7104
rect 6188 7039 6508 7040
rect 11432 7104 11752 7105
rect 11432 7040 11440 7104
rect 11504 7040 11520 7104
rect 11584 7040 11600 7104
rect 11664 7040 11680 7104
rect 11744 7040 11752 7104
rect 11432 7039 11752 7040
rect 3566 6560 3886 6561
rect 3566 6496 3574 6560
rect 3638 6496 3654 6560
rect 3718 6496 3734 6560
rect 3798 6496 3814 6560
rect 3878 6496 3886 6560
rect 3566 6495 3886 6496
rect 8810 6560 9130 6561
rect 8810 6496 8818 6560
rect 8882 6496 8898 6560
rect 8962 6496 8978 6560
rect 9042 6496 9058 6560
rect 9122 6496 9130 6560
rect 8810 6495 9130 6496
rect 14054 6560 14374 6561
rect 14054 6496 14062 6560
rect 14126 6496 14142 6560
rect 14206 6496 14222 6560
rect 14286 6496 14302 6560
rect 14366 6496 14374 6560
rect 14054 6495 14374 6496
rect 16481 6218 16547 6221
rect 17227 6218 18027 6248
rect 16481 6216 18027 6218
rect 16481 6160 16486 6216
rect 16542 6160 18027 6216
rect 16481 6158 18027 6160
rect 16481 6155 16547 6158
rect 17227 6128 18027 6158
rect 6188 6016 6508 6017
rect 6188 5952 6196 6016
rect 6260 5952 6276 6016
rect 6340 5952 6356 6016
rect 6420 5952 6436 6016
rect 6500 5952 6508 6016
rect 6188 5951 6508 5952
rect 11432 6016 11752 6017
rect 11432 5952 11440 6016
rect 11504 5952 11520 6016
rect 11584 5952 11600 6016
rect 11664 5952 11680 6016
rect 11744 5952 11752 6016
rect 11432 5951 11752 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 3566 5472 3886 5473
rect 3566 5408 3574 5472
rect 3638 5408 3654 5472
rect 3718 5408 3734 5472
rect 3798 5408 3814 5472
rect 3878 5408 3886 5472
rect 3566 5407 3886 5408
rect 8810 5472 9130 5473
rect 8810 5408 8818 5472
rect 8882 5408 8898 5472
rect 8962 5408 8978 5472
rect 9042 5408 9058 5472
rect 9122 5408 9130 5472
rect 8810 5407 9130 5408
rect 14054 5472 14374 5473
rect 14054 5408 14062 5472
rect 14126 5408 14142 5472
rect 14206 5408 14222 5472
rect 14286 5408 14302 5472
rect 14366 5408 14374 5472
rect 14054 5407 14374 5408
rect 6188 4928 6508 4929
rect 6188 4864 6196 4928
rect 6260 4864 6276 4928
rect 6340 4864 6356 4928
rect 6420 4864 6436 4928
rect 6500 4864 6508 4928
rect 6188 4863 6508 4864
rect 11432 4928 11752 4929
rect 11432 4864 11440 4928
rect 11504 4864 11520 4928
rect 11584 4864 11600 4928
rect 11664 4864 11680 4928
rect 11744 4864 11752 4928
rect 11432 4863 11752 4864
rect 3566 4384 3886 4385
rect 3566 4320 3574 4384
rect 3638 4320 3654 4384
rect 3718 4320 3734 4384
rect 3798 4320 3814 4384
rect 3878 4320 3886 4384
rect 3566 4319 3886 4320
rect 8810 4384 9130 4385
rect 8810 4320 8818 4384
rect 8882 4320 8898 4384
rect 8962 4320 8978 4384
rect 9042 4320 9058 4384
rect 9122 4320 9130 4384
rect 8810 4319 9130 4320
rect 14054 4384 14374 4385
rect 14054 4320 14062 4384
rect 14126 4320 14142 4384
rect 14206 4320 14222 4384
rect 14286 4320 14302 4384
rect 14366 4320 14374 4384
rect 14054 4319 14374 4320
rect 6188 3840 6508 3841
rect 6188 3776 6196 3840
rect 6260 3776 6276 3840
rect 6340 3776 6356 3840
rect 6420 3776 6436 3840
rect 6500 3776 6508 3840
rect 6188 3775 6508 3776
rect 11432 3840 11752 3841
rect 11432 3776 11440 3840
rect 11504 3776 11520 3840
rect 11584 3776 11600 3840
rect 11664 3776 11680 3840
rect 11744 3776 11752 3840
rect 11432 3775 11752 3776
rect 16481 3498 16547 3501
rect 17227 3498 18027 3528
rect 16481 3496 18027 3498
rect 16481 3440 16486 3496
rect 16542 3440 18027 3496
rect 16481 3438 18027 3440
rect 16481 3435 16547 3438
rect 17227 3408 18027 3438
rect 3566 3296 3886 3297
rect 3566 3232 3574 3296
rect 3638 3232 3654 3296
rect 3718 3232 3734 3296
rect 3798 3232 3814 3296
rect 3878 3232 3886 3296
rect 3566 3231 3886 3232
rect 8810 3296 9130 3297
rect 8810 3232 8818 3296
rect 8882 3232 8898 3296
rect 8962 3232 8978 3296
rect 9042 3232 9058 3296
rect 9122 3232 9130 3296
rect 8810 3231 9130 3232
rect 14054 3296 14374 3297
rect 14054 3232 14062 3296
rect 14126 3232 14142 3296
rect 14206 3232 14222 3296
rect 14286 3232 14302 3296
rect 14366 3232 14374 3296
rect 14054 3231 14374 3232
rect 7005 2954 7071 2957
rect 8753 2954 8819 2957
rect 7005 2952 8819 2954
rect 7005 2896 7010 2952
rect 7066 2896 8758 2952
rect 8814 2896 8819 2952
rect 7005 2894 8819 2896
rect 7005 2891 7071 2894
rect 8753 2891 8819 2894
rect 0 2818 800 2848
rect 1393 2818 1459 2821
rect 0 2816 1459 2818
rect 0 2760 1398 2816
rect 1454 2760 1459 2816
rect 0 2758 1459 2760
rect 0 2728 800 2758
rect 1393 2755 1459 2758
rect 6188 2752 6508 2753
rect 6188 2688 6196 2752
rect 6260 2688 6276 2752
rect 6340 2688 6356 2752
rect 6420 2688 6436 2752
rect 6500 2688 6508 2752
rect 6188 2687 6508 2688
rect 11432 2752 11752 2753
rect 11432 2688 11440 2752
rect 11504 2688 11520 2752
rect 11584 2688 11600 2752
rect 11664 2688 11680 2752
rect 11744 2688 11752 2752
rect 11432 2687 11752 2688
rect 3566 2208 3886 2209
rect 3566 2144 3574 2208
rect 3638 2144 3654 2208
rect 3718 2144 3734 2208
rect 3798 2144 3814 2208
rect 3878 2144 3886 2208
rect 3566 2143 3886 2144
rect 8810 2208 9130 2209
rect 8810 2144 8818 2208
rect 8882 2144 8898 2208
rect 8962 2144 8978 2208
rect 9042 2144 9058 2208
rect 9122 2144 9130 2208
rect 8810 2143 9130 2144
rect 14054 2208 14374 2209
rect 14054 2144 14062 2208
rect 14126 2144 14142 2208
rect 14206 2144 14222 2208
rect 14286 2144 14302 2208
rect 14366 2144 14374 2208
rect 14054 2143 14374 2144
rect 16481 1458 16547 1461
rect 17227 1458 18027 1488
rect 16481 1456 18027 1458
rect 16481 1400 16486 1456
rect 16542 1400 18027 1456
rect 16481 1398 18027 1400
rect 16481 1395 16547 1398
rect 17227 1368 18027 1398
<< via3 >>
rect 6196 17980 6260 17984
rect 6196 17924 6200 17980
rect 6200 17924 6256 17980
rect 6256 17924 6260 17980
rect 6196 17920 6260 17924
rect 6276 17980 6340 17984
rect 6276 17924 6280 17980
rect 6280 17924 6336 17980
rect 6336 17924 6340 17980
rect 6276 17920 6340 17924
rect 6356 17980 6420 17984
rect 6356 17924 6360 17980
rect 6360 17924 6416 17980
rect 6416 17924 6420 17980
rect 6356 17920 6420 17924
rect 6436 17980 6500 17984
rect 6436 17924 6440 17980
rect 6440 17924 6496 17980
rect 6496 17924 6500 17980
rect 6436 17920 6500 17924
rect 11440 17980 11504 17984
rect 11440 17924 11444 17980
rect 11444 17924 11500 17980
rect 11500 17924 11504 17980
rect 11440 17920 11504 17924
rect 11520 17980 11584 17984
rect 11520 17924 11524 17980
rect 11524 17924 11580 17980
rect 11580 17924 11584 17980
rect 11520 17920 11584 17924
rect 11600 17980 11664 17984
rect 11600 17924 11604 17980
rect 11604 17924 11660 17980
rect 11660 17924 11664 17980
rect 11600 17920 11664 17924
rect 11680 17980 11744 17984
rect 11680 17924 11684 17980
rect 11684 17924 11740 17980
rect 11740 17924 11744 17980
rect 11680 17920 11744 17924
rect 3574 17436 3638 17440
rect 3574 17380 3578 17436
rect 3578 17380 3634 17436
rect 3634 17380 3638 17436
rect 3574 17376 3638 17380
rect 3654 17436 3718 17440
rect 3654 17380 3658 17436
rect 3658 17380 3714 17436
rect 3714 17380 3718 17436
rect 3654 17376 3718 17380
rect 3734 17436 3798 17440
rect 3734 17380 3738 17436
rect 3738 17380 3794 17436
rect 3794 17380 3798 17436
rect 3734 17376 3798 17380
rect 3814 17436 3878 17440
rect 3814 17380 3818 17436
rect 3818 17380 3874 17436
rect 3874 17380 3878 17436
rect 3814 17376 3878 17380
rect 8818 17436 8882 17440
rect 8818 17380 8822 17436
rect 8822 17380 8878 17436
rect 8878 17380 8882 17436
rect 8818 17376 8882 17380
rect 8898 17436 8962 17440
rect 8898 17380 8902 17436
rect 8902 17380 8958 17436
rect 8958 17380 8962 17436
rect 8898 17376 8962 17380
rect 8978 17436 9042 17440
rect 8978 17380 8982 17436
rect 8982 17380 9038 17436
rect 9038 17380 9042 17436
rect 8978 17376 9042 17380
rect 9058 17436 9122 17440
rect 9058 17380 9062 17436
rect 9062 17380 9118 17436
rect 9118 17380 9122 17436
rect 9058 17376 9122 17380
rect 14062 17436 14126 17440
rect 14062 17380 14066 17436
rect 14066 17380 14122 17436
rect 14122 17380 14126 17436
rect 14062 17376 14126 17380
rect 14142 17436 14206 17440
rect 14142 17380 14146 17436
rect 14146 17380 14202 17436
rect 14202 17380 14206 17436
rect 14142 17376 14206 17380
rect 14222 17436 14286 17440
rect 14222 17380 14226 17436
rect 14226 17380 14282 17436
rect 14282 17380 14286 17436
rect 14222 17376 14286 17380
rect 14302 17436 14366 17440
rect 14302 17380 14306 17436
rect 14306 17380 14362 17436
rect 14362 17380 14366 17436
rect 14302 17376 14366 17380
rect 6196 16892 6260 16896
rect 6196 16836 6200 16892
rect 6200 16836 6256 16892
rect 6256 16836 6260 16892
rect 6196 16832 6260 16836
rect 6276 16892 6340 16896
rect 6276 16836 6280 16892
rect 6280 16836 6336 16892
rect 6336 16836 6340 16892
rect 6276 16832 6340 16836
rect 6356 16892 6420 16896
rect 6356 16836 6360 16892
rect 6360 16836 6416 16892
rect 6416 16836 6420 16892
rect 6356 16832 6420 16836
rect 6436 16892 6500 16896
rect 6436 16836 6440 16892
rect 6440 16836 6496 16892
rect 6496 16836 6500 16892
rect 6436 16832 6500 16836
rect 11440 16892 11504 16896
rect 11440 16836 11444 16892
rect 11444 16836 11500 16892
rect 11500 16836 11504 16892
rect 11440 16832 11504 16836
rect 11520 16892 11584 16896
rect 11520 16836 11524 16892
rect 11524 16836 11580 16892
rect 11580 16836 11584 16892
rect 11520 16832 11584 16836
rect 11600 16892 11664 16896
rect 11600 16836 11604 16892
rect 11604 16836 11660 16892
rect 11660 16836 11664 16892
rect 11600 16832 11664 16836
rect 11680 16892 11744 16896
rect 11680 16836 11684 16892
rect 11684 16836 11740 16892
rect 11740 16836 11744 16892
rect 11680 16832 11744 16836
rect 3574 16348 3638 16352
rect 3574 16292 3578 16348
rect 3578 16292 3634 16348
rect 3634 16292 3638 16348
rect 3574 16288 3638 16292
rect 3654 16348 3718 16352
rect 3654 16292 3658 16348
rect 3658 16292 3714 16348
rect 3714 16292 3718 16348
rect 3654 16288 3718 16292
rect 3734 16348 3798 16352
rect 3734 16292 3738 16348
rect 3738 16292 3794 16348
rect 3794 16292 3798 16348
rect 3734 16288 3798 16292
rect 3814 16348 3878 16352
rect 3814 16292 3818 16348
rect 3818 16292 3874 16348
rect 3874 16292 3878 16348
rect 3814 16288 3878 16292
rect 8818 16348 8882 16352
rect 8818 16292 8822 16348
rect 8822 16292 8878 16348
rect 8878 16292 8882 16348
rect 8818 16288 8882 16292
rect 8898 16348 8962 16352
rect 8898 16292 8902 16348
rect 8902 16292 8958 16348
rect 8958 16292 8962 16348
rect 8898 16288 8962 16292
rect 8978 16348 9042 16352
rect 8978 16292 8982 16348
rect 8982 16292 9038 16348
rect 9038 16292 9042 16348
rect 8978 16288 9042 16292
rect 9058 16348 9122 16352
rect 9058 16292 9062 16348
rect 9062 16292 9118 16348
rect 9118 16292 9122 16348
rect 9058 16288 9122 16292
rect 14062 16348 14126 16352
rect 14062 16292 14066 16348
rect 14066 16292 14122 16348
rect 14122 16292 14126 16348
rect 14062 16288 14126 16292
rect 14142 16348 14206 16352
rect 14142 16292 14146 16348
rect 14146 16292 14202 16348
rect 14202 16292 14206 16348
rect 14142 16288 14206 16292
rect 14222 16348 14286 16352
rect 14222 16292 14226 16348
rect 14226 16292 14282 16348
rect 14282 16292 14286 16348
rect 14222 16288 14286 16292
rect 14302 16348 14366 16352
rect 14302 16292 14306 16348
rect 14306 16292 14362 16348
rect 14362 16292 14366 16348
rect 14302 16288 14366 16292
rect 6196 15804 6260 15808
rect 6196 15748 6200 15804
rect 6200 15748 6256 15804
rect 6256 15748 6260 15804
rect 6196 15744 6260 15748
rect 6276 15804 6340 15808
rect 6276 15748 6280 15804
rect 6280 15748 6336 15804
rect 6336 15748 6340 15804
rect 6276 15744 6340 15748
rect 6356 15804 6420 15808
rect 6356 15748 6360 15804
rect 6360 15748 6416 15804
rect 6416 15748 6420 15804
rect 6356 15744 6420 15748
rect 6436 15804 6500 15808
rect 6436 15748 6440 15804
rect 6440 15748 6496 15804
rect 6496 15748 6500 15804
rect 6436 15744 6500 15748
rect 11440 15804 11504 15808
rect 11440 15748 11444 15804
rect 11444 15748 11500 15804
rect 11500 15748 11504 15804
rect 11440 15744 11504 15748
rect 11520 15804 11584 15808
rect 11520 15748 11524 15804
rect 11524 15748 11580 15804
rect 11580 15748 11584 15804
rect 11520 15744 11584 15748
rect 11600 15804 11664 15808
rect 11600 15748 11604 15804
rect 11604 15748 11660 15804
rect 11660 15748 11664 15804
rect 11600 15744 11664 15748
rect 11680 15804 11744 15808
rect 11680 15748 11684 15804
rect 11684 15748 11740 15804
rect 11740 15748 11744 15804
rect 11680 15744 11744 15748
rect 3574 15260 3638 15264
rect 3574 15204 3578 15260
rect 3578 15204 3634 15260
rect 3634 15204 3638 15260
rect 3574 15200 3638 15204
rect 3654 15260 3718 15264
rect 3654 15204 3658 15260
rect 3658 15204 3714 15260
rect 3714 15204 3718 15260
rect 3654 15200 3718 15204
rect 3734 15260 3798 15264
rect 3734 15204 3738 15260
rect 3738 15204 3794 15260
rect 3794 15204 3798 15260
rect 3734 15200 3798 15204
rect 3814 15260 3878 15264
rect 3814 15204 3818 15260
rect 3818 15204 3874 15260
rect 3874 15204 3878 15260
rect 3814 15200 3878 15204
rect 8818 15260 8882 15264
rect 8818 15204 8822 15260
rect 8822 15204 8878 15260
rect 8878 15204 8882 15260
rect 8818 15200 8882 15204
rect 8898 15260 8962 15264
rect 8898 15204 8902 15260
rect 8902 15204 8958 15260
rect 8958 15204 8962 15260
rect 8898 15200 8962 15204
rect 8978 15260 9042 15264
rect 8978 15204 8982 15260
rect 8982 15204 9038 15260
rect 9038 15204 9042 15260
rect 8978 15200 9042 15204
rect 9058 15260 9122 15264
rect 9058 15204 9062 15260
rect 9062 15204 9118 15260
rect 9118 15204 9122 15260
rect 9058 15200 9122 15204
rect 14062 15260 14126 15264
rect 14062 15204 14066 15260
rect 14066 15204 14122 15260
rect 14122 15204 14126 15260
rect 14062 15200 14126 15204
rect 14142 15260 14206 15264
rect 14142 15204 14146 15260
rect 14146 15204 14202 15260
rect 14202 15204 14206 15260
rect 14142 15200 14206 15204
rect 14222 15260 14286 15264
rect 14222 15204 14226 15260
rect 14226 15204 14282 15260
rect 14282 15204 14286 15260
rect 14222 15200 14286 15204
rect 14302 15260 14366 15264
rect 14302 15204 14306 15260
rect 14306 15204 14362 15260
rect 14362 15204 14366 15260
rect 14302 15200 14366 15204
rect 6196 14716 6260 14720
rect 6196 14660 6200 14716
rect 6200 14660 6256 14716
rect 6256 14660 6260 14716
rect 6196 14656 6260 14660
rect 6276 14716 6340 14720
rect 6276 14660 6280 14716
rect 6280 14660 6336 14716
rect 6336 14660 6340 14716
rect 6276 14656 6340 14660
rect 6356 14716 6420 14720
rect 6356 14660 6360 14716
rect 6360 14660 6416 14716
rect 6416 14660 6420 14716
rect 6356 14656 6420 14660
rect 6436 14716 6500 14720
rect 6436 14660 6440 14716
rect 6440 14660 6496 14716
rect 6496 14660 6500 14716
rect 6436 14656 6500 14660
rect 11440 14716 11504 14720
rect 11440 14660 11444 14716
rect 11444 14660 11500 14716
rect 11500 14660 11504 14716
rect 11440 14656 11504 14660
rect 11520 14716 11584 14720
rect 11520 14660 11524 14716
rect 11524 14660 11580 14716
rect 11580 14660 11584 14716
rect 11520 14656 11584 14660
rect 11600 14716 11664 14720
rect 11600 14660 11604 14716
rect 11604 14660 11660 14716
rect 11660 14660 11664 14716
rect 11600 14656 11664 14660
rect 11680 14716 11744 14720
rect 11680 14660 11684 14716
rect 11684 14660 11740 14716
rect 11740 14660 11744 14716
rect 11680 14656 11744 14660
rect 3574 14172 3638 14176
rect 3574 14116 3578 14172
rect 3578 14116 3634 14172
rect 3634 14116 3638 14172
rect 3574 14112 3638 14116
rect 3654 14172 3718 14176
rect 3654 14116 3658 14172
rect 3658 14116 3714 14172
rect 3714 14116 3718 14172
rect 3654 14112 3718 14116
rect 3734 14172 3798 14176
rect 3734 14116 3738 14172
rect 3738 14116 3794 14172
rect 3794 14116 3798 14172
rect 3734 14112 3798 14116
rect 3814 14172 3878 14176
rect 3814 14116 3818 14172
rect 3818 14116 3874 14172
rect 3874 14116 3878 14172
rect 3814 14112 3878 14116
rect 8818 14172 8882 14176
rect 8818 14116 8822 14172
rect 8822 14116 8878 14172
rect 8878 14116 8882 14172
rect 8818 14112 8882 14116
rect 8898 14172 8962 14176
rect 8898 14116 8902 14172
rect 8902 14116 8958 14172
rect 8958 14116 8962 14172
rect 8898 14112 8962 14116
rect 8978 14172 9042 14176
rect 8978 14116 8982 14172
rect 8982 14116 9038 14172
rect 9038 14116 9042 14172
rect 8978 14112 9042 14116
rect 9058 14172 9122 14176
rect 9058 14116 9062 14172
rect 9062 14116 9118 14172
rect 9118 14116 9122 14172
rect 9058 14112 9122 14116
rect 14062 14172 14126 14176
rect 14062 14116 14066 14172
rect 14066 14116 14122 14172
rect 14122 14116 14126 14172
rect 14062 14112 14126 14116
rect 14142 14172 14206 14176
rect 14142 14116 14146 14172
rect 14146 14116 14202 14172
rect 14202 14116 14206 14172
rect 14142 14112 14206 14116
rect 14222 14172 14286 14176
rect 14222 14116 14226 14172
rect 14226 14116 14282 14172
rect 14282 14116 14286 14172
rect 14222 14112 14286 14116
rect 14302 14172 14366 14176
rect 14302 14116 14306 14172
rect 14306 14116 14362 14172
rect 14362 14116 14366 14172
rect 14302 14112 14366 14116
rect 6196 13628 6260 13632
rect 6196 13572 6200 13628
rect 6200 13572 6256 13628
rect 6256 13572 6260 13628
rect 6196 13568 6260 13572
rect 6276 13628 6340 13632
rect 6276 13572 6280 13628
rect 6280 13572 6336 13628
rect 6336 13572 6340 13628
rect 6276 13568 6340 13572
rect 6356 13628 6420 13632
rect 6356 13572 6360 13628
rect 6360 13572 6416 13628
rect 6416 13572 6420 13628
rect 6356 13568 6420 13572
rect 6436 13628 6500 13632
rect 6436 13572 6440 13628
rect 6440 13572 6496 13628
rect 6496 13572 6500 13628
rect 6436 13568 6500 13572
rect 11440 13628 11504 13632
rect 11440 13572 11444 13628
rect 11444 13572 11500 13628
rect 11500 13572 11504 13628
rect 11440 13568 11504 13572
rect 11520 13628 11584 13632
rect 11520 13572 11524 13628
rect 11524 13572 11580 13628
rect 11580 13572 11584 13628
rect 11520 13568 11584 13572
rect 11600 13628 11664 13632
rect 11600 13572 11604 13628
rect 11604 13572 11660 13628
rect 11660 13572 11664 13628
rect 11600 13568 11664 13572
rect 11680 13628 11744 13632
rect 11680 13572 11684 13628
rect 11684 13572 11740 13628
rect 11740 13572 11744 13628
rect 11680 13568 11744 13572
rect 3574 13084 3638 13088
rect 3574 13028 3578 13084
rect 3578 13028 3634 13084
rect 3634 13028 3638 13084
rect 3574 13024 3638 13028
rect 3654 13084 3718 13088
rect 3654 13028 3658 13084
rect 3658 13028 3714 13084
rect 3714 13028 3718 13084
rect 3654 13024 3718 13028
rect 3734 13084 3798 13088
rect 3734 13028 3738 13084
rect 3738 13028 3794 13084
rect 3794 13028 3798 13084
rect 3734 13024 3798 13028
rect 3814 13084 3878 13088
rect 3814 13028 3818 13084
rect 3818 13028 3874 13084
rect 3874 13028 3878 13084
rect 3814 13024 3878 13028
rect 8818 13084 8882 13088
rect 8818 13028 8822 13084
rect 8822 13028 8878 13084
rect 8878 13028 8882 13084
rect 8818 13024 8882 13028
rect 8898 13084 8962 13088
rect 8898 13028 8902 13084
rect 8902 13028 8958 13084
rect 8958 13028 8962 13084
rect 8898 13024 8962 13028
rect 8978 13084 9042 13088
rect 8978 13028 8982 13084
rect 8982 13028 9038 13084
rect 9038 13028 9042 13084
rect 8978 13024 9042 13028
rect 9058 13084 9122 13088
rect 9058 13028 9062 13084
rect 9062 13028 9118 13084
rect 9118 13028 9122 13084
rect 9058 13024 9122 13028
rect 14062 13084 14126 13088
rect 14062 13028 14066 13084
rect 14066 13028 14122 13084
rect 14122 13028 14126 13084
rect 14062 13024 14126 13028
rect 14142 13084 14206 13088
rect 14142 13028 14146 13084
rect 14146 13028 14202 13084
rect 14202 13028 14206 13084
rect 14142 13024 14206 13028
rect 14222 13084 14286 13088
rect 14222 13028 14226 13084
rect 14226 13028 14282 13084
rect 14282 13028 14286 13084
rect 14222 13024 14286 13028
rect 14302 13084 14366 13088
rect 14302 13028 14306 13084
rect 14306 13028 14362 13084
rect 14362 13028 14366 13084
rect 14302 13024 14366 13028
rect 6196 12540 6260 12544
rect 6196 12484 6200 12540
rect 6200 12484 6256 12540
rect 6256 12484 6260 12540
rect 6196 12480 6260 12484
rect 6276 12540 6340 12544
rect 6276 12484 6280 12540
rect 6280 12484 6336 12540
rect 6336 12484 6340 12540
rect 6276 12480 6340 12484
rect 6356 12540 6420 12544
rect 6356 12484 6360 12540
rect 6360 12484 6416 12540
rect 6416 12484 6420 12540
rect 6356 12480 6420 12484
rect 6436 12540 6500 12544
rect 6436 12484 6440 12540
rect 6440 12484 6496 12540
rect 6496 12484 6500 12540
rect 6436 12480 6500 12484
rect 11440 12540 11504 12544
rect 11440 12484 11444 12540
rect 11444 12484 11500 12540
rect 11500 12484 11504 12540
rect 11440 12480 11504 12484
rect 11520 12540 11584 12544
rect 11520 12484 11524 12540
rect 11524 12484 11580 12540
rect 11580 12484 11584 12540
rect 11520 12480 11584 12484
rect 11600 12540 11664 12544
rect 11600 12484 11604 12540
rect 11604 12484 11660 12540
rect 11660 12484 11664 12540
rect 11600 12480 11664 12484
rect 11680 12540 11744 12544
rect 11680 12484 11684 12540
rect 11684 12484 11740 12540
rect 11740 12484 11744 12540
rect 11680 12480 11744 12484
rect 3574 11996 3638 12000
rect 3574 11940 3578 11996
rect 3578 11940 3634 11996
rect 3634 11940 3638 11996
rect 3574 11936 3638 11940
rect 3654 11996 3718 12000
rect 3654 11940 3658 11996
rect 3658 11940 3714 11996
rect 3714 11940 3718 11996
rect 3654 11936 3718 11940
rect 3734 11996 3798 12000
rect 3734 11940 3738 11996
rect 3738 11940 3794 11996
rect 3794 11940 3798 11996
rect 3734 11936 3798 11940
rect 3814 11996 3878 12000
rect 3814 11940 3818 11996
rect 3818 11940 3874 11996
rect 3874 11940 3878 11996
rect 3814 11936 3878 11940
rect 8818 11996 8882 12000
rect 8818 11940 8822 11996
rect 8822 11940 8878 11996
rect 8878 11940 8882 11996
rect 8818 11936 8882 11940
rect 8898 11996 8962 12000
rect 8898 11940 8902 11996
rect 8902 11940 8958 11996
rect 8958 11940 8962 11996
rect 8898 11936 8962 11940
rect 8978 11996 9042 12000
rect 8978 11940 8982 11996
rect 8982 11940 9038 11996
rect 9038 11940 9042 11996
rect 8978 11936 9042 11940
rect 9058 11996 9122 12000
rect 9058 11940 9062 11996
rect 9062 11940 9118 11996
rect 9118 11940 9122 11996
rect 9058 11936 9122 11940
rect 14062 11996 14126 12000
rect 14062 11940 14066 11996
rect 14066 11940 14122 11996
rect 14122 11940 14126 11996
rect 14062 11936 14126 11940
rect 14142 11996 14206 12000
rect 14142 11940 14146 11996
rect 14146 11940 14202 11996
rect 14202 11940 14206 11996
rect 14142 11936 14206 11940
rect 14222 11996 14286 12000
rect 14222 11940 14226 11996
rect 14226 11940 14282 11996
rect 14282 11940 14286 11996
rect 14222 11936 14286 11940
rect 14302 11996 14366 12000
rect 14302 11940 14306 11996
rect 14306 11940 14362 11996
rect 14362 11940 14366 11996
rect 14302 11936 14366 11940
rect 6196 11452 6260 11456
rect 6196 11396 6200 11452
rect 6200 11396 6256 11452
rect 6256 11396 6260 11452
rect 6196 11392 6260 11396
rect 6276 11452 6340 11456
rect 6276 11396 6280 11452
rect 6280 11396 6336 11452
rect 6336 11396 6340 11452
rect 6276 11392 6340 11396
rect 6356 11452 6420 11456
rect 6356 11396 6360 11452
rect 6360 11396 6416 11452
rect 6416 11396 6420 11452
rect 6356 11392 6420 11396
rect 6436 11452 6500 11456
rect 6436 11396 6440 11452
rect 6440 11396 6496 11452
rect 6496 11396 6500 11452
rect 6436 11392 6500 11396
rect 11440 11452 11504 11456
rect 11440 11396 11444 11452
rect 11444 11396 11500 11452
rect 11500 11396 11504 11452
rect 11440 11392 11504 11396
rect 11520 11452 11584 11456
rect 11520 11396 11524 11452
rect 11524 11396 11580 11452
rect 11580 11396 11584 11452
rect 11520 11392 11584 11396
rect 11600 11452 11664 11456
rect 11600 11396 11604 11452
rect 11604 11396 11660 11452
rect 11660 11396 11664 11452
rect 11600 11392 11664 11396
rect 11680 11452 11744 11456
rect 11680 11396 11684 11452
rect 11684 11396 11740 11452
rect 11740 11396 11744 11452
rect 11680 11392 11744 11396
rect 3574 10908 3638 10912
rect 3574 10852 3578 10908
rect 3578 10852 3634 10908
rect 3634 10852 3638 10908
rect 3574 10848 3638 10852
rect 3654 10908 3718 10912
rect 3654 10852 3658 10908
rect 3658 10852 3714 10908
rect 3714 10852 3718 10908
rect 3654 10848 3718 10852
rect 3734 10908 3798 10912
rect 3734 10852 3738 10908
rect 3738 10852 3794 10908
rect 3794 10852 3798 10908
rect 3734 10848 3798 10852
rect 3814 10908 3878 10912
rect 3814 10852 3818 10908
rect 3818 10852 3874 10908
rect 3874 10852 3878 10908
rect 3814 10848 3878 10852
rect 8818 10908 8882 10912
rect 8818 10852 8822 10908
rect 8822 10852 8878 10908
rect 8878 10852 8882 10908
rect 8818 10848 8882 10852
rect 8898 10908 8962 10912
rect 8898 10852 8902 10908
rect 8902 10852 8958 10908
rect 8958 10852 8962 10908
rect 8898 10848 8962 10852
rect 8978 10908 9042 10912
rect 8978 10852 8982 10908
rect 8982 10852 9038 10908
rect 9038 10852 9042 10908
rect 8978 10848 9042 10852
rect 9058 10908 9122 10912
rect 9058 10852 9062 10908
rect 9062 10852 9118 10908
rect 9118 10852 9122 10908
rect 9058 10848 9122 10852
rect 14062 10908 14126 10912
rect 14062 10852 14066 10908
rect 14066 10852 14122 10908
rect 14122 10852 14126 10908
rect 14062 10848 14126 10852
rect 14142 10908 14206 10912
rect 14142 10852 14146 10908
rect 14146 10852 14202 10908
rect 14202 10852 14206 10908
rect 14142 10848 14206 10852
rect 14222 10908 14286 10912
rect 14222 10852 14226 10908
rect 14226 10852 14282 10908
rect 14282 10852 14286 10908
rect 14222 10848 14286 10852
rect 14302 10908 14366 10912
rect 14302 10852 14306 10908
rect 14306 10852 14362 10908
rect 14362 10852 14366 10908
rect 14302 10848 14366 10852
rect 6196 10364 6260 10368
rect 6196 10308 6200 10364
rect 6200 10308 6256 10364
rect 6256 10308 6260 10364
rect 6196 10304 6260 10308
rect 6276 10364 6340 10368
rect 6276 10308 6280 10364
rect 6280 10308 6336 10364
rect 6336 10308 6340 10364
rect 6276 10304 6340 10308
rect 6356 10364 6420 10368
rect 6356 10308 6360 10364
rect 6360 10308 6416 10364
rect 6416 10308 6420 10364
rect 6356 10304 6420 10308
rect 6436 10364 6500 10368
rect 6436 10308 6440 10364
rect 6440 10308 6496 10364
rect 6496 10308 6500 10364
rect 6436 10304 6500 10308
rect 11440 10364 11504 10368
rect 11440 10308 11444 10364
rect 11444 10308 11500 10364
rect 11500 10308 11504 10364
rect 11440 10304 11504 10308
rect 11520 10364 11584 10368
rect 11520 10308 11524 10364
rect 11524 10308 11580 10364
rect 11580 10308 11584 10364
rect 11520 10304 11584 10308
rect 11600 10364 11664 10368
rect 11600 10308 11604 10364
rect 11604 10308 11660 10364
rect 11660 10308 11664 10364
rect 11600 10304 11664 10308
rect 11680 10364 11744 10368
rect 11680 10308 11684 10364
rect 11684 10308 11740 10364
rect 11740 10308 11744 10364
rect 11680 10304 11744 10308
rect 3574 9820 3638 9824
rect 3574 9764 3578 9820
rect 3578 9764 3634 9820
rect 3634 9764 3638 9820
rect 3574 9760 3638 9764
rect 3654 9820 3718 9824
rect 3654 9764 3658 9820
rect 3658 9764 3714 9820
rect 3714 9764 3718 9820
rect 3654 9760 3718 9764
rect 3734 9820 3798 9824
rect 3734 9764 3738 9820
rect 3738 9764 3794 9820
rect 3794 9764 3798 9820
rect 3734 9760 3798 9764
rect 3814 9820 3878 9824
rect 3814 9764 3818 9820
rect 3818 9764 3874 9820
rect 3874 9764 3878 9820
rect 3814 9760 3878 9764
rect 8818 9820 8882 9824
rect 8818 9764 8822 9820
rect 8822 9764 8878 9820
rect 8878 9764 8882 9820
rect 8818 9760 8882 9764
rect 8898 9820 8962 9824
rect 8898 9764 8902 9820
rect 8902 9764 8958 9820
rect 8958 9764 8962 9820
rect 8898 9760 8962 9764
rect 8978 9820 9042 9824
rect 8978 9764 8982 9820
rect 8982 9764 9038 9820
rect 9038 9764 9042 9820
rect 8978 9760 9042 9764
rect 9058 9820 9122 9824
rect 9058 9764 9062 9820
rect 9062 9764 9118 9820
rect 9118 9764 9122 9820
rect 9058 9760 9122 9764
rect 14062 9820 14126 9824
rect 14062 9764 14066 9820
rect 14066 9764 14122 9820
rect 14122 9764 14126 9820
rect 14062 9760 14126 9764
rect 14142 9820 14206 9824
rect 14142 9764 14146 9820
rect 14146 9764 14202 9820
rect 14202 9764 14206 9820
rect 14142 9760 14206 9764
rect 14222 9820 14286 9824
rect 14222 9764 14226 9820
rect 14226 9764 14282 9820
rect 14282 9764 14286 9820
rect 14222 9760 14286 9764
rect 14302 9820 14366 9824
rect 14302 9764 14306 9820
rect 14306 9764 14362 9820
rect 14362 9764 14366 9820
rect 14302 9760 14366 9764
rect 6196 9276 6260 9280
rect 6196 9220 6200 9276
rect 6200 9220 6256 9276
rect 6256 9220 6260 9276
rect 6196 9216 6260 9220
rect 6276 9276 6340 9280
rect 6276 9220 6280 9276
rect 6280 9220 6336 9276
rect 6336 9220 6340 9276
rect 6276 9216 6340 9220
rect 6356 9276 6420 9280
rect 6356 9220 6360 9276
rect 6360 9220 6416 9276
rect 6416 9220 6420 9276
rect 6356 9216 6420 9220
rect 6436 9276 6500 9280
rect 6436 9220 6440 9276
rect 6440 9220 6496 9276
rect 6496 9220 6500 9276
rect 6436 9216 6500 9220
rect 11440 9276 11504 9280
rect 11440 9220 11444 9276
rect 11444 9220 11500 9276
rect 11500 9220 11504 9276
rect 11440 9216 11504 9220
rect 11520 9276 11584 9280
rect 11520 9220 11524 9276
rect 11524 9220 11580 9276
rect 11580 9220 11584 9276
rect 11520 9216 11584 9220
rect 11600 9276 11664 9280
rect 11600 9220 11604 9276
rect 11604 9220 11660 9276
rect 11660 9220 11664 9276
rect 11600 9216 11664 9220
rect 11680 9276 11744 9280
rect 11680 9220 11684 9276
rect 11684 9220 11740 9276
rect 11740 9220 11744 9276
rect 11680 9216 11744 9220
rect 3574 8732 3638 8736
rect 3574 8676 3578 8732
rect 3578 8676 3634 8732
rect 3634 8676 3638 8732
rect 3574 8672 3638 8676
rect 3654 8732 3718 8736
rect 3654 8676 3658 8732
rect 3658 8676 3714 8732
rect 3714 8676 3718 8732
rect 3654 8672 3718 8676
rect 3734 8732 3798 8736
rect 3734 8676 3738 8732
rect 3738 8676 3794 8732
rect 3794 8676 3798 8732
rect 3734 8672 3798 8676
rect 3814 8732 3878 8736
rect 3814 8676 3818 8732
rect 3818 8676 3874 8732
rect 3874 8676 3878 8732
rect 3814 8672 3878 8676
rect 8818 8732 8882 8736
rect 8818 8676 8822 8732
rect 8822 8676 8878 8732
rect 8878 8676 8882 8732
rect 8818 8672 8882 8676
rect 8898 8732 8962 8736
rect 8898 8676 8902 8732
rect 8902 8676 8958 8732
rect 8958 8676 8962 8732
rect 8898 8672 8962 8676
rect 8978 8732 9042 8736
rect 8978 8676 8982 8732
rect 8982 8676 9038 8732
rect 9038 8676 9042 8732
rect 8978 8672 9042 8676
rect 9058 8732 9122 8736
rect 9058 8676 9062 8732
rect 9062 8676 9118 8732
rect 9118 8676 9122 8732
rect 9058 8672 9122 8676
rect 14062 8732 14126 8736
rect 14062 8676 14066 8732
rect 14066 8676 14122 8732
rect 14122 8676 14126 8732
rect 14062 8672 14126 8676
rect 14142 8732 14206 8736
rect 14142 8676 14146 8732
rect 14146 8676 14202 8732
rect 14202 8676 14206 8732
rect 14142 8672 14206 8676
rect 14222 8732 14286 8736
rect 14222 8676 14226 8732
rect 14226 8676 14282 8732
rect 14282 8676 14286 8732
rect 14222 8672 14286 8676
rect 14302 8732 14366 8736
rect 14302 8676 14306 8732
rect 14306 8676 14362 8732
rect 14362 8676 14366 8732
rect 14302 8672 14366 8676
rect 6196 8188 6260 8192
rect 6196 8132 6200 8188
rect 6200 8132 6256 8188
rect 6256 8132 6260 8188
rect 6196 8128 6260 8132
rect 6276 8188 6340 8192
rect 6276 8132 6280 8188
rect 6280 8132 6336 8188
rect 6336 8132 6340 8188
rect 6276 8128 6340 8132
rect 6356 8188 6420 8192
rect 6356 8132 6360 8188
rect 6360 8132 6416 8188
rect 6416 8132 6420 8188
rect 6356 8128 6420 8132
rect 6436 8188 6500 8192
rect 6436 8132 6440 8188
rect 6440 8132 6496 8188
rect 6496 8132 6500 8188
rect 6436 8128 6500 8132
rect 11440 8188 11504 8192
rect 11440 8132 11444 8188
rect 11444 8132 11500 8188
rect 11500 8132 11504 8188
rect 11440 8128 11504 8132
rect 11520 8188 11584 8192
rect 11520 8132 11524 8188
rect 11524 8132 11580 8188
rect 11580 8132 11584 8188
rect 11520 8128 11584 8132
rect 11600 8188 11664 8192
rect 11600 8132 11604 8188
rect 11604 8132 11660 8188
rect 11660 8132 11664 8188
rect 11600 8128 11664 8132
rect 11680 8188 11744 8192
rect 11680 8132 11684 8188
rect 11684 8132 11740 8188
rect 11740 8132 11744 8188
rect 11680 8128 11744 8132
rect 3574 7644 3638 7648
rect 3574 7588 3578 7644
rect 3578 7588 3634 7644
rect 3634 7588 3638 7644
rect 3574 7584 3638 7588
rect 3654 7644 3718 7648
rect 3654 7588 3658 7644
rect 3658 7588 3714 7644
rect 3714 7588 3718 7644
rect 3654 7584 3718 7588
rect 3734 7644 3798 7648
rect 3734 7588 3738 7644
rect 3738 7588 3794 7644
rect 3794 7588 3798 7644
rect 3734 7584 3798 7588
rect 3814 7644 3878 7648
rect 3814 7588 3818 7644
rect 3818 7588 3874 7644
rect 3874 7588 3878 7644
rect 3814 7584 3878 7588
rect 8818 7644 8882 7648
rect 8818 7588 8822 7644
rect 8822 7588 8878 7644
rect 8878 7588 8882 7644
rect 8818 7584 8882 7588
rect 8898 7644 8962 7648
rect 8898 7588 8902 7644
rect 8902 7588 8958 7644
rect 8958 7588 8962 7644
rect 8898 7584 8962 7588
rect 8978 7644 9042 7648
rect 8978 7588 8982 7644
rect 8982 7588 9038 7644
rect 9038 7588 9042 7644
rect 8978 7584 9042 7588
rect 9058 7644 9122 7648
rect 9058 7588 9062 7644
rect 9062 7588 9118 7644
rect 9118 7588 9122 7644
rect 9058 7584 9122 7588
rect 14062 7644 14126 7648
rect 14062 7588 14066 7644
rect 14066 7588 14122 7644
rect 14122 7588 14126 7644
rect 14062 7584 14126 7588
rect 14142 7644 14206 7648
rect 14142 7588 14146 7644
rect 14146 7588 14202 7644
rect 14202 7588 14206 7644
rect 14142 7584 14206 7588
rect 14222 7644 14286 7648
rect 14222 7588 14226 7644
rect 14226 7588 14282 7644
rect 14282 7588 14286 7644
rect 14222 7584 14286 7588
rect 14302 7644 14366 7648
rect 14302 7588 14306 7644
rect 14306 7588 14362 7644
rect 14362 7588 14366 7644
rect 14302 7584 14366 7588
rect 6196 7100 6260 7104
rect 6196 7044 6200 7100
rect 6200 7044 6256 7100
rect 6256 7044 6260 7100
rect 6196 7040 6260 7044
rect 6276 7100 6340 7104
rect 6276 7044 6280 7100
rect 6280 7044 6336 7100
rect 6336 7044 6340 7100
rect 6276 7040 6340 7044
rect 6356 7100 6420 7104
rect 6356 7044 6360 7100
rect 6360 7044 6416 7100
rect 6416 7044 6420 7100
rect 6356 7040 6420 7044
rect 6436 7100 6500 7104
rect 6436 7044 6440 7100
rect 6440 7044 6496 7100
rect 6496 7044 6500 7100
rect 6436 7040 6500 7044
rect 11440 7100 11504 7104
rect 11440 7044 11444 7100
rect 11444 7044 11500 7100
rect 11500 7044 11504 7100
rect 11440 7040 11504 7044
rect 11520 7100 11584 7104
rect 11520 7044 11524 7100
rect 11524 7044 11580 7100
rect 11580 7044 11584 7100
rect 11520 7040 11584 7044
rect 11600 7100 11664 7104
rect 11600 7044 11604 7100
rect 11604 7044 11660 7100
rect 11660 7044 11664 7100
rect 11600 7040 11664 7044
rect 11680 7100 11744 7104
rect 11680 7044 11684 7100
rect 11684 7044 11740 7100
rect 11740 7044 11744 7100
rect 11680 7040 11744 7044
rect 3574 6556 3638 6560
rect 3574 6500 3578 6556
rect 3578 6500 3634 6556
rect 3634 6500 3638 6556
rect 3574 6496 3638 6500
rect 3654 6556 3718 6560
rect 3654 6500 3658 6556
rect 3658 6500 3714 6556
rect 3714 6500 3718 6556
rect 3654 6496 3718 6500
rect 3734 6556 3798 6560
rect 3734 6500 3738 6556
rect 3738 6500 3794 6556
rect 3794 6500 3798 6556
rect 3734 6496 3798 6500
rect 3814 6556 3878 6560
rect 3814 6500 3818 6556
rect 3818 6500 3874 6556
rect 3874 6500 3878 6556
rect 3814 6496 3878 6500
rect 8818 6556 8882 6560
rect 8818 6500 8822 6556
rect 8822 6500 8878 6556
rect 8878 6500 8882 6556
rect 8818 6496 8882 6500
rect 8898 6556 8962 6560
rect 8898 6500 8902 6556
rect 8902 6500 8958 6556
rect 8958 6500 8962 6556
rect 8898 6496 8962 6500
rect 8978 6556 9042 6560
rect 8978 6500 8982 6556
rect 8982 6500 9038 6556
rect 9038 6500 9042 6556
rect 8978 6496 9042 6500
rect 9058 6556 9122 6560
rect 9058 6500 9062 6556
rect 9062 6500 9118 6556
rect 9118 6500 9122 6556
rect 9058 6496 9122 6500
rect 14062 6556 14126 6560
rect 14062 6500 14066 6556
rect 14066 6500 14122 6556
rect 14122 6500 14126 6556
rect 14062 6496 14126 6500
rect 14142 6556 14206 6560
rect 14142 6500 14146 6556
rect 14146 6500 14202 6556
rect 14202 6500 14206 6556
rect 14142 6496 14206 6500
rect 14222 6556 14286 6560
rect 14222 6500 14226 6556
rect 14226 6500 14282 6556
rect 14282 6500 14286 6556
rect 14222 6496 14286 6500
rect 14302 6556 14366 6560
rect 14302 6500 14306 6556
rect 14306 6500 14362 6556
rect 14362 6500 14366 6556
rect 14302 6496 14366 6500
rect 6196 6012 6260 6016
rect 6196 5956 6200 6012
rect 6200 5956 6256 6012
rect 6256 5956 6260 6012
rect 6196 5952 6260 5956
rect 6276 6012 6340 6016
rect 6276 5956 6280 6012
rect 6280 5956 6336 6012
rect 6336 5956 6340 6012
rect 6276 5952 6340 5956
rect 6356 6012 6420 6016
rect 6356 5956 6360 6012
rect 6360 5956 6416 6012
rect 6416 5956 6420 6012
rect 6356 5952 6420 5956
rect 6436 6012 6500 6016
rect 6436 5956 6440 6012
rect 6440 5956 6496 6012
rect 6496 5956 6500 6012
rect 6436 5952 6500 5956
rect 11440 6012 11504 6016
rect 11440 5956 11444 6012
rect 11444 5956 11500 6012
rect 11500 5956 11504 6012
rect 11440 5952 11504 5956
rect 11520 6012 11584 6016
rect 11520 5956 11524 6012
rect 11524 5956 11580 6012
rect 11580 5956 11584 6012
rect 11520 5952 11584 5956
rect 11600 6012 11664 6016
rect 11600 5956 11604 6012
rect 11604 5956 11660 6012
rect 11660 5956 11664 6012
rect 11600 5952 11664 5956
rect 11680 6012 11744 6016
rect 11680 5956 11684 6012
rect 11684 5956 11740 6012
rect 11740 5956 11744 6012
rect 11680 5952 11744 5956
rect 3574 5468 3638 5472
rect 3574 5412 3578 5468
rect 3578 5412 3634 5468
rect 3634 5412 3638 5468
rect 3574 5408 3638 5412
rect 3654 5468 3718 5472
rect 3654 5412 3658 5468
rect 3658 5412 3714 5468
rect 3714 5412 3718 5468
rect 3654 5408 3718 5412
rect 3734 5468 3798 5472
rect 3734 5412 3738 5468
rect 3738 5412 3794 5468
rect 3794 5412 3798 5468
rect 3734 5408 3798 5412
rect 3814 5468 3878 5472
rect 3814 5412 3818 5468
rect 3818 5412 3874 5468
rect 3874 5412 3878 5468
rect 3814 5408 3878 5412
rect 8818 5468 8882 5472
rect 8818 5412 8822 5468
rect 8822 5412 8878 5468
rect 8878 5412 8882 5468
rect 8818 5408 8882 5412
rect 8898 5468 8962 5472
rect 8898 5412 8902 5468
rect 8902 5412 8958 5468
rect 8958 5412 8962 5468
rect 8898 5408 8962 5412
rect 8978 5468 9042 5472
rect 8978 5412 8982 5468
rect 8982 5412 9038 5468
rect 9038 5412 9042 5468
rect 8978 5408 9042 5412
rect 9058 5468 9122 5472
rect 9058 5412 9062 5468
rect 9062 5412 9118 5468
rect 9118 5412 9122 5468
rect 9058 5408 9122 5412
rect 14062 5468 14126 5472
rect 14062 5412 14066 5468
rect 14066 5412 14122 5468
rect 14122 5412 14126 5468
rect 14062 5408 14126 5412
rect 14142 5468 14206 5472
rect 14142 5412 14146 5468
rect 14146 5412 14202 5468
rect 14202 5412 14206 5468
rect 14142 5408 14206 5412
rect 14222 5468 14286 5472
rect 14222 5412 14226 5468
rect 14226 5412 14282 5468
rect 14282 5412 14286 5468
rect 14222 5408 14286 5412
rect 14302 5468 14366 5472
rect 14302 5412 14306 5468
rect 14306 5412 14362 5468
rect 14362 5412 14366 5468
rect 14302 5408 14366 5412
rect 6196 4924 6260 4928
rect 6196 4868 6200 4924
rect 6200 4868 6256 4924
rect 6256 4868 6260 4924
rect 6196 4864 6260 4868
rect 6276 4924 6340 4928
rect 6276 4868 6280 4924
rect 6280 4868 6336 4924
rect 6336 4868 6340 4924
rect 6276 4864 6340 4868
rect 6356 4924 6420 4928
rect 6356 4868 6360 4924
rect 6360 4868 6416 4924
rect 6416 4868 6420 4924
rect 6356 4864 6420 4868
rect 6436 4924 6500 4928
rect 6436 4868 6440 4924
rect 6440 4868 6496 4924
rect 6496 4868 6500 4924
rect 6436 4864 6500 4868
rect 11440 4924 11504 4928
rect 11440 4868 11444 4924
rect 11444 4868 11500 4924
rect 11500 4868 11504 4924
rect 11440 4864 11504 4868
rect 11520 4924 11584 4928
rect 11520 4868 11524 4924
rect 11524 4868 11580 4924
rect 11580 4868 11584 4924
rect 11520 4864 11584 4868
rect 11600 4924 11664 4928
rect 11600 4868 11604 4924
rect 11604 4868 11660 4924
rect 11660 4868 11664 4924
rect 11600 4864 11664 4868
rect 11680 4924 11744 4928
rect 11680 4868 11684 4924
rect 11684 4868 11740 4924
rect 11740 4868 11744 4924
rect 11680 4864 11744 4868
rect 3574 4380 3638 4384
rect 3574 4324 3578 4380
rect 3578 4324 3634 4380
rect 3634 4324 3638 4380
rect 3574 4320 3638 4324
rect 3654 4380 3718 4384
rect 3654 4324 3658 4380
rect 3658 4324 3714 4380
rect 3714 4324 3718 4380
rect 3654 4320 3718 4324
rect 3734 4380 3798 4384
rect 3734 4324 3738 4380
rect 3738 4324 3794 4380
rect 3794 4324 3798 4380
rect 3734 4320 3798 4324
rect 3814 4380 3878 4384
rect 3814 4324 3818 4380
rect 3818 4324 3874 4380
rect 3874 4324 3878 4380
rect 3814 4320 3878 4324
rect 8818 4380 8882 4384
rect 8818 4324 8822 4380
rect 8822 4324 8878 4380
rect 8878 4324 8882 4380
rect 8818 4320 8882 4324
rect 8898 4380 8962 4384
rect 8898 4324 8902 4380
rect 8902 4324 8958 4380
rect 8958 4324 8962 4380
rect 8898 4320 8962 4324
rect 8978 4380 9042 4384
rect 8978 4324 8982 4380
rect 8982 4324 9038 4380
rect 9038 4324 9042 4380
rect 8978 4320 9042 4324
rect 9058 4380 9122 4384
rect 9058 4324 9062 4380
rect 9062 4324 9118 4380
rect 9118 4324 9122 4380
rect 9058 4320 9122 4324
rect 14062 4380 14126 4384
rect 14062 4324 14066 4380
rect 14066 4324 14122 4380
rect 14122 4324 14126 4380
rect 14062 4320 14126 4324
rect 14142 4380 14206 4384
rect 14142 4324 14146 4380
rect 14146 4324 14202 4380
rect 14202 4324 14206 4380
rect 14142 4320 14206 4324
rect 14222 4380 14286 4384
rect 14222 4324 14226 4380
rect 14226 4324 14282 4380
rect 14282 4324 14286 4380
rect 14222 4320 14286 4324
rect 14302 4380 14366 4384
rect 14302 4324 14306 4380
rect 14306 4324 14362 4380
rect 14362 4324 14366 4380
rect 14302 4320 14366 4324
rect 6196 3836 6260 3840
rect 6196 3780 6200 3836
rect 6200 3780 6256 3836
rect 6256 3780 6260 3836
rect 6196 3776 6260 3780
rect 6276 3836 6340 3840
rect 6276 3780 6280 3836
rect 6280 3780 6336 3836
rect 6336 3780 6340 3836
rect 6276 3776 6340 3780
rect 6356 3836 6420 3840
rect 6356 3780 6360 3836
rect 6360 3780 6416 3836
rect 6416 3780 6420 3836
rect 6356 3776 6420 3780
rect 6436 3836 6500 3840
rect 6436 3780 6440 3836
rect 6440 3780 6496 3836
rect 6496 3780 6500 3836
rect 6436 3776 6500 3780
rect 11440 3836 11504 3840
rect 11440 3780 11444 3836
rect 11444 3780 11500 3836
rect 11500 3780 11504 3836
rect 11440 3776 11504 3780
rect 11520 3836 11584 3840
rect 11520 3780 11524 3836
rect 11524 3780 11580 3836
rect 11580 3780 11584 3836
rect 11520 3776 11584 3780
rect 11600 3836 11664 3840
rect 11600 3780 11604 3836
rect 11604 3780 11660 3836
rect 11660 3780 11664 3836
rect 11600 3776 11664 3780
rect 11680 3836 11744 3840
rect 11680 3780 11684 3836
rect 11684 3780 11740 3836
rect 11740 3780 11744 3836
rect 11680 3776 11744 3780
rect 3574 3292 3638 3296
rect 3574 3236 3578 3292
rect 3578 3236 3634 3292
rect 3634 3236 3638 3292
rect 3574 3232 3638 3236
rect 3654 3292 3718 3296
rect 3654 3236 3658 3292
rect 3658 3236 3714 3292
rect 3714 3236 3718 3292
rect 3654 3232 3718 3236
rect 3734 3292 3798 3296
rect 3734 3236 3738 3292
rect 3738 3236 3794 3292
rect 3794 3236 3798 3292
rect 3734 3232 3798 3236
rect 3814 3292 3878 3296
rect 3814 3236 3818 3292
rect 3818 3236 3874 3292
rect 3874 3236 3878 3292
rect 3814 3232 3878 3236
rect 8818 3292 8882 3296
rect 8818 3236 8822 3292
rect 8822 3236 8878 3292
rect 8878 3236 8882 3292
rect 8818 3232 8882 3236
rect 8898 3292 8962 3296
rect 8898 3236 8902 3292
rect 8902 3236 8958 3292
rect 8958 3236 8962 3292
rect 8898 3232 8962 3236
rect 8978 3292 9042 3296
rect 8978 3236 8982 3292
rect 8982 3236 9038 3292
rect 9038 3236 9042 3292
rect 8978 3232 9042 3236
rect 9058 3292 9122 3296
rect 9058 3236 9062 3292
rect 9062 3236 9118 3292
rect 9118 3236 9122 3292
rect 9058 3232 9122 3236
rect 14062 3292 14126 3296
rect 14062 3236 14066 3292
rect 14066 3236 14122 3292
rect 14122 3236 14126 3292
rect 14062 3232 14126 3236
rect 14142 3292 14206 3296
rect 14142 3236 14146 3292
rect 14146 3236 14202 3292
rect 14202 3236 14206 3292
rect 14142 3232 14206 3236
rect 14222 3292 14286 3296
rect 14222 3236 14226 3292
rect 14226 3236 14282 3292
rect 14282 3236 14286 3292
rect 14222 3232 14286 3236
rect 14302 3292 14366 3296
rect 14302 3236 14306 3292
rect 14306 3236 14362 3292
rect 14362 3236 14366 3292
rect 14302 3232 14366 3236
rect 6196 2748 6260 2752
rect 6196 2692 6200 2748
rect 6200 2692 6256 2748
rect 6256 2692 6260 2748
rect 6196 2688 6260 2692
rect 6276 2748 6340 2752
rect 6276 2692 6280 2748
rect 6280 2692 6336 2748
rect 6336 2692 6340 2748
rect 6276 2688 6340 2692
rect 6356 2748 6420 2752
rect 6356 2692 6360 2748
rect 6360 2692 6416 2748
rect 6416 2692 6420 2748
rect 6356 2688 6420 2692
rect 6436 2748 6500 2752
rect 6436 2692 6440 2748
rect 6440 2692 6496 2748
rect 6496 2692 6500 2748
rect 6436 2688 6500 2692
rect 11440 2748 11504 2752
rect 11440 2692 11444 2748
rect 11444 2692 11500 2748
rect 11500 2692 11504 2748
rect 11440 2688 11504 2692
rect 11520 2748 11584 2752
rect 11520 2692 11524 2748
rect 11524 2692 11580 2748
rect 11580 2692 11584 2748
rect 11520 2688 11584 2692
rect 11600 2748 11664 2752
rect 11600 2692 11604 2748
rect 11604 2692 11660 2748
rect 11660 2692 11664 2748
rect 11600 2688 11664 2692
rect 11680 2748 11744 2752
rect 11680 2692 11684 2748
rect 11684 2692 11740 2748
rect 11740 2692 11744 2748
rect 11680 2688 11744 2692
rect 3574 2204 3638 2208
rect 3574 2148 3578 2204
rect 3578 2148 3634 2204
rect 3634 2148 3638 2204
rect 3574 2144 3638 2148
rect 3654 2204 3718 2208
rect 3654 2148 3658 2204
rect 3658 2148 3714 2204
rect 3714 2148 3718 2204
rect 3654 2144 3718 2148
rect 3734 2204 3798 2208
rect 3734 2148 3738 2204
rect 3738 2148 3794 2204
rect 3794 2148 3798 2204
rect 3734 2144 3798 2148
rect 3814 2204 3878 2208
rect 3814 2148 3818 2204
rect 3818 2148 3874 2204
rect 3874 2148 3878 2204
rect 3814 2144 3878 2148
rect 8818 2204 8882 2208
rect 8818 2148 8822 2204
rect 8822 2148 8878 2204
rect 8878 2148 8882 2204
rect 8818 2144 8882 2148
rect 8898 2204 8962 2208
rect 8898 2148 8902 2204
rect 8902 2148 8958 2204
rect 8958 2148 8962 2204
rect 8898 2144 8962 2148
rect 8978 2204 9042 2208
rect 8978 2148 8982 2204
rect 8982 2148 9038 2204
rect 9038 2148 9042 2204
rect 8978 2144 9042 2148
rect 9058 2204 9122 2208
rect 9058 2148 9062 2204
rect 9062 2148 9118 2204
rect 9118 2148 9122 2204
rect 9058 2144 9122 2148
rect 14062 2204 14126 2208
rect 14062 2148 14066 2204
rect 14066 2148 14122 2204
rect 14122 2148 14126 2204
rect 14062 2144 14126 2148
rect 14142 2204 14206 2208
rect 14142 2148 14146 2204
rect 14146 2148 14202 2204
rect 14202 2148 14206 2204
rect 14142 2144 14206 2148
rect 14222 2204 14286 2208
rect 14222 2148 14226 2204
rect 14226 2148 14282 2204
rect 14282 2148 14286 2204
rect 14222 2144 14286 2148
rect 14302 2204 14366 2208
rect 14302 2148 14306 2204
rect 14306 2148 14362 2204
rect 14362 2148 14366 2204
rect 14302 2144 14366 2148
<< metal4 >>
rect 3566 17440 3886 18000
rect 3566 17376 3574 17440
rect 3638 17376 3654 17440
rect 3718 17376 3734 17440
rect 3798 17376 3814 17440
rect 3878 17376 3886 17440
rect 3566 16352 3886 17376
rect 3566 16288 3574 16352
rect 3638 16288 3654 16352
rect 3718 16288 3734 16352
rect 3798 16288 3814 16352
rect 3878 16288 3886 16352
rect 3566 15392 3886 16288
rect 3566 15264 3608 15392
rect 3844 15264 3886 15392
rect 3566 15200 3574 15264
rect 3878 15200 3886 15264
rect 3566 15156 3608 15200
rect 3844 15156 3886 15200
rect 3566 14176 3886 15156
rect 3566 14112 3574 14176
rect 3638 14112 3654 14176
rect 3718 14112 3734 14176
rect 3798 14112 3814 14176
rect 3878 14112 3886 14176
rect 3566 13088 3886 14112
rect 3566 13024 3574 13088
rect 3638 13024 3654 13088
rect 3718 13024 3734 13088
rect 3798 13024 3814 13088
rect 3878 13024 3886 13088
rect 3566 12000 3886 13024
rect 3566 11936 3574 12000
rect 3638 11936 3654 12000
rect 3718 11936 3734 12000
rect 3798 11936 3814 12000
rect 3878 11936 3886 12000
rect 3566 10912 3886 11936
rect 3566 10848 3574 10912
rect 3638 10848 3654 10912
rect 3718 10848 3734 10912
rect 3798 10848 3814 10912
rect 3878 10848 3886 10912
rect 3566 10134 3886 10848
rect 3566 9898 3608 10134
rect 3844 9898 3886 10134
rect 3566 9824 3886 9898
rect 3566 9760 3574 9824
rect 3638 9760 3654 9824
rect 3718 9760 3734 9824
rect 3798 9760 3814 9824
rect 3878 9760 3886 9824
rect 3566 8736 3886 9760
rect 3566 8672 3574 8736
rect 3638 8672 3654 8736
rect 3718 8672 3734 8736
rect 3798 8672 3814 8736
rect 3878 8672 3886 8736
rect 3566 7648 3886 8672
rect 3566 7584 3574 7648
rect 3638 7584 3654 7648
rect 3718 7584 3734 7648
rect 3798 7584 3814 7648
rect 3878 7584 3886 7648
rect 3566 6560 3886 7584
rect 3566 6496 3574 6560
rect 3638 6496 3654 6560
rect 3718 6496 3734 6560
rect 3798 6496 3814 6560
rect 3878 6496 3886 6560
rect 3566 5472 3886 6496
rect 3566 5408 3574 5472
rect 3638 5408 3654 5472
rect 3718 5408 3734 5472
rect 3798 5408 3814 5472
rect 3878 5408 3886 5472
rect 3566 4875 3886 5408
rect 3566 4639 3608 4875
rect 3844 4639 3886 4875
rect 3566 4384 3886 4639
rect 3566 4320 3574 4384
rect 3638 4320 3654 4384
rect 3718 4320 3734 4384
rect 3798 4320 3814 4384
rect 3878 4320 3886 4384
rect 3566 3296 3886 4320
rect 3566 3232 3574 3296
rect 3638 3232 3654 3296
rect 3718 3232 3734 3296
rect 3798 3232 3814 3296
rect 3878 3232 3886 3296
rect 3566 2208 3886 3232
rect 3566 2144 3574 2208
rect 3638 2144 3654 2208
rect 3718 2144 3734 2208
rect 3798 2144 3814 2208
rect 3878 2144 3886 2208
rect 3566 2128 3886 2144
rect 6188 17984 6508 18000
rect 6188 17920 6196 17984
rect 6260 17920 6276 17984
rect 6340 17920 6356 17984
rect 6420 17920 6436 17984
rect 6500 17920 6508 17984
rect 6188 16896 6508 17920
rect 6188 16832 6196 16896
rect 6260 16832 6276 16896
rect 6340 16832 6356 16896
rect 6420 16832 6436 16896
rect 6500 16832 6508 16896
rect 6188 15808 6508 16832
rect 6188 15744 6196 15808
rect 6260 15744 6276 15808
rect 6340 15744 6356 15808
rect 6420 15744 6436 15808
rect 6500 15744 6508 15808
rect 6188 14720 6508 15744
rect 6188 14656 6196 14720
rect 6260 14656 6276 14720
rect 6340 14656 6356 14720
rect 6420 14656 6436 14720
rect 6500 14656 6508 14720
rect 6188 13632 6508 14656
rect 6188 13568 6196 13632
rect 6260 13568 6276 13632
rect 6340 13568 6356 13632
rect 6420 13568 6436 13632
rect 6500 13568 6508 13632
rect 6188 12763 6508 13568
rect 6188 12544 6230 12763
rect 6466 12544 6508 12763
rect 6188 12480 6196 12544
rect 6260 12480 6276 12527
rect 6340 12480 6356 12527
rect 6420 12480 6436 12527
rect 6500 12480 6508 12544
rect 6188 11456 6508 12480
rect 6188 11392 6196 11456
rect 6260 11392 6276 11456
rect 6340 11392 6356 11456
rect 6420 11392 6436 11456
rect 6500 11392 6508 11456
rect 6188 10368 6508 11392
rect 6188 10304 6196 10368
rect 6260 10304 6276 10368
rect 6340 10304 6356 10368
rect 6420 10304 6436 10368
rect 6500 10304 6508 10368
rect 6188 9280 6508 10304
rect 6188 9216 6196 9280
rect 6260 9216 6276 9280
rect 6340 9216 6356 9280
rect 6420 9216 6436 9280
rect 6500 9216 6508 9280
rect 6188 8192 6508 9216
rect 6188 8128 6196 8192
rect 6260 8128 6276 8192
rect 6340 8128 6356 8192
rect 6420 8128 6436 8192
rect 6500 8128 6508 8192
rect 6188 7504 6508 8128
rect 6188 7268 6230 7504
rect 6466 7268 6508 7504
rect 6188 7104 6508 7268
rect 6188 7040 6196 7104
rect 6260 7040 6276 7104
rect 6340 7040 6356 7104
rect 6420 7040 6436 7104
rect 6500 7040 6508 7104
rect 6188 6016 6508 7040
rect 6188 5952 6196 6016
rect 6260 5952 6276 6016
rect 6340 5952 6356 6016
rect 6420 5952 6436 6016
rect 6500 5952 6508 6016
rect 6188 4928 6508 5952
rect 6188 4864 6196 4928
rect 6260 4864 6276 4928
rect 6340 4864 6356 4928
rect 6420 4864 6436 4928
rect 6500 4864 6508 4928
rect 6188 3840 6508 4864
rect 6188 3776 6196 3840
rect 6260 3776 6276 3840
rect 6340 3776 6356 3840
rect 6420 3776 6436 3840
rect 6500 3776 6508 3840
rect 6188 2752 6508 3776
rect 6188 2688 6196 2752
rect 6260 2688 6276 2752
rect 6340 2688 6356 2752
rect 6420 2688 6436 2752
rect 6500 2688 6508 2752
rect 6188 2128 6508 2688
rect 8810 17440 9130 18000
rect 8810 17376 8818 17440
rect 8882 17376 8898 17440
rect 8962 17376 8978 17440
rect 9042 17376 9058 17440
rect 9122 17376 9130 17440
rect 8810 16352 9130 17376
rect 8810 16288 8818 16352
rect 8882 16288 8898 16352
rect 8962 16288 8978 16352
rect 9042 16288 9058 16352
rect 9122 16288 9130 16352
rect 8810 15392 9130 16288
rect 8810 15264 8852 15392
rect 9088 15264 9130 15392
rect 8810 15200 8818 15264
rect 9122 15200 9130 15264
rect 8810 15156 8852 15200
rect 9088 15156 9130 15200
rect 8810 14176 9130 15156
rect 8810 14112 8818 14176
rect 8882 14112 8898 14176
rect 8962 14112 8978 14176
rect 9042 14112 9058 14176
rect 9122 14112 9130 14176
rect 8810 13088 9130 14112
rect 8810 13024 8818 13088
rect 8882 13024 8898 13088
rect 8962 13024 8978 13088
rect 9042 13024 9058 13088
rect 9122 13024 9130 13088
rect 8810 12000 9130 13024
rect 8810 11936 8818 12000
rect 8882 11936 8898 12000
rect 8962 11936 8978 12000
rect 9042 11936 9058 12000
rect 9122 11936 9130 12000
rect 8810 10912 9130 11936
rect 8810 10848 8818 10912
rect 8882 10848 8898 10912
rect 8962 10848 8978 10912
rect 9042 10848 9058 10912
rect 9122 10848 9130 10912
rect 8810 10134 9130 10848
rect 8810 9898 8852 10134
rect 9088 9898 9130 10134
rect 8810 9824 9130 9898
rect 8810 9760 8818 9824
rect 8882 9760 8898 9824
rect 8962 9760 8978 9824
rect 9042 9760 9058 9824
rect 9122 9760 9130 9824
rect 8810 8736 9130 9760
rect 8810 8672 8818 8736
rect 8882 8672 8898 8736
rect 8962 8672 8978 8736
rect 9042 8672 9058 8736
rect 9122 8672 9130 8736
rect 8810 7648 9130 8672
rect 8810 7584 8818 7648
rect 8882 7584 8898 7648
rect 8962 7584 8978 7648
rect 9042 7584 9058 7648
rect 9122 7584 9130 7648
rect 8810 6560 9130 7584
rect 8810 6496 8818 6560
rect 8882 6496 8898 6560
rect 8962 6496 8978 6560
rect 9042 6496 9058 6560
rect 9122 6496 9130 6560
rect 8810 5472 9130 6496
rect 8810 5408 8818 5472
rect 8882 5408 8898 5472
rect 8962 5408 8978 5472
rect 9042 5408 9058 5472
rect 9122 5408 9130 5472
rect 8810 4875 9130 5408
rect 8810 4639 8852 4875
rect 9088 4639 9130 4875
rect 8810 4384 9130 4639
rect 8810 4320 8818 4384
rect 8882 4320 8898 4384
rect 8962 4320 8978 4384
rect 9042 4320 9058 4384
rect 9122 4320 9130 4384
rect 8810 3296 9130 4320
rect 8810 3232 8818 3296
rect 8882 3232 8898 3296
rect 8962 3232 8978 3296
rect 9042 3232 9058 3296
rect 9122 3232 9130 3296
rect 8810 2208 9130 3232
rect 8810 2144 8818 2208
rect 8882 2144 8898 2208
rect 8962 2144 8978 2208
rect 9042 2144 9058 2208
rect 9122 2144 9130 2208
rect 8810 2128 9130 2144
rect 11432 17984 11752 18000
rect 11432 17920 11440 17984
rect 11504 17920 11520 17984
rect 11584 17920 11600 17984
rect 11664 17920 11680 17984
rect 11744 17920 11752 17984
rect 11432 16896 11752 17920
rect 11432 16832 11440 16896
rect 11504 16832 11520 16896
rect 11584 16832 11600 16896
rect 11664 16832 11680 16896
rect 11744 16832 11752 16896
rect 11432 15808 11752 16832
rect 11432 15744 11440 15808
rect 11504 15744 11520 15808
rect 11584 15744 11600 15808
rect 11664 15744 11680 15808
rect 11744 15744 11752 15808
rect 11432 14720 11752 15744
rect 11432 14656 11440 14720
rect 11504 14656 11520 14720
rect 11584 14656 11600 14720
rect 11664 14656 11680 14720
rect 11744 14656 11752 14720
rect 11432 13632 11752 14656
rect 11432 13568 11440 13632
rect 11504 13568 11520 13632
rect 11584 13568 11600 13632
rect 11664 13568 11680 13632
rect 11744 13568 11752 13632
rect 11432 12763 11752 13568
rect 11432 12544 11474 12763
rect 11710 12544 11752 12763
rect 11432 12480 11440 12544
rect 11504 12480 11520 12527
rect 11584 12480 11600 12527
rect 11664 12480 11680 12527
rect 11744 12480 11752 12544
rect 11432 11456 11752 12480
rect 11432 11392 11440 11456
rect 11504 11392 11520 11456
rect 11584 11392 11600 11456
rect 11664 11392 11680 11456
rect 11744 11392 11752 11456
rect 11432 10368 11752 11392
rect 11432 10304 11440 10368
rect 11504 10304 11520 10368
rect 11584 10304 11600 10368
rect 11664 10304 11680 10368
rect 11744 10304 11752 10368
rect 11432 9280 11752 10304
rect 11432 9216 11440 9280
rect 11504 9216 11520 9280
rect 11584 9216 11600 9280
rect 11664 9216 11680 9280
rect 11744 9216 11752 9280
rect 11432 8192 11752 9216
rect 11432 8128 11440 8192
rect 11504 8128 11520 8192
rect 11584 8128 11600 8192
rect 11664 8128 11680 8192
rect 11744 8128 11752 8192
rect 11432 7504 11752 8128
rect 11432 7268 11474 7504
rect 11710 7268 11752 7504
rect 11432 7104 11752 7268
rect 11432 7040 11440 7104
rect 11504 7040 11520 7104
rect 11584 7040 11600 7104
rect 11664 7040 11680 7104
rect 11744 7040 11752 7104
rect 11432 6016 11752 7040
rect 11432 5952 11440 6016
rect 11504 5952 11520 6016
rect 11584 5952 11600 6016
rect 11664 5952 11680 6016
rect 11744 5952 11752 6016
rect 11432 4928 11752 5952
rect 11432 4864 11440 4928
rect 11504 4864 11520 4928
rect 11584 4864 11600 4928
rect 11664 4864 11680 4928
rect 11744 4864 11752 4928
rect 11432 3840 11752 4864
rect 11432 3776 11440 3840
rect 11504 3776 11520 3840
rect 11584 3776 11600 3840
rect 11664 3776 11680 3840
rect 11744 3776 11752 3840
rect 11432 2752 11752 3776
rect 11432 2688 11440 2752
rect 11504 2688 11520 2752
rect 11584 2688 11600 2752
rect 11664 2688 11680 2752
rect 11744 2688 11752 2752
rect 11432 2128 11752 2688
rect 14054 17440 14374 18000
rect 14054 17376 14062 17440
rect 14126 17376 14142 17440
rect 14206 17376 14222 17440
rect 14286 17376 14302 17440
rect 14366 17376 14374 17440
rect 14054 16352 14374 17376
rect 14054 16288 14062 16352
rect 14126 16288 14142 16352
rect 14206 16288 14222 16352
rect 14286 16288 14302 16352
rect 14366 16288 14374 16352
rect 14054 15392 14374 16288
rect 14054 15264 14096 15392
rect 14332 15264 14374 15392
rect 14054 15200 14062 15264
rect 14366 15200 14374 15264
rect 14054 15156 14096 15200
rect 14332 15156 14374 15200
rect 14054 14176 14374 15156
rect 14054 14112 14062 14176
rect 14126 14112 14142 14176
rect 14206 14112 14222 14176
rect 14286 14112 14302 14176
rect 14366 14112 14374 14176
rect 14054 13088 14374 14112
rect 14054 13024 14062 13088
rect 14126 13024 14142 13088
rect 14206 13024 14222 13088
rect 14286 13024 14302 13088
rect 14366 13024 14374 13088
rect 14054 12000 14374 13024
rect 14054 11936 14062 12000
rect 14126 11936 14142 12000
rect 14206 11936 14222 12000
rect 14286 11936 14302 12000
rect 14366 11936 14374 12000
rect 14054 10912 14374 11936
rect 14054 10848 14062 10912
rect 14126 10848 14142 10912
rect 14206 10848 14222 10912
rect 14286 10848 14302 10912
rect 14366 10848 14374 10912
rect 14054 10134 14374 10848
rect 14054 9898 14096 10134
rect 14332 9898 14374 10134
rect 14054 9824 14374 9898
rect 14054 9760 14062 9824
rect 14126 9760 14142 9824
rect 14206 9760 14222 9824
rect 14286 9760 14302 9824
rect 14366 9760 14374 9824
rect 14054 8736 14374 9760
rect 14054 8672 14062 8736
rect 14126 8672 14142 8736
rect 14206 8672 14222 8736
rect 14286 8672 14302 8736
rect 14366 8672 14374 8736
rect 14054 7648 14374 8672
rect 14054 7584 14062 7648
rect 14126 7584 14142 7648
rect 14206 7584 14222 7648
rect 14286 7584 14302 7648
rect 14366 7584 14374 7648
rect 14054 6560 14374 7584
rect 14054 6496 14062 6560
rect 14126 6496 14142 6560
rect 14206 6496 14222 6560
rect 14286 6496 14302 6560
rect 14366 6496 14374 6560
rect 14054 5472 14374 6496
rect 14054 5408 14062 5472
rect 14126 5408 14142 5472
rect 14206 5408 14222 5472
rect 14286 5408 14302 5472
rect 14366 5408 14374 5472
rect 14054 4875 14374 5408
rect 14054 4639 14096 4875
rect 14332 4639 14374 4875
rect 14054 4384 14374 4639
rect 14054 4320 14062 4384
rect 14126 4320 14142 4384
rect 14206 4320 14222 4384
rect 14286 4320 14302 4384
rect 14366 4320 14374 4384
rect 14054 3296 14374 4320
rect 14054 3232 14062 3296
rect 14126 3232 14142 3296
rect 14206 3232 14222 3296
rect 14286 3232 14302 3296
rect 14366 3232 14374 3296
rect 14054 2208 14374 3232
rect 14054 2144 14062 2208
rect 14126 2144 14142 2208
rect 14206 2144 14222 2208
rect 14286 2144 14302 2208
rect 14366 2144 14374 2208
rect 14054 2128 14374 2144
<< via4 >>
rect 3608 15264 3844 15392
rect 3608 15200 3638 15264
rect 3638 15200 3654 15264
rect 3654 15200 3718 15264
rect 3718 15200 3734 15264
rect 3734 15200 3798 15264
rect 3798 15200 3814 15264
rect 3814 15200 3844 15264
rect 3608 15156 3844 15200
rect 3608 9898 3844 10134
rect 3608 4639 3844 4875
rect 6230 12544 6466 12763
rect 6230 12527 6260 12544
rect 6260 12527 6276 12544
rect 6276 12527 6340 12544
rect 6340 12527 6356 12544
rect 6356 12527 6420 12544
rect 6420 12527 6436 12544
rect 6436 12527 6466 12544
rect 6230 7268 6466 7504
rect 8852 15264 9088 15392
rect 8852 15200 8882 15264
rect 8882 15200 8898 15264
rect 8898 15200 8962 15264
rect 8962 15200 8978 15264
rect 8978 15200 9042 15264
rect 9042 15200 9058 15264
rect 9058 15200 9088 15264
rect 8852 15156 9088 15200
rect 8852 9898 9088 10134
rect 8852 4639 9088 4875
rect 11474 12544 11710 12763
rect 11474 12527 11504 12544
rect 11504 12527 11520 12544
rect 11520 12527 11584 12544
rect 11584 12527 11600 12544
rect 11600 12527 11664 12544
rect 11664 12527 11680 12544
rect 11680 12527 11710 12544
rect 11474 7268 11710 7504
rect 14096 15264 14332 15392
rect 14096 15200 14126 15264
rect 14126 15200 14142 15264
rect 14142 15200 14206 15264
rect 14206 15200 14222 15264
rect 14222 15200 14286 15264
rect 14286 15200 14302 15264
rect 14302 15200 14332 15264
rect 14096 15156 14332 15200
rect 14096 9898 14332 10134
rect 14096 4639 14332 4875
<< metal5 >>
rect 1104 15392 16836 15435
rect 1104 15156 3608 15392
rect 3844 15156 8852 15392
rect 9088 15156 14096 15392
rect 14332 15156 16836 15392
rect 1104 15114 16836 15156
rect 1104 12763 16836 12805
rect 1104 12527 6230 12763
rect 6466 12527 11474 12763
rect 11710 12527 16836 12763
rect 1104 12485 16836 12527
rect 1104 10134 16836 10176
rect 1104 9898 3608 10134
rect 3844 9898 8852 10134
rect 9088 9898 14096 10134
rect 14332 9898 16836 10134
rect 1104 9856 16836 9898
rect 1104 7504 16836 7547
rect 1104 7268 6230 7504
rect 6466 7268 11474 7504
rect 11710 7268 16836 7504
rect 1104 7226 16836 7268
rect 1104 4875 16836 4917
rect 1104 4639 3608 4875
rect 3844 4639 8852 4875
rect 9088 4639 14096 4875
rect 14332 4639 16836 4875
rect 1104 4597 16836 4639
use sky130_fd_sc_hd__dfrtp_4  _361_
timestamp 1623854003
transform 1 0 1380 0 1 2720
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1623854003
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1623854003
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1623854003
transform 1 0 1840 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1623854003
transform -1 0 1656 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6
timestamp 1623854003
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_11
timestamp 1623854003
transform 1 0 2116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23
timestamp 1623854003
transform 1 0 3220 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _184_
timestamp 1623854003
transform -1 0 4508 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _199_
timestamp 1623854003
transform -1 0 5060 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _200_
timestamp 1623854003
transform 1 0 5336 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _376_
timestamp 1623854003
transform 1 0 3496 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1623854003
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1623854003
transform 1 0 3496 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1623854003
transform 1 0 5060 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37
timestamp 1623854003
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46
timestamp 1623854003
transform 1 0 5336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1623854003
transform 1 0 5704 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1623854003
transform -1 0 6348 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1623854003
transform -1 0 6440 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53
timestamp 1623854003
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__a31o_1  _274_
timestamp 1623854003
transform 1 0 6808 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1623854003
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1623854003
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output36
timestamp 1623854003
transform 1 0 6624 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59
timestamp 1623854003
transform 1 0 6532 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_58
timestamp 1623854003
transform 1 0 6440 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _267_
timestamp 1623854003
transform -1 0 7452 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1623854003
transform 1 0 7452 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _273_
timestamp 1623854003
transform -1 0 7820 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1623854003
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _275_
timestamp 1623854003
transform 1 0 8372 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1623854003
transform 1 0 8280 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73
timestamp 1623854003
transform 1 0 7820 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77
timestamp 1623854003
transform 1 0 8188 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81
timestamp 1623854003
transform 1 0 8556 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_72
timestamp 1623854003
transform 1 0 7728 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_78
timestamp 1623854003
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1623854003
transform -1 0 10120 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _276_
timestamp 1623854003
transform 1 0 9200 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1623854003
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1623854003
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_93
timestamp 1623854003
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _360_
timestamp 1623854003
transform 1 0 9200 0 -1 2720
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_1  _321_
timestamp 1623854003
transform -1 0 10396 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1623854003
transform -1 0 10672 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_104
timestamp 1623854003
transform 1 0 10672 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _206_
timestamp 1623854003
transform 1 0 10948 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1623854003
transform -1 0 11776 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_111
timestamp 1623854003
transform 1 0 11316 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__o2bb2a_1  _194_
timestamp 1623854003
transform 1 0 11868 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _195_
timestamp 1623854003
transform 1 0 11684 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1623854003
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1623854003
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _185_
timestamp 1623854003
transform 1 0 12420 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _375_
timestamp 1623854003
transform -1 0 14444 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1623854003
transform -1 0 13616 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_122
timestamp 1623854003
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_130
timestamp 1623854003
transform 1 0 13064 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_136
timestamp 1623854003
transform 1 0 13616 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _306_
timestamp 1623854003
transform 1 0 14536 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1623854003
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1623854003
transform -1 0 15456 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_149
timestamp 1623854003
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _323_
timestamp 1623854003
transform -1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1623854003
transform 1 0 16284 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1623854003
transform 1 0 16008 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1623854003
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_160
timestamp 1623854003
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _358_
timestamp 1623854003
transform 1 0 14720 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1623854003
transform -1 0 16836 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1623854003
transform -1 0 16836 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _305_
timestamp 1623854003
transform -1 0 3404 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 1623854003
transform -1 0 2576 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1623854003
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1623854003
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6
timestamp 1623854003
transform 1 0 1656 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_12
timestamp 1623854003
transform 1 0 2208 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_16
timestamp 1623854003
transform 1 0 2576 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _192_
timestamp 1623854003
transform 1 0 5152 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _197_
timestamp 1623854003
transform 1 0 4416 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1623854003
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_25
timestamp 1623854003
transform 1 0 3404 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_30
timestamp 1623854003
transform 1 0 3864 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_47
timestamp 1623854003
transform 1 0 5428 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _272_
timestamp 1623854003
transform 1 0 6900 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_59
timestamp 1623854003
transform 1 0 6532 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_70
timestamp 1623854003
transform 1 0 7544 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1623854003
transform -1 0 8648 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1623854003
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_78
timestamp 1623854003
transform 1 0 8280 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_82
timestamp 1623854003
transform 1 0 8648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_87
timestamp 1623854003
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _193_
timestamp 1623854003
transform 1 0 11960 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _208_
timestamp 1623854003
transform 1 0 10764 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_2_99
timestamp 1623854003
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1623854003
transform -1 0 13064 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1623854003
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_130
timestamp 1623854003
transform 1 0 13064 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_142
timestamp 1623854003
transform 1 0 14168 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _178_
timestamp 1623854003
transform -1 0 16560 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_2_144
timestamp 1623854003
transform 1 0 14352 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1623854003
transform -1 0 16836 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1623854003
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1623854003
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1623854003
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__a22oi_2  _201_
timestamp 1623854003
transform -1 0 5796 0 1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1623854003
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_39
timestamp 1623854003
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__a311o_1  _277_
timestamp 1623854003
transform -1 0 7360 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _359_
timestamp 1623854003
transform 1 0 7360 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1623854003
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1623854003
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_58
timestamp 1623854003
transform 1 0 6440 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_88
timestamp 1623854003
transform 1 0 9200 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _186_
timestamp 1623854003
transform 1 0 12052 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _209_
timestamp 1623854003
transform 1 0 11224 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1623854003
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_100
timestamp 1623854003
transform 1 0 10304 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_108
timestamp 1623854003
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1623854003
transform 1 0 11500 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1623854003
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _374_
timestamp 1623854003
transform 1 0 12696 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _357_
timestamp 1623854003
transform 1 0 14536 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1623854003
transform 1 0 16376 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1623854003
transform -1 0 16836 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1623854003
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1623854003
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1623854003
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_1  _198_
timestamp 1623854003
transform -1 0 4692 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _204_
timestamp 1623854003
transform -1 0 5980 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1623854003
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1623854003
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1623854003
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_39
timestamp 1623854003
transform 1 0 4692 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _202_
timestamp 1623854003
transform 1 0 5980 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_4_58
timestamp 1623854003
transform 1 0 6440 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_70
timestamp 1623854003
transform 1 0 7544 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1623854003
transform 1 0 9568 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _216_
timestamp 1623854003
transform 1 0 9108 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1623854003
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_82
timestamp 1623854003
transform 1 0 8648 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_95
timestamp 1623854003
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _210_
timestamp 1623854003
transform -1 0 12788 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o2111ai_4  _225_
timestamp 1623854003
transform 1 0 10028 0 -1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _307_
timestamp 1623854003
transform 1 0 13800 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1623854003
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_127
timestamp 1623854003
transform 1 0 12788 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_135
timestamp 1623854003
transform 1 0 13524 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1623854003
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp 1623854003
transform -1 0 15732 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1623854003
transform -1 0 16560 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144
timestamp 1623854003
transform 1 0 14352 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_159
timestamp 1623854003
transform 1 0 15732 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1623854003
transform -1 0 16836 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _377_
timestamp 1623854003
transform 1 0 1564 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1623854003
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1623854003
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_1  _191_
timestamp 1623854003
transform 1 0 4508 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _213_
timestamp 1623854003
transform -1 0 4508 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_25
timestamp 1623854003
transform 1 0 3404 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_43
timestamp 1623854003
transform 1 0 5060 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _269_
timestamp 1623854003
transform -1 0 7544 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _271_
timestamp 1623854003
transform -1 0 7268 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _319_
timestamp 1623854003
transform -1 0 6348 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1623854003
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_51
timestamp 1623854003
transform 1 0 5796 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_70
timestamp 1623854003
transform 1 0 7544 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _214_
timestamp 1623854003
transform 1 0 8832 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _215_
timestamp 1623854003
transform -1 0 8832 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _217_
timestamp 1623854003
transform -1 0 10304 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_89
timestamp 1623854003
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1623854003
transform -1 0 11960 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _205_
timestamp 1623854003
transform -1 0 10580 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _207_
timestamp 1623854003
transform 1 0 11960 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _211_
timestamp 1623854003
transform 1 0 11224 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1623854003
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_103
timestamp 1623854003
transform 1 0 10580 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_109
timestamp 1623854003
transform 1 0 11132 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _316_
timestamp 1623854003
transform -1 0 13248 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_121
timestamp 1623854003
transform 1 0 12236 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_132
timestamp 1623854003
transform 1 0 13248 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_144
timestamp 1623854003
transform 1 0 14352 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_156
timestamp 1623854003
transform 1 0 15456 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1623854003
transform -1 0 16836 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1623854003
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1623854003
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1623854003
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1623854003
transform 1 0 1380 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp 1623854003
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _183_
timestamp 1623854003
transform -1 0 3772 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp 1623854003
transform -1 0 2576 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_18
timestamp 1623854003
transform 1 0 2760 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_6
timestamp 1623854003
transform 1 0 1656 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_16
timestamp 1623854003
transform 1 0 2576 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_4  _179_
timestamp 1623854003
transform 1 0 5060 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _190_
timestamp 1623854003
transform -1 0 4232 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1623854003
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_30
timestamp 1623854003
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_34
timestamp 1623854003
transform 1 0 4232 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_46
timestamp 1623854003
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_28
timestamp 1623854003
transform 1 0 3680 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_40
timestamp 1623854003
transform 1 0 4784 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1623854003
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _362_
timestamp 1623854003
transform -1 0 7452 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1623854003
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_69
timestamp 1623854003
transform 1 0 7452 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1623854003
transform 1 0 5704 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_56
timestamp 1623854003
transform 1 0 6256 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_58
timestamp 1623854003
transform 1 0 6440 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_65
timestamp 1623854003
transform 1 0 7084 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1623854003
transform 1 0 8740 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _212_
timestamp 1623854003
transform -1 0 8648 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_6_81
timestamp 1623854003
transform 1 0 8556 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_73
timestamp 1623854003
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_82
timestamp 1623854003
transform 1 0 8648 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1623854003
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1623854003
transform 1 0 8924 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_86
timestamp 1623854003
transform 1 0 9016 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_94
timestamp 1623854003
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__o221ai_2  _218_
timestamp 1623854003
transform -1 0 10212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _219_
timestamp 1623854003
transform 1 0 10764 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _233_
timestamp 1623854003
transform -1 0 12144 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _234_
timestamp 1623854003
transform 1 0 9936 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _365_
timestamp 1623854003
transform 1 0 11960 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1623854003
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_99
timestamp 1623854003
transform 1 0 10212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_111
timestamp 1623854003
transform 1 0 11316 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_117
timestamp 1623854003
transform 1 0 11868 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_112
timestamp 1623854003
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1623854003
transform -1 0 13524 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _364_
timestamp 1623854003
transform 1 0 13524 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1623854003
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_138
timestamp 1623854003
transform 1 0 13800 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_142
timestamp 1623854003
transform 1 0 14168 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_120
timestamp 1623854003
transform 1 0 12144 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _317_
timestamp 1623854003
transform -1 0 14720 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _325_
timestamp 1623854003
transform -1 0 16008 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _356_
timestamp 1623854003
transform -1 0 16560 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1623854003
transform 1 0 16284 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_144
timestamp 1623854003
transform 1 0 14352 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_155
timestamp 1623854003
transform 1 0 15364 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_162
timestamp 1623854003
transform 1 0 16008 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1623854003
transform -1 0 16836 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1623854003
transform -1 0 16836 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _372_
timestamp 1623854003
transform 1 0 1472 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1623854003
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1623854003
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _373_
timestamp 1623854003
transform 1 0 3956 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1623854003
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1623854003
transform 1 0 3312 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_28
timestamp 1623854003
transform 1 0 3680 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1623854003
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_1  _270_
timestamp 1623854003
transform 1 0 6256 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_51
timestamp 1623854003
transform 1 0 5796 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_55
timestamp 1623854003
transform 1 0 6164 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_60
timestamp 1623854003
transform 1 0 6624 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _180_
timestamp 1623854003
transform 1 0 7728 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1623854003
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_79
timestamp 1623854003
transform 1 0 8372 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1623854003
transform 1 0 8924 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1623854003
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1623854003
transform 1 0 10396 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _264_
timestamp 1623854003
transform 1 0 11776 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o22ai_1  _265_
timestamp 1623854003
transform 1 0 11316 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_8_99
timestamp 1623854003
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_104
timestamp 1623854003
transform 1 0 10672 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_110
timestamp 1623854003
transform 1 0 11224 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1623854003
transform -1 0 12788 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _266_
timestamp 1623854003
transform 1 0 13524 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1623854003
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_127
timestamp 1623854003
transform 1 0 12788 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_142
timestamp 1623854003
transform 1 0 14168 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1623854003
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_156
timestamp 1623854003
transform 1 0 15456 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1623854003
transform -1 0 16836 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _188_
timestamp 1623854003
transform -1 0 3864 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _371_
timestamp 1623854003
transform 1 0 1380 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1623854003
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _187_
timestamp 1623854003
transform -1 0 4508 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _226_
timestamp 1623854003
transform 1 0 4508 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _308_
timestamp 1623854003
transform 1 0 5152 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1623854003
transform 1 0 5428 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _363_
timestamp 1623854003
transform 1 0 6440 0 1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1623854003
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_55
timestamp 1623854003
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _378_
timestamp 1623854003
transform -1 0 10212 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__o31a_4  _235_
timestamp 1623854003
transform 1 0 10212 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _237_
timestamp 1623854003
transform -1 0 12512 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1623854003
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1623854003
transform 1 0 11500 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_115
timestamp 1623854003
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__or3_1  _224_
timestamp 1623854003
transform 1 0 12512 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _249_
timestamp 1623854003
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _250_
timestamp 1623854003
transform -1 0 14628 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_129
timestamp 1623854003
transform 1 0 12972 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_2  _370_
timestamp 1623854003
transform 1 0 14628 0 1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1623854003
transform -1 0 16836 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _189_
timestamp 1623854003
transform -1 0 3220 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp 1623854003
transform -1 0 2576 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1623854003
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1623854003
transform -1 0 1656 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_6
timestamp 1623854003
transform 1 0 1656 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_12
timestamp 1623854003
transform 1 0 2208 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_16
timestamp 1623854003
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_23
timestamp 1623854003
transform 1 0 3220 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1623854003
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1623854003
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1623854003
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1623854003
transform -1 0 6900 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_54
timestamp 1623854003
transform 1 0 6072 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_63
timestamp 1623854003
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1623854003
transform 1 0 9108 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1623854003
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_75
timestamp 1623854003
transform 1 0 8004 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_83
timestamp 1623854003
transform 1 0 8740 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_90
timestamp 1623854003
transform 1 0 9384 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _238_
timestamp 1623854003
transform 1 0 11592 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_10_102
timestamp 1623854003
transform 1 0 10488 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _247_
timestamp 1623854003
transform -1 0 14168 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1623854003
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1623854003
transform 1 0 12236 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_133
timestamp 1623854003
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_142
timestamp 1623854003
transform 1 0 14168 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1623854003
transform 1 0 14352 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1623854003
transform 1 0 14628 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _311_
timestamp 1623854003
transform -1 0 15916 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_150
timestamp 1623854003
transform 1 0 14904 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_161
timestamp 1623854003
transform 1 0 15916 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1623854003
transform -1 0 16836 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_167
timestamp 1623854003
transform 1 0 16468 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1623854003
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1623854003
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1623854003
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1623854003
transform 1 0 4784 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1623854003
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_39
timestamp 1623854003
transform 1 0 4692 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_43
timestamp 1623854003
transform 1 0 5060 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__o2bb2a_1  _261_
timestamp 1623854003
transform 1 0 6808 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1623854003
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_55
timestamp 1623854003
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_58
timestamp 1623854003
transform 1 0 6440 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_70
timestamp 1623854003
transform 1 0 7544 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _315_
timestamp 1623854003
transform 1 0 8464 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_78
timestamp 1623854003
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_83
timestamp 1623854003
transform 1 0 8740 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_95
timestamp 1623854003
transform 1 0 9844 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _259_
timestamp 1623854003
transform 1 0 9936 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1623854003
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_105
timestamp 1623854003
transform 1 0 10764 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1623854003
transform 1 0 11500 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_115
timestamp 1623854003
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1623854003
transform 1 0 13892 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_127
timestamp 1623854003
transform 1 0 12788 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_142
timestamp 1623854003
transform 1 0 14168 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1623854003
transform 1 0 16284 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_154
timestamp 1623854003
transform 1 0 15272 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_162
timestamp 1623854003
transform 1 0 16008 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1623854003
transform -1 0 16836 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _349_
timestamp 1623854003
transform -1 0 3680 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01
timestamp 1623854003
transform -1 0 2576 0 -1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1623854003
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_16
timestamp 1623854003
transform 1 0 2576 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1623854003
transform 1 0 4508 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp 1623854003
transform -1 0 5612 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb1
timestamp 1623854003
transform 1 0 3864 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1623854003
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_28
timestamp 1623854003
transform 1 0 3680 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_40
timestamp 1623854003
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _314_
timestamp 1623854003
transform -1 0 7084 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _348_
timestamp 1623854003
transform 1 0 5796 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _366_
timestamp 1623854003
transform 1 0 7084 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_12_49
timestamp 1623854003
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_60
timestamp 1623854003
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1623854003
transform 1 0 9384 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _260_
timestamp 1623854003
transform 1 0 9660 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1623854003
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_87
timestamp 1623854003
transform 1 0 9108 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _258_
timestamp 1623854003
transform -1 0 11592 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _262_
timestamp 1623854003
transform -1 0 11868 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _263_
timestamp 1623854003
transform 1 0 10396 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_117
timestamp 1623854003
transform 1 0 11868 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _256_
timestamp 1623854003
transform -1 0 13432 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _257_
timestamp 1623854003
transform -1 0 13156 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1623854003
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_134
timestamp 1623854003
transform 1 0 13432 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_142
timestamp 1623854003
transform 1 0 14168 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _368_
timestamp 1623854003
transform 1 0 14628 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_12_144
timestamp 1623854003
transform 1 0 14352 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1623854003
transform -1 0 16836 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_8  _182_
timestamp 1623854003
transform -1 0 3404 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00
timestamp 1623854003
transform -1 0 2300 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1
timestamp 1623854003
transform -1 0 2576 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1623854003
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1623854003
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1623854003
transform -1 0 1656 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1623854003
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_16
timestamp 1623854003
transform 1 0 2576 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_6
timestamp 1623854003
transform 1 0 1656 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1623854003
transform -1 0 5520 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen1
timestamp 1623854003
transform 1 0 3496 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb0
timestamp 1623854003
transform -1 0 5152 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1623854003
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_24
timestamp 1623854003
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_31
timestamp 1623854003
transform 1 0 3956 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_25
timestamp 1623854003
transform 1 0 3404 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1623854003
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1623854003
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _367_
timestamp 1623854003
transform 1 0 6440 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1623854003
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_48
timestamp 1623854003
transform 1 0 5520 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_56
timestamp 1623854003
transform 1 0 6256 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_54
timestamp 1623854003
transform 1 0 6072 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_66
timestamp 1623854003
transform 1 0 7176 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1623854003
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_79
timestamp 1623854003
transform 1 0 8372 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_91
timestamp 1623854003
transform 1 0 9476 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_78
timestamp 1623854003
transform 1 0 8280 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_87
timestamp 1623854003
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _240_
timestamp 1623854003
transform 1 0 10028 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _241_
timestamp 1623854003
transform -1 0 11592 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _242_
timestamp 1623854003
transform 1 0 11960 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1623854003
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_104
timestamp 1623854003
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_115
timestamp 1623854003
transform 1 0 11684 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_99
timestamp 1623854003
transform 1 0 10212 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_111
timestamp 1623854003
transform 1 0 11316 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _243_
timestamp 1623854003
transform -1 0 14076 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _245_
timestamp 1623854003
transform -1 0 13800 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _251_
timestamp 1623854003
transform -1 0 13064 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _252_
timestamp 1623854003
transform 1 0 12420 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _254_
timestamp 1623854003
transform 1 0 13800 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1623854003
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_127
timestamp 1623854003
transform 1 0 12788 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_133
timestamp 1623854003
transform 1 0 13340 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1623854003
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1623854003
transform 1 0 14536 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1623854003
transform 1 0 14352 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _313_
timestamp 1623854003
transform -1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _369_
timestamp 1623854003
transform 1 0 14628 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_13_149
timestamp 1623854003
transform 1 0 14812 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1623854003
transform 1 0 15824 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1623854003
transform -1 0 16836 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1623854003
transform -1 0 16836 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1623854003
transform -1 0 3772 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.reseten0
timestamp 1623854003
transform 1 0 1932 0 1 10336
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1623854003
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1623854003
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen0
timestamp 1623854003
transform 1 0 4416 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb0
timestamp 1623854003
transform 1 0 3772 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1623854003
transform -1 0 5152 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_44
timestamp 1623854003
transform 1 0 5152 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _287_
timestamp 1623854003
transform 1 0 6440 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _289_
timestamp 1623854003
transform 1 0 5704 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _345_
timestamp 1623854003
transform 1 0 7268 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1623854003
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__o41a_2  _296_
timestamp 1623854003
transform 1 0 8832 0 1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _297_
timestamp 1623854003
transform -1 0 10580 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _298_
timestamp 1623854003
transform 1 0 8096 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1623854003
transform -1 0 11500 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _227_
timestamp 1623854003
transform 1 0 10580 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _239_
timestamp 1623854003
transform 1 0 11684 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _280_
timestamp 1623854003
transform -1 0 12696 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1623854003
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1623854003
transform 1 0 11500 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_118
timestamp 1623854003
transform 1 0 11960 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1623854003
transform -1 0 12972 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _255_
timestamp 1623854003
transform 1 0 14168 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_129
timestamp 1623854003
transform 1 0 12972 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_141
timestamp 1623854003
transform 1 0 14076 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp 1623854003
transform -1 0 15916 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_146
timestamp 1623854003
transform 1 0 14536 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1623854003
transform 1 0 15916 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1623854003
transform -1 0 16836 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1623854003
transform 1 0 16468 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _181_
timestamp 1623854003
transform 1 0 1564 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _330_
timestamp 1623854003
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1623854003
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1623854003
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_23
timestamp 1623854003
transform 1 0 3220 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen1
timestamp 1623854003
transform 1 0 5152 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb1
timestamp 1623854003
transform -1 0 5152 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1623854003
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_30
timestamp 1623854003
transform 1 0 3864 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_36
timestamp 1623854003
transform 1 0 4416 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1623854003
transform 1 0 7360 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1623854003
transform 1 0 5612 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_52
timestamp 1623854003
transform 1 0 5888 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_64
timestamp 1623854003
transform 1 0 6992 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _300_
timestamp 1623854003
transform 1 0 8188 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1623854003
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_87
timestamp 1623854003
transform 1 0 9108 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_95
timestamp 1623854003
transform 1 0 9844 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1623854003
transform 1 0 9936 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _221_
timestamp 1623854003
transform 1 0 10304 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _223_
timestamp 1623854003
transform 1 0 11408 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1623854003
transform 1 0 11132 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_99
timestamp 1623854003
transform 1 0 10212 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_105
timestamp 1623854003
transform 1 0 10764 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1623854003
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1623854003
transform 1 0 13984 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1623854003
transform 1 0 13156 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1623854003
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_129
timestamp 1623854003
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_134
timestamp 1623854003
transform 1 0 13432 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _301_
timestamp 1623854003
transform 1 0 14352 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _343_
timestamp 1623854003
transform 1 0 14812 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1623854003
transform 1 0 16284 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_147
timestamp 1623854003
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_158
timestamp 1623854003
transform 1 0 15640 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_164
timestamp 1623854003
transform 1 0 16192 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1623854003
transform -1 0 16836 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb0
timestamp 1623854003
transform 1 0 1564 0 1 11424
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1623854003
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1623854003
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_16
timestamp 1623854003
transform 1 0 2576 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1623854003
transform 1 0 4876 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_28
timestamp 1623854003
transform 1 0 3680 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_40
timestamp 1623854003
transform 1 0 4784 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_45
timestamp 1623854003
transform 1 0 5244 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__o31a_1  _303_
timestamp 1623854003
transform -1 0 7084 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1623854003
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_65
timestamp 1623854003
transform 1 0 7084 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_2  _294_
timestamp 1623854003
transform -1 0 10120 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _295_
timestamp 1623854003
transform 1 0 8832 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_77
timestamp 1623854003
transform 1 0 8188 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_83
timestamp 1623854003
transform 1 0 8740 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o31a_1  _281_
timestamp 1623854003
transform -1 0 12604 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1623854003
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1623854003
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_110
timestamp 1623854003
transform 1 0 11224 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_115
timestamp 1623854003
transform 1 0 11684 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _285_
timestamp 1623854003
transform 1 0 12604 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _336_
timestamp 1623854003
transform 1 0 13708 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_134
timestamp 1623854003
transform 1 0 13432 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _170_
timestamp 1623854003
transform 1 0 14536 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _339_
timestamp 1623854003
transform 1 0 15364 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_153
timestamp 1623854003
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1623854003
transform 1 0 16192 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1623854003
transform -1 0 16836 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0
timestamp 1623854003
transform -1 0 2116 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1623854003
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1623854003
transform -1 0 1656 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_11
timestamp 1623854003
transform 1 0 2116 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_23
timestamp 1623854003
transform 1 0 3220 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1623854003
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1623854003
transform 1 0 3864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_42
timestamp 1623854003
transform 1 0 4968 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _229_
timestamp 1623854003
transform 1 0 6808 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _284_
timestamp 1623854003
transform -1 0 6624 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _286_
timestamp 1623854003
transform -1 0 8372 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_60
timestamp 1623854003
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_69
timestamp 1623854003
transform 1 0 7452 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o311a_1  _293_
timestamp 1623854003
transform 1 0 9844 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1623854003
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_79
timestamp 1623854003
transform 1 0 8372 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1623854003
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_87
timestamp 1623854003
transform 1 0 9108 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _231_
timestamp 1623854003
transform -1 0 11776 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _292_
timestamp 1623854003
transform 1 0 11776 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _304_
timestamp 1623854003
transform 1 0 10580 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_119
timestamp 1623854003
transform 1 0 12052 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _278_
timestamp 1623854003
transform -1 0 13064 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1623854003
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_130
timestamp 1623854003
transform 1 0 13064 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_142
timestamp 1623854003
transform 1 0 14168 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _290_
timestamp 1623854003
transform 1 0 15456 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_18_144
timestamp 1623854003
transform 1 0 14352 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1623854003
transform 1 0 16100 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1623854003
transform -1 0 16836 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_167
timestamp 1623854003
transform 1 0 16468 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.iss.delayenb1
timestamp 1623854003
transform 1 0 1840 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1623854003
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1623854003
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1623854003
transform 1 0 1380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1623854003
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1623854003
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1623854003
transform 1 0 1748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1623854003
transform 1 0 2944 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.delayen0
timestamp 1623854003
transform 1 0 2300 0 1 12512
box -38 -48 1050 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.delayen1
timestamp 1623854003
transform 1 0 2484 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1623854003
transform 1 0 3220 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0
timestamp 1623854003
transform 1 0 3312 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb0
timestamp 1623854003
transform -1 0 4416 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb1
timestamp 1623854003
transform -1 0 4508 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1623854003
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_28
timestamp 1623854003
transform 1 0 3680 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_26
timestamp 1623854003
transform 1 0 3496 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1623854003
transform 1 0 5336 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1623854003
transform 1 0 4968 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen0
timestamp 1623854003
transform 1 0 4416 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen1
timestamp 1623854003
transform 1 0 4508 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_20_45
timestamp 1623854003
transform 1 0 5244 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_41
timestamp 1623854003
transform 1 0 4876 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _291_
timestamp 1623854003
transform 1 0 6440 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _302_
timestamp 1623854003
transform -1 0 7544 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _344_
timestamp 1623854003
transform 1 0 7544 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1623854003
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_53
timestamp 1623854003
transform 1 0 5980 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_55
timestamp 1623854003
transform 1 0 6164 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_67
timestamp 1623854003
transform 1 0 7268 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _337_
timestamp 1623854003
transform -1 0 10212 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1623854003
transform 1 0 8188 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1623854003
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  repeater38
timestamp 1623854003
transform -1 0 10856 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_79
timestamp 1623854003
transform 1 0 8372 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_91
timestamp 1623854003
transform 1 0 9476 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_75
timestamp 1623854003
transform 1 0 8004 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_87
timestamp 1623854003
transform 1 0 9108 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _232_
timestamp 1623854003
transform 1 0 10856 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _329_
timestamp 1623854003
transform 1 0 11684 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _347_
timestamp 1623854003
transform 1 0 11776 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _355_
timestamp 1623854003
transform 1 0 10212 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1623854003
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_111
timestamp 1623854003
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_108
timestamp 1623854003
transform 1 0 11040 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen1
timestamp 1623854003
transform 1 0 14076 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb1
timestamp 1623854003
transform 1 0 13432 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1623854003
transform 1 0 13984 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1623854003
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_124
timestamp 1623854003
transform 1 0 12512 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1623854003
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_125
timestamp 1623854003
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1623854003
transform 1 0 13708 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _338_
timestamp 1623854003
transform 1 0 15364 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1623854003
transform 1 0 14536 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_149
timestamp 1623854003
transform 1 0 14812 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1623854003
transform 1 0 16192 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1623854003
transform 1 0 14352 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_156
timestamp 1623854003
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1623854003
transform -1 0 16836 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1623854003
transform -1 0 16836 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1623854003
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1623854003
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1623854003
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 1623854003
transform 1 0 4692 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1623854003
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_42
timestamp 1623854003
transform 1 0 4968 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1623854003
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb1
timestamp 1623854003
transform 1 0 7268 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1623854003
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_50
timestamp 1623854003
transform 1 0 5704 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_58
timestamp 1623854003
transform 1 0 6440 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_66
timestamp 1623854003
transform 1 0 7176 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1623854003
transform 1 0 8372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen1
timestamp 1623854003
transform 1 0 7912 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_21_82
timestamp 1623854003
transform 1 0 8648 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_94
timestamp 1623854003
transform 1 0 9752 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _299_
timestamp 1623854003
transform 1 0 11684 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1623854003
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_106
timestamp 1623854003
transform 1 0 10856 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen0
timestamp 1623854003
transform 1 0 13708 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb0
timestamp 1623854003
transform 1 0 13064 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_21_120
timestamp 1623854003
transform 1 0 12144 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_128
timestamp 1623854003
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_142
timestamp 1623854003
transform 1 0 14168 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen0
timestamp 1623854003
transform 1 0 15548 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb0
timestamp 1623854003
transform -1 0 15548 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1623854003
transform -1 0 16376 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1623854003
transform 1 0 16376 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1623854003
transform -1 0 16836 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_4  ringosc.dstage\[11\].id.delayen0
timestamp 1623854003
transform 1 0 1840 0 -1 14688
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1623854003
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1623854003
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1623854003
transform 1 0 1748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 1623854003
transform 1 0 2852 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _354_
timestamp 1623854003
transform 1 0 3864 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1623854003
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1623854003
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_39
timestamp 1623854003
transform 1 0 4692 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_47
timestamp 1623854003
transform 1 0 5428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _282_
timestamp 1623854003
transform 1 0 5704 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _283_
timestamp 1623854003
transform 1 0 6348 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb0
timestamp 1623854003
transform 1 0 7452 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_22_64
timestamp 1623854003
transform 1 0 6992 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_68
timestamp 1623854003
transform 1 0 7360 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb0
timestamp 1623854003
transform -1 0 9844 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen0
timestamp 1623854003
transform 1 0 8096 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1623854003
transform 1 0 8556 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1623854003
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1623854003
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_87
timestamp 1623854003
transform 1 0 9108 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_95
timestamp 1623854003
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen0
timestamp 1623854003
transform 1 0 10028 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen1
timestamp 1623854003
transform 1 0 11868 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb1
timestamp 1623854003
transform -1 0 11868 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1623854003
transform -1 0 10856 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_106
timestamp 1623854003
transform 1 0 10856 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1623854003
transform 1 0 12328 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1623854003
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1623854003
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_137
timestamp 1623854003
transform 1 0 13708 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1623854003
transform 1 0 16284 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_144
timestamp 1623854003
transform 1 0 14352 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_156
timestamp 1623854003
transform 1 0 15456 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_164
timestamp 1623854003
transform 1 0 16192 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1623854003
transform -1 0 16836 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb0
timestamp 1623854003
transform 1 0 1472 0 1 14688
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1623854003
transform 1 0 2484 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1623854003
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1623854003
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_18
timestamp 1623854003
transform 1 0 2760 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _288_
timestamp 1623854003
transform -1 0 5888 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _332_
timestamp 1623854003
transform 1 0 3956 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_30
timestamp 1623854003
transform 1 0 3864 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_40
timestamp 1623854003
transform 1 0 4784 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_46
timestamp 1623854003
transform 1 0 5336 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _279_
timestamp 1623854003
transform 1 0 5888 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _340_
timestamp 1623854003
transform -1 0 7268 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1623854003
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_67
timestamp 1623854003
transform 1 0 7268 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_79
timestamp 1623854003
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_91
timestamp 1623854003
transform 1 0 9476 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _346_
timestamp 1623854003
transform 1 0 11684 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1623854003
transform -1 0 11592 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1623854003
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_103
timestamp 1623854003
transform 1 0 10580 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1623854003
transform 1 0 13892 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_124
timestamp 1623854003
transform 1 0 12512 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_136
timestamp 1623854003
transform 1 0 13616 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_143
timestamp 1623854003
transform 1 0 14260 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1623854003
transform 1 0 16192 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen1
timestamp 1623854003
transform 1 0 15732 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb1
timestamp 1623854003
transform 1 0 15088 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_23_151
timestamp 1623854003
transform 1 0 14996 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1623854003
transform -1 0 16836 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1623854003
transform 1 0 16468 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1623854003
transform -1 0 3404 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[11\].id.delayen1
timestamp 1623854003
transform 1 0 2392 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[11\].id.delayenb1
timestamp 1623854003
transform 1 0 1748 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1623854003
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1623854003
transform -1 0 1656 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_6
timestamp 1623854003
transform 1 0 1656 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_19
timestamp 1623854003
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1623854003
transform 1 0 3404 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1623854003
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_28
timestamp 1623854003
transform 1 0 3680 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1623854003
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_42
timestamp 1623854003
transform 1 0 4968 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_54
timestamp 1623854003
transform 1 0 6072 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_66
timestamp 1623854003
transform 1 0 7176 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1623854003
transform 1 0 8464 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1623854003
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_78
timestamp 1623854003
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1623854003
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_87
timestamp 1623854003
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1623854003
transform 1 0 11592 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_99
timestamp 1623854003
transform 1 0 10212 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_111
timestamp 1623854003
transform 1 0 11316 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_118
timestamp 1623854003
transform 1 0 11960 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _335_
timestamp 1623854003
transform -1 0 13800 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen1
timestamp 1623854003
transform 1 0 13800 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1623854003
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_126
timestamp 1623854003
transform 1 0 12696 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1623854003
transform 1 0 15732 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1623854003
transform 1 0 14352 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1623854003
transform 1 0 16284 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_147
timestamp 1623854003
transform 1 0 14628 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_162
timestamp 1623854003
transform 1 0 16008 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1623854003
transform -1 0 16836 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _331_
timestamp 1623854003
transform 1 0 1748 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1623854003
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1623854003
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_16
timestamp 1623854003
transform 1 0 2576 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen0
timestamp 1623854003
transform 1 0 4416 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb0
timestamp 1623854003
transform 1 0 3772 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_25_28
timestamp 1623854003
transform 1 0 3680 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_41
timestamp 1623854003
transform 1 0 4876 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1623854003
transform 1 0 5612 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[5\].id.delayenb1
timestamp 1623854003
transform 1 0 7636 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1623854003
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1623854003
transform 1 0 5888 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_56
timestamp 1623854003
transform 1 0 6256 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_58
timestamp 1623854003
transform 1 0 6440 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_70
timestamp 1623854003
transform 1 0 7544 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1623854003
transform 1 0 8740 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[5\].id.delayen1
timestamp 1623854003
transform 1 0 8280 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb0
timestamp 1623854003
transform 1 0 9476 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_25_86
timestamp 1623854003
transform 1 0 9016 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_90
timestamp 1623854003
transform 1 0 9384 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen0
timestamp 1623854003
transform 1 0 10120 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1623854003
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_103
timestamp 1623854003
transform 1 0 10580 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_111
timestamp 1623854003
transform 1 0 11316 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1623854003
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb1
timestamp 1623854003
transform 1 0 13064 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1623854003
transform 1 0 13708 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_127
timestamp 1623854003
transform 1 0 12788 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_140
timestamp 1623854003
transform 1 0 13984 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_152
timestamp 1623854003
transform 1 0 15088 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1623854003
transform 1 0 16192 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1623854003
transform -1 0 16836 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1623854003
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1623854003
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1623854003
transform -1 0 1656 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1623854003
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1623854003
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_6
timestamp 1623854003
transform 1 0 1656 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_18
timestamp 1623854003
transform 1 0 2760 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _333_
timestamp 1623854003
transform -1 0 4508 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1623854003
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1623854003
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_30
timestamp 1623854003
transform 1 0 3864 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_26
timestamp 1623854003
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1623854003
transform 1 0 4876 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb1
timestamp 1623854003
transform 1 0 4508 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1623854003
transform 1 0 4600 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_44
timestamp 1623854003
transform 1 0 5152 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_44
timestamp 1623854003
transform 1 0 5152 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _342_
timestamp 1623854003
transform -1 0 6624 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1623854003
transform -1 0 5980 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  ringosc.ibufp11
timestamp 1623854003
transform -1 0 6716 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1623854003
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_50
timestamp 1623854003
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_48
timestamp 1623854003
transform 1 0 5520 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_53
timestamp 1623854003
transform 1 0 5980 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1623854003
transform 1 0 7176 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb0
timestamp 1623854003
transform 1 0 7636 0 1 16864
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_1  ringosc.ibufp10
timestamp 1623854003
transform -1 0 7176 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_60
timestamp 1623854003
transform 1 0 6624 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_61
timestamp 1623854003
transform 1 0 6716 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_66
timestamp 1623854003
transform 1 0 7176 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_70
timestamp 1623854003
transform 1 0 7544 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1623854003
transform -1 0 8188 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1623854003
transform 1 0 9568 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1623854003
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_73
timestamp 1623854003
transform 1 0 7820 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_77
timestamp 1623854003
transform 1 0 8188 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1623854003
transform 1 0 8924 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1623854003
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_82
timestamp 1623854003
transform 1 0 8648 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_90
timestamp 1623854003
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen1
timestamp 1623854003
transform 1 0 10580 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb1
timestamp 1623854003
transform -1 0 10580 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1623854003
transform -1 0 10856 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_99
timestamp 1623854003
transform 1 0 10212 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1623854003
transform 1 0 11684 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1623854003
transform 1 0 11040 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1623854003
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_118
timestamp 1623854003
transform 1 0 11960 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_111
timestamp 1623854003
transform 1 0 11316 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_106
timestamp 1623854003
transform 1 0 10856 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _334_
timestamp 1623854003
transform 1 0 12512 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 1623854003
transform 1 0 13432 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[9\].id.delayenb0
timestamp 1623854003
transform 1 0 12420 0 -1 16864
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1623854003
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_122
timestamp 1623854003
transform 1 0 12328 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1623854003
transform 1 0 14076 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_133
timestamp 1623854003
transform 1 0 13340 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1623854003
transform 1 0 14352 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_156
timestamp 1623854003
transform 1 0 15456 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_145
timestamp 1623854003
transform 1 0 14444 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_157
timestamp 1623854003
transform 1 0 15548 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1623854003
transform 1 0 16284 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1623854003
transform -1 0 16836 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1623854003
transform -1 0 16836 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1623854003
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1623854003
transform -1 0 2576 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1623854003
transform -1 0 1656 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_6
timestamp 1623854003
transform 1 0 1656 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_12
timestamp 1623854003
transform 1 0 2208 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_16
timestamp 1623854003
transform 1 0 2576 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen1
timestamp 1623854003
transform 1 0 4140 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1623854003
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1623854003
transform -1 0 4140 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_28
timestamp 1623854003
transform 1 0 3680 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_38
timestamp 1623854003
transform 1 0 4600 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_46
timestamp 1623854003
transform 1 0 5336 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1623854003
transform 1 0 6440 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1623854003
transform -1 0 5796 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output37
timestamp 1623854003
transform -1 0 7268 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_51
timestamp 1623854003
transform 1 0 5796 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_57
timestamp 1623854003
transform 1 0 6348 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_59
timestamp 1623854003
transform 1 0 6532 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_67
timestamp 1623854003
transform 1 0 7268 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1623854003
transform 1 0 9108 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1623854003
transform 1 0 8740 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_79
timestamp 1623854003
transform 1 0 8372 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_86
timestamp 1623854003
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_88
timestamp 1623854003
transform 1 0 9200 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1623854003
transform 1 0 11776 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1623854003
transform 1 0 10120 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1623854003
transform -1 0 12236 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_96
timestamp 1623854003
transform 1 0 9936 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_104
timestamp 1623854003
transform 1 0 10672 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_117
timestamp 1623854003
transform 1 0 11868 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1623854003
transform -1 0 14076 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1623854003
transform 1 0 12236 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_133
timestamp 1623854003
transform 1 0 13340 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_137
timestamp 1623854003
transform 1 0 13708 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1623854003
transform 1 0 14076 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1623854003
transform 1 0 14444 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1623854003
transform -1 0 16560 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1623854003
transform 1 0 15180 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1623854003
transform 1 0 15916 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_146
timestamp 1623854003
transform 1 0 14536 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1623854003
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_156
timestamp 1623854003
transform 1 0 15456 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_160
timestamp 1623854003
transform 1 0 15824 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1623854003
transform -1 0 16836 0 -1 17952
box -38 -48 314 592
<< labels >>
rlabel metal2 s 6918 0 6974 800 4 clockp[0]
port 1 nsew
rlabel metal2 s 6918 19371 6974 20171 4 clockp[1]
port 2 nsew
rlabel metal2 s 10138 19371 10194 20171 4 dco
port 3 nsew
rlabel metal2 s 13818 19371 13874 20171 4 div[0]
port 4 nsew
rlabel metal3 s 17227 3408 18027 3528 4 div[1]
port 5 nsew
rlabel metal3 s 0 2728 800 2848 4 div[2]
port 6 nsew
rlabel metal2 s 1858 0 1914 800 4 div[3]
port 7 nsew
rlabel metal2 s 15198 0 15254 800 4 div[4]
port 8 nsew
rlabel metal2 s 17038 19371 17094 20171 4 enable
port 9 nsew
rlabel metal2 s 8758 19371 8814 20171 4 ext_trim[0]
port 10 nsew
rlabel metal3 s 0 14968 800 15088 4 ext_trim[10]
port 11 nsew
rlabel metal2 s 478 0 534 800 4 ext_trim[11]
port 12 nsew
rlabel metal2 s 3698 19371 3754 20171 4 ext_trim[12]
port 13 nsew
rlabel metal2 s 5538 19371 5594 20171 4 ext_trim[13]
port 14 nsew
rlabel metal2 s 8298 0 8354 800 4 ext_trim[14]
port 15 nsew
rlabel metal3 s 0 7488 800 7608 4 ext_trim[15]
port 16 nsew
rlabel metal3 s 17227 10888 18027 11008 4 ext_trim[16]
port 17 nsew
rlabel metal2 s 3698 0 3754 800 4 ext_trim[17]
port 18 nsew
rlabel metal3 s 17227 1368 18027 1488 4 ext_trim[18]
port 19 nsew
rlabel metal2 s 15198 19371 15254 20171 4 ext_trim[19]
port 20 nsew
rlabel metal3 s 0 10208 800 10328 4 ext_trim[1]
port 21 nsew
rlabel metal2 s 16578 0 16634 800 4 ext_trim[20]
port 22 nsew
rlabel metal3 s 0 12248 800 12368 4 ext_trim[21]
port 23 nsew
rlabel metal3 s 17227 15648 18027 15768 4 ext_trim[22]
port 24 nsew
rlabel metal2 s 2318 19371 2374 20171 4 ext_trim[23]
port 25 nsew
rlabel metal2 s 478 19371 534 20171 4 ext_trim[24]
port 26 nsew
rlabel metal2 s 10138 0 10194 800 4 ext_trim[25]
port 27 nsew
rlabel metal2 s 13358 0 13414 800 4 ext_trim[2]
port 28 nsew
rlabel metal2 s 11978 19371 12034 20171 4 ext_trim[3]
port 29 nsew
rlabel metal2 s 11518 0 11574 800 4 ext_trim[4]
port 30 nsew
rlabel metal3 s 0 17008 800 17128 4 ext_trim[5]
port 31 nsew
rlabel metal2 s 5078 0 5134 800 4 ext_trim[6]
port 32 nsew
rlabel metal3 s 17227 13608 18027 13728 4 ext_trim[7]
port 33 nsew
rlabel metal3 s 17227 6128 18027 6248 4 ext_trim[8]
port 34 nsew
rlabel metal3 s 17227 18368 18027 18488 4 ext_trim[9]
port 35 nsew
rlabel metal3 s 17227 8168 18027 8288 4 osc
port 36 nsew
rlabel metal3 s 0 5448 800 5568 4 resetb
port 37 nsew
rlabel metal4 s 14054 2128 14374 18000 4 VPWR
port 38 nsew
rlabel metal4 s 8810 2128 9130 18000 4 VPWR
port 38 nsew
rlabel metal4 s 3566 2128 3886 18000 4 VPWR
port 38 nsew
rlabel metal5 s 1104 15115 16836 15435 4 VPWR
port 38 nsew
rlabel metal5 s 1104 9856 16836 10176 4 VPWR
port 38 nsew
rlabel metal5 s 1104 4597 16836 4917 4 VPWR
port 38 nsew
rlabel metal4 s 11432 2128 11752 18000 4 VGND
port 39 nsew
rlabel metal4 s 6188 2128 6508 18000 4 VGND
port 39 nsew
rlabel metal5 s 1104 12485 16836 12805 4 VGND
port 39 nsew
rlabel metal5 s 1104 7227 16836 7547 4 VGND
port 39 nsew
<< properties >>
string FIXED_BBOX 0 0 18027 20171
<< end >>
