* NGSPICE file created from digital_pll.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_1 abstract view
.subckt sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_2 abstract view
.subckt sky130_fd_sc_hd__einvn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_4 abstract view
.subckt sky130_fd_sc_hd__einvn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_2 abstract view
.subckt sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_4 abstract view
.subckt sky130_fd_sc_hd__einvp_4 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt digital_pll clockp[0] clockp[1] dco div[0] div[1] div[2] div[3] div[4] enable
+ ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12] ext_trim[13] ext_trim[14] ext_trim[15]
+ ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19] ext_trim[1] ext_trim[20] ext_trim[21]
+ ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25] ext_trim[2] ext_trim[3] ext_trim[4]
+ ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8] ext_trim[9] osc resetb VPWR VGND
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_294_ _297_/C _302_/C _301_/A VGND VGND VPWR VPWR _294_/X sky130_fd_sc_hd__or3_2
X_363_ _328_/A _363_/D _318_/X VGND VGND VPWR VPWR _363_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[1\].id.delayint0 ringosc.dstage\[1\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_346_ _288_/B _346_/A1 _355_/S VGND VGND VPWR VPWR _346_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_277_ _362_/Q _272_/B _363_/Q _267_/B _226_/B VGND VGND VPWR VPWR _359_/D sky130_fd_sc_hd__a311o_1
X_200_ _196_/A _199_/Y _196_/A _199_/Y VGND VGND VPWR VPWR _200_/X sky130_fd_sc_hd__a2bb2o_1
Xringosc.dstage\[11\].id.delayen1 ringosc.dstage\[11\].id.delayen1/A _331_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[11\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
X_329_ _292_/B _232_/B _370_/Q VGND VGND VPWR VPWR _329_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[10\].id.delayenb0 ringosc.dstage\[10\].id.delayenb1/A _332_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[9\].id.delayenb0 ringosc.dstage\[9\].id.delayenb1/A _334_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[9\].id.delayen0/Z sky130_fd_sc_hd__einvn_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_293_ _367_/Q _221_/B _302_/B _370_/Q _232_/B VGND VGND VPWR VPWR _293_/X sky130_fd_sc_hd__o311a_1
X_362_ _328_/A _362_/D _319_/X VGND VGND VPWR VPWR _362_/Q sky130_fd_sc_hd__dfrtp_2
X_345_ _300_/X _345_/A1 _354_/S VGND VGND VPWR VPWR _345_/X sky130_fd_sc_hd__mux2_1
X_276_ _276_/A _276_/B VGND VGND VPWR VPWR _360_/D sky130_fd_sc_hd__or2_1
X_328_ _328_/A VGND VGND VPWR VPWR _328_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_259_ _366_/Q _220_/Y _262_/A VGND VGND VPWR VPWR _259_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[10\].id.delayenb1 ringosc.dstage\[10\].id.delayenb1/A _333_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
Xringosc.dstage\[9\].id.delayenb1 ringosc.dstage\[9\].id.delayenb1/A _335_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[9\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
XFILLER_6_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_292_ _301_/A _292_/B VGND VGND VPWR VPWR _299_/B sky130_fd_sc_hd__nand2_1
X_361_ _328_/A _361_/D _320_/X VGND VGND VPWR VPWR _361_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_344_ _286_/X _344_/A1 _354_/S VGND VGND VPWR VPWR _344_/X sky130_fd_sc_hd__mux2_1
X_275_ _267_/A _267_/B _360_/Q _359_/Q _272_/D VGND VGND VPWR VPWR _276_/B sky130_fd_sc_hd__o221a_1
Xringosc.dstage\[4\].id.delayen0 ringosc.dstage\[4\].id.delayen0/A _344_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_189_ _371_/Q _226_/B VGND VGND VPWR VPWR _371_/D sky130_fd_sc_hd__or2_1
X_327_ _327_/A VGND VGND VPWR VPWR _327_/X sky130_fd_sc_hd__clkbuf_1
X_258_ _262_/A _262_/B VGND VGND VPWR VPWR _258_/X sky130_fd_sc_hd__or2_1
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[5\].id.delayenb0 ringosc.dstage\[5\].id.delayenb1/A _342_/X VGND
+ VGND VPWR VPWR ringosc.ibufp10/A sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[10\].id.delaybuf0 ringosc.dstage\[9\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[9\].id.delaybuf0 ringosc.dstage\[8\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_291_ _369_/Q _368_/Q _367_/Q _370_/Q VGND VGND VPWR VPWR _291_/X sky130_fd_sc_hd__a31o_1
X_360_ _328_/A _360_/D _321_/X VGND VGND VPWR VPWR _360_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_343_ _301_/Y _343_/A1 _355_/S VGND VGND VPWR VPWR _343_/X sky130_fd_sc_hd__mux2_2
X_274_ _272_/D _268_/A _273_/Y _276_/A VGND VGND VPWR VPWR _361_/D sky130_fd_sc_hd__a31o_1
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[4\].id.delayen1 ringosc.dstage\[4\].id.delayen1/A _345_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
X_326_ _370_/Q VGND VGND VPWR VPWR _326_/X sky130_fd_sc_hd__clkbuf_1
X_188_ _372_/Q _272_/D _371_/Q _226_/B VGND VGND VPWR VPWR _372_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_257_ _236_/A _251_/X _256_/Y _368_/Q _236_/Y VGND VGND VPWR VPWR _368_/D sky130_fd_sc_hd__a32o_1
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_309_ _327_/A VGND VGND VPWR VPWR _309_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[10\].id.delaybuf1 ringosc.dstage\[10\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[5\].id.delayenb1 ringosc.dstage\[5\].id.delayenb1/A _343_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[5\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
Xringosc.dstage\[9\].id.delaybuf1 ringosc.dstage\[9\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_290_ _369_/Q _368_/Q _297_/C _370_/Q VGND VGND VPWR VPWR _290_/X sky130_fd_sc_hd__a31o_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_342_ _283_/X _342_/A1 _354_/S VGND VGND VPWR VPWR _342_/X sky130_fd_sc_hd__mux2_2
X_273_ _267_/A _267_/B _267_/C VGND VGND VPWR VPWR _273_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_325_ _327_/A VGND VGND VPWR VPWR _325_/X sky130_fd_sc_hd__clkbuf_1
X_187_ _372_/Q _226_/B _373_/Q _272_/D VGND VGND VPWR VPWR _373_/D sky130_fd_sc_hd__a22o_1
X_256_ _256_/A _256_/B VGND VGND VPWR VPWR _256_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_239_ _288_/A _239_/B VGND VGND VPWR VPWR _239_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_308_ _327_/A VGND VGND VPWR VPWR _308_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[5\].id.delaybuf0 ringosc.dstage\[4\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_341_ _299_/B _341_/A1 _355_/S VGND VGND VPWR VPWR _341_/X sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[1\].id.delayenb0 ringosc.dstage\[1\].id.delayenb1/A _350_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[1\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
X_272_ _362_/Q _272_/B _363_/Q _272_/D VGND VGND VPWR VPWR _276_/A sky130_fd_sc_hd__and4_1
Xringosc.dstage\[8\].id.delayint0 ringosc.dstage\[8\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_5_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_255_ _297_/A _236_/A _254_/X VGND VGND VPWR VPWR _369_/D sky130_fd_sc_hd__o21ai_1
XFILLER_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_186_ _374_/Q _272_/D _359_/Q _226_/B VGND VGND VPWR VPWR _374_/D sky130_fd_sc_hd__a22o_1
X_324_ _327_/A VGND VGND VPWR VPWR _324_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_169_ _374_/Q VGND VGND VPWR VPWR _193_/B sky130_fd_sc_hd__inv_2
X_307_ _327_/A VGND VGND VPWR VPWR _307_/X sky130_fd_sc_hd__clkbuf_1
X_238_ _224_/A _220_/A _224_/B _237_/X VGND VGND VPWR VPWR _262_/A sky130_fd_sc_hd__o22a_1
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput36 _328_/X VGND VGND VPWR VPWR clockp[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[5\].id.delaybuf1 ringosc.dstage\[5\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[1\].id.delayenb1 ringosc.dstage\[1\].id.delayenb1/A _351_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[1\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
XFILLER_12_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_340_ _279_/X _340_/A1 _354_/S VGND VGND VPWR VPWR _340_/X sky130_fd_sc_hd__mux2_1
X_271_ _362_/Q _272_/B _363_/Q _269_/Y _272_/D VGND VGND VPWR VPWR _362_/D sky130_fd_sc_hd__o221a_1
Xringosc.dstage\[1\].id.delayen0 ringosc.dstage\[1\].id.delayen0/A _350_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
X_254_ _244_/Y _253_/A _244_/A _253_/Y _236_/Y VGND VGND VPWR VPWR _254_/X sky130_fd_sc_hd__a221o_1
X_323_ _327_/A VGND VGND VPWR VPWR _323_/X sky130_fd_sc_hd__clkbuf_1
X_185_ _375_/Q _272_/D _360_/Q _226_/B VGND VGND VPWR VPWR _375_/D sky130_fd_sc_hd__a22o_1
X_306_ _327_/A VGND VGND VPWR VPWR _306_/X sky130_fd_sc_hd__clkbuf_1
X_168_ _359_/Q VGND VGND VPWR VPWR _267_/B sky130_fd_sc_hd__inv_2
X_237_ _365_/Q _220_/Y _224_/A _220_/A VGND VGND VPWR VPWR _237_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput37 output37/A VGND VGND VPWR VPWR clockp[1] sky130_fd_sc_hd__clkbuf_2
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_270_ _164_/Y _269_/Y _226_/B VGND VGND VPWR VPWR _363_/D sky130_fd_sc_hd__a21oi_1
Xringosc.dstage\[1\].id.delayen1 ringosc.dstage\[1\].id.delayen1/A _351_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_4_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[1\].id.delaybuf0 ringosc.dstage\[0\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_322_ _327_/A VGND VGND VPWR VPWR _322_/X sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[4\].id.delayint0 ringosc.dstage\[4\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_253_ _253_/A VGND VGND VPWR VPWR _253_/Y sky130_fd_sc_hd__inv_2
X_184_ _376_/Q _272_/D _361_/Q _226_/B VGND VGND VPWR VPWR _376_/D sky130_fd_sc_hd__a22o_1
X_305_ _327_/A VGND VGND VPWR VPWR _305_/X sky130_fd_sc_hd__clkbuf_1
X_167_ _360_/Q VGND VGND VPWR VPWR _267_/A sky130_fd_sc_hd__inv_2
X_236_ _236_/A VGND VGND VPWR VPWR _236_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_219_ _219_/A _219_/B VGND VGND VPWR VPWR _220_/A sky130_fd_sc_hd__or2_4
Xringosc.dstage\[9\].id.delayen0 ringosc.dstage\[9\].id.delayen0/A _334_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[1\].id.delaybuf1 ringosc.dstage\[1\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_252_ _280_/B _220_/A _251_/X VGND VGND VPWR VPWR _253_/A sky130_fd_sc_hd__o21ai_1
X_321_ _327_/A VGND VGND VPWR VPWR _321_/X sky130_fd_sc_hd__clkbuf_1
X_183_ _377_/Q _272_/D _362_/Q _226_/B VGND VGND VPWR VPWR _377_/D sky130_fd_sc_hd__a22o_1
X_304_ _288_/A _239_/B _302_/B _370_/Q _232_/B VGND VGND VPWR VPWR _304_/X sky130_fd_sc_hd__o311a_1
X_235_ _301_/A _220_/Y _224_/X _234_/X VGND VGND VPWR VPWR _236_/A sky130_fd_sc_hd__o31a_4
X_166_ _361_/Q VGND VGND VPWR VPWR _267_/C sky130_fd_sc_hd__inv_2
X_218_ _164_/Y _165_/Y _216_/A _216_/B _214_/X VGND VGND VPWR VPWR _219_/B sky130_fd_sc_hd__o221ai_2
Xringosc.dstage\[9\].id.delayen1 ringosc.dstage\[9\].id.delayen1/A _335_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_251_ _256_/A _256_/B VGND VGND VPWR VPWR _251_/X sky130_fd_sc_hd__or2_1
X_182_ _354_/S _182_/B VGND VGND VPWR VPWR _327_/A sky130_fd_sc_hd__nor2_8
X_320_ _327_/A VGND VGND VPWR VPWR _320_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_303_ _297_/A _368_/Q _367_/Q _302_/X VGND VGND VPWR VPWR _303_/X sky130_fd_sc_hd__o31a_1
X_165_ _378_/Q VGND VGND VPWR VPWR _165_/Y sky130_fd_sc_hd__inv_2
X_234_ _219_/B _225_/Y _220_/A _233_/X _226_/X VGND VGND VPWR VPWR _234_/X sky130_fd_sc_hd__o221a_1
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[0\].id.delayint0 ringosc.dstage\[0\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.iss.reseten0 ringosc.iss.const1/HI _182_/B VGND VGND VPWR VPWR ringosc.ibufp00/A
+ sky130_fd_sc_hd__einvp_4
X_217_ _201_/Y _203_/Y _205_/Y _211_/Y _216_/Y VGND VGND VPWR VPWR _219_/A sky130_fd_sc_hd__o221a_1
XFILLER_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[8\].id.delayenb0 ringosc.dstage\[8\].id.delayenb1/A _336_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[8\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
X_181_ _181_/A _181_/B VGND VGND VPWR VPWR _182_/B sky130_fd_sc_hd__nand2_4
X_250_ _301_/A _236_/A _249_/X VGND VGND VPWR VPWR _370_/D sky130_fd_sc_hd__o21ai_1
XFILLER_24_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_302_ _370_/Q _302_/B _302_/C VGND VGND VPWR VPWR _302_/X sky130_fd_sc_hd__and3_1
X_164_ _363_/Q VGND VGND VPWR VPWR _164_/Y sky130_fd_sc_hd__inv_2
X_233_ _365_/Q _364_/Q _233_/C VGND VGND VPWR VPWR _233_/X sky130_fd_sc_hd__or3_1
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_216_ _216_/A _216_/B VGND VGND VPWR VPWR _216_/Y sky130_fd_sc_hd__nand2_2
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.iss.delayint0 ringosc.iss.delayen1/Z VGND VGND VPWR VPWR ringosc.iss.delayen0/A
+ sky130_fd_sc_hd__clkinv_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater38 _355_/S VGND VGND VPWR VPWR _354_/S sky130_fd_sc_hd__buf_8
XFILLER_16_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[8\].id.delayenb1 ringosc.dstage\[8\].id.delayenb1/A _337_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[8\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
XFILLER_13_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_180_ _378_/Q _272_/D _363_/Q _226_/B VGND VGND VPWR VPWR _378_/D sky130_fd_sc_hd__a22o_1
X_378_ _328_/A _378_/D _327_/X VGND VGND VPWR VPWR _378_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_232_ _370_/Q _232_/B VGND VGND VPWR VPWR _233_/C sky130_fd_sc_hd__or2_1
X_301_ _301_/A _301_/B VGND VGND VPWR VPWR _301_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[6\].id.delayen0 ringosc.dstage\[6\].id.delayen0/A _340_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
X_215_ _214_/A _214_/B _214_/X VGND VGND VPWR VPWR _216_/B sky130_fd_sc_hd__a21bo_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_377_ _328_/A _377_/D _327_/A VGND VGND VPWR VPWR _377_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[4\].id.delayenb0 ringosc.dstage\[4\].id.delayenb1/A _344_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[4\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
Xringosc.dstage\[8\].id.delaybuf0 ringosc.dstage\[7\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_231_ _297_/C _302_/B VGND VGND VPWR VPWR _232_/B sky130_fd_sc_hd__or2_1
X_300_ _221_/A _366_/Q _301_/A _302_/C _296_/X VGND VGND VPWR VPWR _300_/X sky130_fd_sc_hd__o41a_1
Xinput1 dco VGND VGND VPWR VPWR _355_/S sky130_fd_sc_hd__buf_4
Xringosc.dstage\[10\].id.delayen0 ringosc.dstage\[10\].id.delayen0/A _332_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[6\].id.delayen1 ringosc.dstage\[6\].id.delayen1/A _341_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
X_214_ _214_/A _214_/B VGND VGND VPWR VPWR _214_/X sky130_fd_sc_hd__or2_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[4\].id.delayenb1 ringosc.dstage\[4\].id.delayenb1/A _345_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[4\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
Xringosc.dstage\[8\].id.delaybuf1 ringosc.dstage\[8\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_376_ _328_/A _376_/D _305_/X VGND VGND VPWR VPWR _376_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_230_ _302_/B VGND VGND VPWR VPWR _301_/B sky130_fd_sc_hd__inv_2
XFILLER_1_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_359_ _328_/A _359_/D _322_/X VGND VGND VPWR VPWR _359_/Q sky130_fd_sc_hd__dfrtp_1
Xinput2 div[0] VGND VGND VPWR VPWR _177_/A sky130_fd_sc_hd__buf_1
Xringosc.dstage\[10\].id.delayen1 ringosc.dstage\[10\].id.delayen1/A _333_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_10_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_213_ _362_/Q _377_/Q _190_/Y _197_/X VGND VGND VPWR VPWR _214_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_375_ _328_/A _375_/D _306_/X VGND VGND VPWR VPWR _375_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_358_ _328_/A _358_/D _323_/X VGND VGND VPWR VPWR _358_/Q sky130_fd_sc_hd__dfrtp_1
Xringosc.dstage\[4\].id.delaybuf0 ringosc.dstage\[3\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_289_ _297_/A _368_/Q _370_/Q _284_/X VGND VGND VPWR VPWR _289_/X sky130_fd_sc_hd__o31a_1
Xinput3 div[1] VGND VGND VPWR VPWR _207_/A sky130_fd_sc_hd__buf_1
Xringosc.dstage\[7\].id.delayint0 ringosc.dstage\[7\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[0\].id.delayenb0 ringosc.dstage\[0\].id.delayenb1/A _352_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[0\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_212_ _363_/Q _378_/Q _164_/Y _165_/Y VGND VGND VPWR VPWR _214_/A sky130_fd_sc_hd__a22o_1
XFILLER_18_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_374_ _328_/A _374_/D _307_/X VGND VGND VPWR VPWR _374_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_288_ _288_/A _288_/B VGND VGND VPWR VPWR _288_/X sky130_fd_sc_hd__or2_1
Xringosc.dstage\[3\].id.delayen0 ringosc.dstage\[3\].id.delayen0/A _346_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
Xinput4 div[2] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__buf_1
X_357_ _328_/A _357_/D _324_/X VGND VGND VPWR VPWR _358_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[4\].id.delaybuf1 ringosc.dstage\[4\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[0\].id.delayenb1 ringosc.dstage\[0\].id.delayenb1/A _353_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[0\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
X_211_ _207_/A _207_/B _210_/X VGND VGND VPWR VPWR _211_/Y sky130_fd_sc_hd__a21oi_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.iss.delayenb0 ringosc.iss.delayenb1/A ringosc.iss.ctrlen0/X VGND VGND VPWR
+ VPWR ringosc.ibufp00/A sky130_fd_sc_hd__einvn_4
XFILLER_2_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_373_ _328_/A _373_/D _308_/X VGND VGND VPWR VPWR _373_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_287_ _297_/A _368_/Q _370_/Q _288_/A _284_/X VGND VGND VPWR VPWR _287_/X sky130_fd_sc_hd__o41a_1
Xinput5 div[3] VGND VGND VPWR VPWR _202_/A sky130_fd_sc_hd__buf_1
X_356_ _328_/A _356_/D _325_/X VGND VGND VPWR VPWR _357_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_27_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[3\].id.delayen1 ringosc.dstage\[3\].id.delayen1/A _347_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_19_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_210_ _207_/A _207_/B _177_/A _209_/Y _207_/Y VGND VGND VPWR VPWR _210_/X sky130_fd_sc_hd__o221a_1
XFILLER_24_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_339_ _303_/X _339_/A1 _355_/S VGND VGND VPWR VPWR _339_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[0\].id.delaybuf0 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.dstage\[0\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
Xringosc.iss.delayenb1 ringosc.iss.delayenb1/A _355_/X VGND VGND VPWR VPWR ringosc.iss.delayen1/Z
+ sky130_fd_sc_hd__einvn_2
XFILLER_7_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[3\].id.delayint0 ringosc.dstage\[3\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput30 ext_trim[6] VGND VGND VPWR VPWR _340_/A1 sky130_fd_sc_hd__buf_1
XFILLER_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_372_ _328_/A _372_/D _309_/X VGND VGND VPWR VPWR _372_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_355_ _304_/X _355_/A1 _355_/S VGND VGND VPWR VPWR _355_/X sky130_fd_sc_hd__mux2_2
X_286_ _297_/A _368_/Q _370_/Q _367_/Q _284_/X VGND VGND VPWR VPWR _286_/X sky130_fd_sc_hd__o41a_1
Xinput6 div[4] VGND VGND VPWR VPWR _216_/A sky130_fd_sc_hd__buf_1
XFILLER_10_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ _290_/X _338_/A1 _355_/S VGND VGND VPWR VPWR _338_/X sky130_fd_sc_hd__mux2_1
X_269_ _362_/Q _272_/B VGND VGND VPWR VPWR _269_/Y sky130_fd_sc_hd__nand2_1
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[0\].id.delaybuf1 ringosc.dstage\[0\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xinput31 ext_trim[7] VGND VGND VPWR VPWR _338_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput20 ext_trim[20] VGND VGND VPWR VPWR _339_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.iss.delaybuf0 ringosc.iss.delayenb1/A VGND VGND VPWR VPWR ringosc.iss.delayen1/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_371_ _328_/A _371_/D _310_/X VGND VGND VPWR VPWR _371_/Q sky130_fd_sc_hd__dfrtp_1
X_354_ _282_/X _354_/A1 _354_/S VGND VGND VPWR VPWR _354_/X sky130_fd_sc_hd__mux2_1
X_285_ _297_/A _368_/Q _370_/Q _297_/C _284_/X VGND VGND VPWR VPWR _285_/X sky130_fd_sc_hd__o41a_1
XFILLER_6_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput7 enable VGND VGND VPWR VPWR _181_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_337_ _293_/X _337_/A1 _355_/S VGND VGND VPWR VPWR _337_/X sky130_fd_sc_hd__mux2_1
X_268_ _268_/A VGND VGND VPWR VPWR _272_/B sky130_fd_sc_hd__inv_2
X_199_ _361_/Q _376_/Q _192_/Y VGND VGND VPWR VPWR _199_/Y sky130_fd_sc_hd__a21oi_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput21 ext_trim[21] VGND VGND VPWR VPWR _337_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput10 ext_trim[11] VGND VGND VPWR VPWR _330_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput32 ext_trim[8] VGND VGND VPWR VPWR _336_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_370_ _328_/A _370_/D _311_/X VGND VGND VPWR VPWR _370_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_353_ _291_/X _353_/A1 _354_/S VGND VGND VPWR VPWR _353_/X sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[0\].id.delayen0 ringosc.dstage\[0\].id.delayen0/A _352_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
X_284_ _370_/Q _302_/C _288_/B VGND VGND VPWR VPWR _284_/X sky130_fd_sc_hd__o21a_1
Xinput8 ext_trim[0] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[7\].id.delayenb0 ringosc.dstage\[7\].id.delayenb1/A _338_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[7\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
X_336_ _281_/X _336_/A1 _355_/S VGND VGND VPWR VPWR _336_/X sky130_fd_sc_hd__mux2_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_267_ _267_/A _267_/B _267_/C VGND VGND VPWR VPWR _268_/A sky130_fd_sc_hd__or3_1
X_198_ _191_/X _197_/X _191_/X _197_/X VGND VGND VPWR VPWR _202_/B sky130_fd_sc_hd__a2bb2o_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput33 ext_trim[9] VGND VGND VPWR VPWR _334_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput11 ext_trim[12] VGND VGND VPWR VPWR _354_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput22 ext_trim[22] VGND VGND VPWR VPWR _335_/A1 sky130_fd_sc_hd__clkbuf_1
X_319_ _327_/A VGND VGND VPWR VPWR _319_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[0\].id.delayen1 ringosc.dstage\[0\].id.delayen1/A _353_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
Xinput9 ext_trim[10] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
X_283_ _370_/Q _302_/C _288_/A _288_/B VGND VGND VPWR VPWR _283_/X sky130_fd_sc_hd__o31a_1
X_352_ _233_/C input8/X _354_/S VGND VGND VPWR VPWR _352_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_335_ _296_/X _335_/A1 _355_/S VGND VGND VPWR VPWR _335_/X sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[7\].id.delayenb1 ringosc.dstage\[7\].id.delayenb1/A _339_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[7\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_197_ _361_/Q _376_/Q _192_/Y _196_/Y VGND VGND VPWR VPWR _197_/X sky130_fd_sc_hd__o2bb2a_1
XPHY_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_266_ _364_/Q _236_/A _224_/B _236_/Y VGND VGND VPWR VPWR _364_/D sky130_fd_sc_hd__o22a_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 ext_trim[13] VGND VGND VPWR VPWR _353_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput23 ext_trim[23] VGND VGND VPWR VPWR _333_/A1 sky130_fd_sc_hd__clkbuf_1
X_249_ _246_/Y _248_/A _246_/A _248_/Y _236_/Y VGND VGND VPWR VPWR _249_/X sky130_fd_sc_hd__a221o_1
X_318_ _327_/A VGND VGND VPWR VPWR _318_/X sky130_fd_sc_hd__clkbuf_1
Xinput34 osc VGND VGND VPWR VPWR _356_/D sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[8\].id.delayen0 ringosc.dstage\[8\].id.delayen0/A _336_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[8\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_282_ _370_/Q _302_/C _367_/Q _288_/B VGND VGND VPWR VPWR _282_/X sky130_fd_sc_hd__o31a_1
X_351_ _298_/X _351_/A1 _354_/S VGND VGND VPWR VPWR _351_/X sky130_fd_sc_hd__mux2_1
X_334_ _285_/X _334_/A1 _355_/S VGND VGND VPWR VPWR _334_/X sky130_fd_sc_hd__mux2_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_196_ _196_/A VGND VGND VPWR VPWR _196_/Y sky130_fd_sc_hd__inv_2
X_265_ _224_/A _236_/A _236_/Y _264_/X VGND VGND VPWR VPWR _365_/D sky130_fd_sc_hd__o22ai_1
Xinput24 ext_trim[24] VGND VGND VPWR VPWR _331_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput13 ext_trim[14] VGND VGND VPWR VPWR _351_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput35 resetb VGND VGND VPWR VPWR _181_/B sky130_fd_sc_hd__buf_1
X_179_ _272_/D VGND VGND VPWR VPWR _226_/B sky130_fd_sc_hd__clkinv_4
X_317_ _327_/A VGND VGND VPWR VPWR _317_/X sky130_fd_sc_hd__clkbuf_1
X_248_ _248_/A VGND VGND VPWR VPWR _248_/Y sky130_fd_sc_hd__inv_2
Xringosc.dstage\[7\].id.delaybuf0 ringosc.dstage\[6\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[3\].id.delayenb0 ringosc.dstage\[3\].id.delayenb1/A _346_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[3\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[11\].id.delayint0 ringosc.dstage\[11\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_22_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[8\].id.delayen1 ringosc.dstage\[8\].id.delayen1/A _337_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[8\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_281_ _297_/C _302_/C _370_/Q _288_/B VGND VGND VPWR VPWR _281_/X sky130_fd_sc_hd__o31a_1
X_350_ _289_/X _350_/A1 _354_/S VGND VGND VPWR VPWR _350_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_333_ _326_/X _333_/A1 _354_/S VGND VGND VPWR VPWR _333_/X sky130_fd_sc_hd__mux2_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_195_ _360_/Q _375_/Q _193_/Y _194_/X VGND VGND VPWR VPWR _196_/A sky130_fd_sc_hd__a22o_1
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_264_ _224_/B _237_/X _224_/B _237_/X VGND VGND VPWR VPWR _264_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput25 ext_trim[25] VGND VGND VPWR VPWR _355_/A1 sky130_fd_sc_hd__clkbuf_1
X_316_ _327_/A VGND VGND VPWR VPWR _316_/X sky130_fd_sc_hd__clkbuf_1
Xinput14 ext_trim[15] VGND VGND VPWR VPWR _349_/A1 sky130_fd_sc_hd__clkbuf_1
X_247_ _370_/Q _220_/Y _301_/A _220_/A VGND VGND VPWR VPWR _248_/A sky130_fd_sc_hd__o22a_1
Xringosc.dstage\[7\].id.delaybuf1 ringosc.dstage\[7\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[3\].id.delayenb1 ringosc.dstage\[3\].id.delayenb1/A _347_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[3\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
XFILLER_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_178_ _358_/D _358_/Q _358_/D _358_/Q VGND VGND VPWR VPWR _272_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_280_ _369_/Q _280_/B VGND VGND VPWR VPWR _302_/C sky130_fd_sc_hd__or2_4
XFILLER_14_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_332_ _288_/X input9/X _354_/S VGND VGND VPWR VPWR _332_/X sky130_fd_sc_hd__mux2_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_194_ _360_/Q _375_/Q _360_/Q _375_/Q VGND VGND VPWR VPWR _194_/X sky130_fd_sc_hd__o2bb2a_1
XPHY_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_263_ _236_/A _258_/X _262_/Y _366_/Q _236_/Y VGND VGND VPWR VPWR _366_/D sky130_fd_sc_hd__a32o_1
XFILLER_23_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput15 ext_trim[16] VGND VGND VPWR VPWR _347_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput26 ext_trim[2] VGND VGND VPWR VPWR _348_/A1 sky130_fd_sc_hd__buf_1
X_177_ _177_/A VGND VGND VPWR VPWR _177_/Y sky130_fd_sc_hd__inv_2
X_246_ _246_/A VGND VGND VPWR VPWR _246_/Y sky130_fd_sc_hd__inv_2
X_315_ _327_/A VGND VGND VPWR VPWR _315_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_229_ _369_/Q _368_/Q VGND VGND VPWR VPWR _302_/B sky130_fd_sc_hd__or2_4
XFILLER_8_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[3\].id.delaybuf0 ringosc.dstage\[2\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[6\].id.delayint0 ringosc.dstage\[6\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_28_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.ibufp10 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.ibufp11/A sky130_fd_sc_hd__inv_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_331_ _302_/X _331_/A1 _354_/S VGND VGND VPWR VPWR _331_/X sky130_fd_sc_hd__mux2_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_193_ _267_/B _193_/B VGND VGND VPWR VPWR _193_/Y sky130_fd_sc_hd__nor2_4
XPHY_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_262_ _262_/A _262_/B VGND VGND VPWR VPWR _262_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput27 ext_trim[3] VGND VGND VPWR VPWR _346_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_245_ _256_/B _244_/A _256_/A _220_/A _301_/B VGND VGND VPWR VPWR _246_/A sky130_fd_sc_hd__o32a_1
XFILLER_14_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput16 ext_trim[17] VGND VGND VPWR VPWR _345_/A1 sky130_fd_sc_hd__buf_1
X_176_ _364_/Q VGND VGND VPWR VPWR _224_/B sky130_fd_sc_hd__inv_2
X_314_ _327_/A VGND VGND VPWR VPWR _314_/X sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[5\].id.delayen0 ringosc.dstage\[5\].id.delayen0/A _342_/X VGND VGND
+ VPWR VPWR ringosc.ibufp10/A sky130_fd_sc_hd__einvp_2
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[3\].id.delaybuf1 ringosc.dstage\[3\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_228_ _297_/C VGND VGND VPWR VPWR _239_/B sky130_fd_sc_hd__inv_2
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.ibufp11 ringosc.ibufp11/A VGND VGND VPWR VPWR output37/A sky130_fd_sc_hd__inv_2
XFILLER_14_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.ibufp00 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.ibufp01/A sky130_fd_sc_hd__clkinv_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ _287_/X _330_/A1 _354_/S VGND VGND VPWR VPWR _330_/X sky130_fd_sc_hd__mux2_2
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_192_ _361_/Q _376_/Q VGND VGND VPWR VPWR _192_/Y sky130_fd_sc_hd__nor2_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ _367_/Q _260_/X _367_/Q _260_/X VGND VGND VPWR VPWR _367_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_313_ _327_/A VGND VGND VPWR VPWR _313_/X sky130_fd_sc_hd__clkbuf_1
X_244_ _244_/A VGND VGND VPWR VPWR _244_/Y sky130_fd_sc_hd__inv_2
Xinput17 ext_trim[18] VGND VGND VPWR VPWR _343_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput28 ext_trim[4] VGND VGND VPWR VPWR _344_/A1 sky130_fd_sc_hd__buf_1
X_175_ _365_/Q VGND VGND VPWR VPWR _224_/A sky130_fd_sc_hd__inv_2
Xringosc.dstage\[5\].id.delayen1 ringosc.dstage\[5\].id.delayen1/A _343_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[5\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_227_ _367_/Q _366_/Q VGND VGND VPWR VPWR _297_/C sky130_fd_sc_hd__or2_4
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[2\].id.delayint0 ringosc.dstage\[2\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.ibufp01 ringosc.ibufp01/A VGND VGND VPWR VPWR _328_/A sky130_fd_sc_hd__clkinv_8
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_260_ _221_/B _220_/A _236_/A _259_/X VGND VGND VPWR VPWR _260_/X sky130_fd_sc_hd__o211a_1
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_191_ _362_/Q _377_/Q _190_/Y VGND VGND VPWR VPWR _191_/X sky130_fd_sc_hd__a21o_1
XFILLER_23_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput18 ext_trim[19] VGND VGND VPWR VPWR _341_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput29 ext_trim[5] VGND VGND VPWR VPWR _342_/A1 sky130_fd_sc_hd__clkbuf_1
X_312_ _327_/A VGND VGND VPWR VPWR _312_/X sky130_fd_sc_hd__clkbuf_1
X_243_ _297_/A _220_/Y _369_/Q _220_/A VGND VGND VPWR VPWR _244_/A sky130_fd_sc_hd__o22a_1
X_174_ _366_/Q VGND VGND VPWR VPWR _221_/B sky130_fd_sc_hd__inv_2
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[11\].id.delayenb0 ringosc.dstage\[11\].id.delayenb1/A _330_/X VGND
+ VGND VPWR VPWR ringosc.iss.delayenb1/A sky130_fd_sc_hd__einvn_4
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_226_ _372_/Q _226_/B _373_/Q _371_/Q VGND VGND VPWR VPWR _226_/X sky130_fd_sc_hd__and4_1
XFILLER_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_209_ _209_/A VGND VGND VPWR VPWR _209_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_190_ _362_/Q _377_/Q VGND VGND VPWR VPWR _190_/Y sky130_fd_sc_hd__nor2_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_173_ _367_/Q VGND VGND VPWR VPWR _221_/A sky130_fd_sc_hd__inv_2
X_242_ _368_/Q _220_/Y _280_/B _220_/A VGND VGND VPWR VPWR _256_/B sky130_fd_sc_hd__a22o_1
Xinput19 ext_trim[1] VGND VGND VPWR VPWR _350_/A1 sky130_fd_sc_hd__clkbuf_1
X_311_ _327_/A VGND VGND VPWR VPWR _311_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[11\].id.delayenb1 ringosc.dstage\[11\].id.delayenb1/A _331_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[11\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
X_225_ _177_/Y _209_/A _210_/X _205_/A _216_/Y VGND VGND VPWR VPWR _225_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_208_ _267_/B _193_/B _193_/Y VGND VGND VPWR VPWR _209_/A sky130_fd_sc_hd__a21oi_4
XFILLER_28_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_310_ _327_/A VGND VGND VPWR VPWR _310_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_172_ _368_/Q VGND VGND VPWR VPWR _280_/B sky130_fd_sc_hd__inv_2
X_241_ _239_/Y _262_/B _262_/A _220_/A _239_/B VGND VGND VPWR VPWR _256_/A sky130_fd_sc_hd__o32a_1
Xringosc.iss.const1 VGND VGND VPWR VPWR ringosc.iss.const1/HI ringosc.iss.const1/LO
+ sky130_fd_sc_hd__conb_1
Xringosc.dstage\[2\].id.delayen0 ringosc.dstage\[2\].id.delayen0/A _348_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_22_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_224_ _224_/A _224_/B _292_/B VGND VGND VPWR VPWR _224_/X sky130_fd_sc_hd__or3_1
Xringosc.dstage\[6\].id.delayenb0 ringosc.dstage\[6\].id.delayenb1/A _340_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[6\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
Xringosc.dstage\[11\].id.delaybuf0 ringosc.dstage\[10\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_207_ _207_/A _207_/B VGND VGND VPWR VPWR _207_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_171_ _369_/Q VGND VGND VPWR VPWR _297_/A sky130_fd_sc_hd__inv_2
XFILLER_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_240_ _366_/Q _220_/Y _221_/B _220_/A VGND VGND VPWR VPWR _262_/B sky130_fd_sc_hd__a22o_1
Xringosc.dstage\[2\].id.delayen1 ringosc.dstage\[2\].id.delayen1/A _349_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_20_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_369_ _328_/A _369_/D _312_/X VGND VGND VPWR VPWR _369_/Q sky130_fd_sc_hd__dfrtp_2
X_223_ _297_/A _280_/B _223_/C VGND VGND VPWR VPWR _292_/B sky130_fd_sc_hd__or3_1
XFILLER_8_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[6\].id.delayenb1 ringosc.dstage\[6\].id.delayenb1/A _341_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[6\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
Xringosc.dstage\[11\].id.delaybuf1 ringosc.dstage\[11\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_206_ _193_/Y _194_/X _193_/Y _194_/X VGND VGND VPWR VPWR _207_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.iss.delayen0 ringosc.iss.delayen0/A _354_/X VGND VGND VPWR VPWR ringosc.ibufp00/A
+ sky130_fd_sc_hd__einvp_4
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_170_ _370_/Q VGND VGND VPWR VPWR _301_/A sky130_fd_sc_hd__clkinv_4
X_299_ _329_/X _299_/B VGND VGND VPWR VPWR _299_/X sky130_fd_sc_hd__and2_1
X_368_ _328_/A _368_/D _313_/X VGND VGND VPWR VPWR _368_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_222_ _223_/C VGND VGND VPWR VPWR _288_/A sky130_fd_sc_hd__inv_2
XFILLER_10_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_205_ _205_/A VGND VGND VPWR VPWR _205_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[6\].id.delaybuf0 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.dstage\[6\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[2\].id.delayenb0 ringosc.dstage\[2\].id.delayenb1/A _348_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[2\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
Xringosc.dstage\[10\].id.delayint0 ringosc.dstage\[10\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[9\].id.delayint0 ringosc.dstage\[9\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_25_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.iss.delayen1 ringosc.iss.delayen1/A _355_/X VGND VGND VPWR VPWR ringosc.iss.delayen1/Z
+ sky130_fd_sc_hd__einvp_1
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_298_ _301_/A _302_/C _221_/A _297_/X _296_/X VGND VGND VPWR VPWR _298_/X sky130_fd_sc_hd__o311a_1
X_367_ _328_/A _367_/D _314_/X VGND VGND VPWR VPWR _367_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_221_ _221_/A _221_/B VGND VGND VPWR VPWR _223_/C sky130_fd_sc_hd__or2_1
XFILLER_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_204_ input4/X _200_/X _203_/A _201_/Y VGND VGND VPWR VPWR _205_/A sky130_fd_sc_hd__o211a_1
XFILLER_24_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[6\].id.delaybuf1 ringosc.dstage\[6\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[2\].id.delayenb1 ringosc.dstage\[2\].id.delayenb1/A _349_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[2\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_297_ _297_/A _368_/Q _297_/C _301_/A VGND VGND VPWR VPWR _297_/X sky130_fd_sc_hd__or4_4
X_366_ _328_/A _366_/D _315_/X VGND VGND VPWR VPWR _366_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_220_ _220_/A VGND VGND VPWR VPWR _220_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_349_ _295_/X _349_/A1 _354_/S VGND VGND VPWR VPWR _349_/X sky130_fd_sc_hd__mux2_1
X_203_ _203_/A VGND VGND VPWR VPWR _203_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.iss.ctrlen0 _182_/B _354_/X VGND VGND VPWR VPWR ringosc.iss.ctrlen0/X sky130_fd_sc_hd__or2_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[2\].id.delaybuf0 ringosc.dstage\[1\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[5\].id.delayint0 ringosc.dstage\[5\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_26_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_296_ _367_/Q _221_/B _302_/C _301_/A _295_/X VGND VGND VPWR VPWR _296_/X sky130_fd_sc_hd__o41a_2
X_365_ _328_/A _365_/D _316_/X VGND VGND VPWR VPWR _365_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_279_ _367_/Q _288_/B VGND VGND VPWR VPWR _279_/X sky130_fd_sc_hd__or2_1
X_348_ _284_/X _348_/A1 _354_/S VGND VGND VPWR VPWR _348_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_202_ _202_/A _202_/B VGND VGND VPWR VPWR _203_/A sky130_fd_sc_hd__or2_1
XFILLER_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[7\].id.delayen0 ringosc.dstage\[7\].id.delayen0/A _338_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[7\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[2\].id.delaybuf1 ringosc.dstage\[2\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_295_ _301_/A _302_/B _221_/A _294_/X _293_/X VGND VGND VPWR VPWR _295_/X sky130_fd_sc_hd__o311a_1
XFILLER_3_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_364_ _328_/A _364_/D _317_/X VGND VGND VPWR VPWR _364_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_347_ _299_/X _347_/A1 _355_/S VGND VGND VPWR VPWR _347_/X sky130_fd_sc_hd__mux2_1
X_278_ _370_/Q _302_/B VGND VGND VPWR VPWR _288_/B sky130_fd_sc_hd__or2_4
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_201_ _202_/A _202_/B input4/X _200_/X VGND VGND VPWR VPWR _201_/Y sky130_fd_sc_hd__a22oi_2
Xringosc.dstage\[11\].id.delayen0 ringosc.dstage\[11\].id.delayen0/A _330_/X VGND
+ VGND VPWR VPWR ringosc.iss.delayenb1/A sky130_fd_sc_hd__einvp_4
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[7\].id.delayen1 ringosc.dstage\[7\].id.delayen1/A _339_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[7\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
.ends

