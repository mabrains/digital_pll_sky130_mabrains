* NGSPICE file created from digital_pll.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_sc_hd__a22o_1 VGND X B1 VPWR B2 A1 A2 VPB VNB
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_1 abstract view
.subckt sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
.ends

.subckt sky130_fd_sc_hd__einvn_2 TE_B VGND Z VPWR A VPB VNB
X0 a_214_120# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X3 Z A a_214_120# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X5 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_27_47# a_214_120# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR TE_B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VGND TE_B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_214_120# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_sc_hd__inv_2 VGND Y VPWR A VPB VNB
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22a_1 VGND X B1 VPWR B2 A1 A2 VPB VNB
X0 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvn_4 TE_B VGND Z VPWR A VPB VNB
X0 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X4 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X5 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X6 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X7 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND TE_B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR TE_B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

.subckt sky130_fd_sc_hd__o32a_1 VGND X B1 VPWR A1 B2 A2 A3 VPB VNB
X0 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_sc_hd__a41o_4 VGND X B1 VPWR A1 A2 A3 A4 VPB VNB
X0 VPWR A2 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_1079_47# A3 a_889_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_79_21# A1 a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_467_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_467_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_889_47# A3 a_1079_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_79_21# B1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A3 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_467_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A4 a_1079_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_467_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_639_47# A2 a_889_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR A4 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_467_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_889_47# A2 a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_639_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_1079_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 RESET_B Q VGND CLK VPWR VPB VNB D
X0 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_sc_hd__buf_6 VGND X VPWR A VPB VNB
X0 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_1 VGND X B1 VPWR A1 A2 VPB VNB
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_sc_hd__a41o_2 VGND X B1 VPWR A1 A2 A3 A4 VPB VNB
X0 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_381_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A4 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_381_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_549_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_381_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_465_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A2 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_79_21# A1 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvp_4 VGND Z VPWR TE A VPB VNB
X0 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X1 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X4 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X5 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X8 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND TE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR TE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 RESET_B Q VGND CLK VPWR VPB VNB D
X0 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X9 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND X VPWR A VPB VNB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_sc_hd__inv_4 VGND Y VPWR A VPB VNB
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrbp_1 abstract view
.subckt sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_sc_hd__einvp_2 VGND Z VPWR TE A VPB VNB
X0 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X1 VGND TE a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_204_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Z A a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X6 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR TE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VGND TE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_204_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VGND Y B1 VPWR A1 A2 VPB VNB
X0 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND X VPWR A VPB B VNB C
X0 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrbp_2 abstract view
.subckt sky130_fd_sc_hd__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

.subckt sky130_fd_sc_hd__or3_4 VGND X VPWR A VPB B VNB C
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_297# C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_2 VGND Y VPWR A VPB B VNB
X0 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__conb_1 HI VGND VPWR VPB VNB
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_sc_hd__nor2_1 VGND Y VPWR A VPB B VNB
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 RESET_B Q VGND CLK VPWR VPB VNB D
X0 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X25 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X26 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt digital_pll clockc clockd[0] clockd[1] clockd[2] clockd[3] clockp[0] clockp[1]
+ dco div[0] div[1] div[2] div[3] div[4] ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12]
+ ext_trim[13] ext_trim[14] ext_trim[15] ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19]
+ ext_trim[1] ext_trim[20] ext_trim[21] ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25]
+ ext_trim[2] ext_trim[3] ext_trim[4] ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8]
+ ext_trim[9] extclk_sel osc reset sel[0] sel[1] sel[2] VPWR VGND
XFILLER_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_294_ _294_/A _294_/B VGND VGND VPWR VPWR _309_/C sky130_fd_sc_hd__or2_1
X_363_ _320_/X _363_/A1 _379_/S VGND VGND VPWR VPWR _363_/X sky130_fd_sc_hd__mux2_2
XFILLER_36_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[1\].id.delayint0 ringosc.dstage\[1\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_12_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_346_ _348_/A VGND VGND VPWR VPWR _346_/X sky130_fd_sc_hd__clkbuf_1
X_277_ _235_/Y _241_/Y _276_/X _390_/Q _235_/A VGND VGND VPWR VPWR _390_/D sky130_fd_sc_hd__a32o_1
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_200_ VGND _400_/D _385_/Q VPWR _233_/B _400_/Q _284_/D VPWR VGND sky130_fd_sc_hd__a22o_1
XFILLER_2_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[11\].id.delayen1 ringosc.dstage\[11\].id.delayen1/A _355_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[11\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_329_ _348_/A VGND VGND VPWR VPWR _329_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[10\].id.delayenb0 _356_/X VGND ringosc.dstage\[10\].id.delayen0/Z
+ VPWR ringosc.dstage\[10\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
Xringosc.dstage\[9\].id.delayenb0 _358_/X VGND ringosc.dstage\[9\].id.delayen0/Z VPWR
+ ringosc.dstage\[9\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput42 idiv8/D VGND VGND VPWR VPWR clockd[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_362_ _305_/X _362_/A1 _377_/S VGND VGND VPWR VPWR _362_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_293_ _395_/Q _392_/Q _315_/B VGND VGND VPWR VPWR _293_/X sky130_fd_sc_hd__or3_1
XFILLER_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_276_ _389_/Q _276_/B VGND VGND VPWR VPWR _276_/X sky130_fd_sc_hd__or2_1
X_345_ _348_/A VGND VGND VPWR VPWR _345_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_259_ VGND _259_/Y VPWR _259_/A VPWR VGND sky130_fd_sc_hd__inv_2
X_328_ _348_/A VGND VGND VPWR VPWR _328_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[10\].id.delayenb1 _357_/X VGND ringosc.dstage\[10\].id.delayen1/Z
+ VPWR ringosc.dstage\[10\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
Xringosc.dstage\[9\].id.delayenb1 _359_/X VGND ringosc.dstage\[9\].id.delayen1/Z VPWR
+ ringosc.dstage\[9\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_15_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput43 idiv16/D VGND VGND VPWR VPWR clockd[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_361_ _314_/X _361_/A1 _377_/S VGND VGND VPWR VPWR _361_/X sky130_fd_sc_hd__mux2_1
X_292_ _395_/Q _292_/B VGND VGND VPWR VPWR _292_/X sky130_fd_sc_hd__or2_1
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_275_ _235_/Y _269_/X _274_/X _391_/Q _235_/A VGND VGND VPWR VPWR _391_/D sky130_fd_sc_hd__a32o_1
X_344_ _348_/A VGND VGND VPWR VPWR _344_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[4\].id.delayen0 ringosc.dstage\[4\].id.delayen0/A _368_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_189_ VGND _221_/A VPWR _189_/A VPWR VGND sky130_fd_sc_hd__inv_2
X_327_ _348_/A VGND VGND VPWR VPWR _327_/X sky130_fd_sc_hd__clkbuf_1
X_258_ VGND _259_/A _313_/A VPWR _239_/A _395_/Q _239_/Y VPWR VGND sky130_fd_sc_hd__o22a_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput44 _349_/X VGND VGND VPWR VPWR clockp[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[10\].id.delaybuf0 ringosc.dstage\[9\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[9\].id.delaybuf0 ringosc.dstage\[8\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[5\].id.delayenb0 _366_/X VGND ringosc.ibufp10/A VPWR ringosc.dstage\[5\].id.delayenb1/A
+ VPWR VGND sky130_fd_sc_hd__einvn_4
XFILLER_26_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_360_ _303_/X _360_/A1 _377_/S VGND VGND VPWR VPWR _360_/X sky130_fd_sc_hd__mux2_1
X_291_ _395_/Q _315_/B VGND VGND VPWR VPWR _291_/X sky130_fd_sc_hd__or2_1
XFILLER_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_343_ _348_/A VGND VGND VPWR VPWR _343_/X sky130_fd_sc_hd__clkbuf_1
X_274_ _274_/A _274_/B VGND VGND VPWR VPWR _274_/X sky130_fd_sc_hd__or2_1
XFILLER_23_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[4\].id.delayen1 ringosc.dstage\[4\].id.delayen1/A _369_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_9_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_326_ _348_/A VGND VGND VPWR VPWR _326_/X sky130_fd_sc_hd__clkbuf_1
X_257_ VGND _257_/Y VPWR _257_/A VPWR VGND sky130_fd_sc_hd__inv_2
X_188_ VGND _188_/Y VPWR _389_/Q VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_309_ _309_/A _311_/C _309_/C VGND VGND VPWR VPWR _313_/B sky130_fd_sc_hd__or3_1
XFILLER_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput45 idiv2/CLK VGND VGND VPWR VPWR clockp[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[10\].id.delaybuf1 ringosc.dstage\[10\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[9\].id.delaybuf1 ringosc.dstage\[9\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[5\].id.delayenb1 _367_/X VGND ringosc.dstage\[5\].id.delayen1/Z VPWR
+ ringosc.dstage\[5\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_290_ _290_/A _315_/B VGND VGND VPWR VPWR _292_/B sky130_fd_sc_hd__or2_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_342_ _348_/A VGND VGND VPWR VPWR _342_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_273_ _294_/A _235_/Y _272_/X VGND VGND VPWR VPWR _392_/D sky130_fd_sc_hd__o21ai_1
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_325_ _325_/A _325_/B _325_/C VGND VGND VPWR VPWR _350_/S sky130_fd_sc_hd__nor3_2
X_256_ VGND _257_/A _239_/A VPWR _267_/B _310_/B _253_/A _267_/A VPWR VGND sky130_fd_sc_hd__o32a_1
X_187_ VGND _187_/Y VPWR _390_/Q VPWR VGND sky130_fd_sc_hd__inv_2
X_308_ _393_/Q _392_/Q _394_/Q _395_/Q VGND VGND VPWR VPWR _308_/X sky130_fd_sc_hd__a31o_1
X_239_ VGND _239_/Y VPWR _239_/A VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_37_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[5\].id.delaybuf0 ringosc.dstage\[4\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[1\].id.delayenb0 _374_/X VGND ringosc.dstage\[1\].id.delayen0/Z VPWR
+ ringosc.dstage\[1\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
X_341_ _348_/A VGND VGND VPWR VPWR _341_/X sky130_fd_sc_hd__clkbuf_1
X_272_ _247_/Y _271_/A _247_/A _271_/Y _235_/A VGND VGND VPWR VPWR _272_/X sky130_fd_sc_hd__a221o_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[8\].id.delayint0 ringosc.dstage\[8\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_324_ _325_/A _325_/B _324_/C VGND VGND VPWR VPWR _351_/S sky130_fd_sc_hd__nor3_2
X_255_ VGND _310_/B VPWR _315_/B VPWR VGND sky130_fd_sc_hd__inv_2
X_186_ VGND _294_/B VPWR _391_/Q VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_1_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_307_ _392_/Q _391_/Q _297_/A _299_/Y VGND VGND VPWR VPWR _307_/X sky130_fd_sc_hd__a31o_1
X_238_ VGND _239_/A _217_/Y VPWR _218_/Y _221_/X _237_/X _236_/Y VPWR VGND sky130_fd_sc_hd__a41o_4
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[5\].id.delaybuf1 ringosc.dstage\[5\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[1\].id.delayenb1 _375_/X VGND ringosc.dstage\[1\].id.delayen1/Z VPWR
+ ringosc.dstage\[1\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_271_ VGND _271_/Y VPWR _271_/A VPWR VGND sky130_fd_sc_hd__inv_2
X_340_ _348_/A VGND VGND VPWR VPWR _340_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[1\].id.delayen0 ringosc.dstage\[1\].id.delayen0/A _374_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XFILLER_23_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_323_ _325_/A _323_/B _325_/C VGND VGND VPWR VPWR _352_/S sky130_fd_sc_hd__nor3_2
X_254_ _394_/Q _393_/Q VGND VGND VPWR VPWR _315_/B sky130_fd_sc_hd__or2_4
X_185_ VGND _294_/A VPWR _392_/Q VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_306_ _315_/B _306_/B _395_/Q VGND VGND VPWR VPWR _306_/X sky130_fd_sc_hd__or3_1
X_237_ _237_/A _237_/B _237_/C VGND VGND VPWR VPWR _237_/X sky130_fd_sc_hd__or3_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_270_ _294_/B _239_/A _269_/X VGND VGND VPWR VPWR _271_/A sky130_fd_sc_hd__o21ai_1
XFILLER_27_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[1\].id.delayen1 ringosc.dstage\[1\].id.delayen1/A _375_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
X_399_ _328_/X _399_/Q VGND _349_/A VPWR VPWR VGND _399_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_4_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[1\].id.delaybuf0 ringosc.dstage\[0\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_322_ _325_/A _323_/B _324_/C VGND VGND VPWR VPWR _353_/S sky130_fd_sc_hd__nor3_2
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_184_ VGND _311_/C VPWR _393_/Q VPWR VGND sky130_fd_sc_hd__inv_2
X_253_ VGND _253_/Y VPWR _253_/A VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[4\].id.delayint0 ringosc.dstage\[4\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_305_ _394_/Q _393_/Q _290_/A _395_/Q VGND VGND VPWR VPWR _305_/X sky130_fd_sc_hd__a31o_1
X_236_ _230_/Y _231_/X _226_/Y VGND VGND VPWR VPWR _236_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_219_ _387_/Q _402_/Q _206_/Y VGND VGND VPWR VPWR _219_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[9\].id.delayen0 ringosc.dstage\[9\].id.delayen0/A _358_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XFILLER_0_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater46 VGND _377_/S VPWR _379_/S VPWR VGND sky130_fd_sc_hd__buf_6
XFILLER_37_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_398_ _329_/X _398_/Q VGND _349_/A VPWR VPWR VGND _398_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[1\].id.delaybuf1 ringosc.dstage\[1\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_321_ VGND _321_/X _395_/Q VPWR _315_/B _306_/B VPWR VGND sky130_fd_sc_hd__o21a_1
X_252_ VGND _253_/A _394_/Q VPWR _239_/A _309_/A _239_/Y VPWR VGND sky130_fd_sc_hd__o22a_1
X_183_ VGND _309_/A VPWR _394_/Q VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_304_ _392_/Q _391_/Q _393_/Q _297_/A VGND VGND VPWR VPWR _304_/X sky130_fd_sc_hd__a31o_1
XFILLER_24_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_235_ VGND _235_/Y VPWR _235_/A VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_1_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_218_ _218_/A _218_/B VGND VGND VPWR VPWR _218_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput39 _353_/X VGND VGND VPWR VPWR clockc sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[9\].id.delayen1 ringosc.dstage\[9\].id.delayen1/A _359_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_397_ _330_/X _397_/Q VGND _349_/A VPWR VPWR VGND _397_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_23_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_320_ _309_/A _393_/Q _313_/A _392_/Q _315_/X VGND VGND VPWR VPWR _320_/X sky130_fd_sc_hd__o41a_1
X_182_ VGND _313_/A VPWR _395_/Q VPWR VGND sky130_fd_sc_hd__inv_2
X_251_ VGND _267_/B _311_/C VPWR _239_/A _393_/Q _239_/Y VPWR VGND sky130_fd_sc_hd__a22o_1
XFILLER_13_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_303_ _391_/Q _315_/B _300_/Y VGND VGND VPWR VPWR _303_/X sky130_fd_sc_hd__a21o_1
X_234_ VGND _235_/A _233_/Y VPWR _218_/Y _232_/Y _226_/Y _217_/A VPWR VGND sky130_fd_sc_hd__a41o_2
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[0\].id.delayint0 ringosc.dstage\[0\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.iss.reseten0 VGND ringosc.ibufp00/A VPWR _197_/B ringosc.iss.const1/HI VPWR
+ VGND sky130_fd_sc_hd__einvp_4
XFILLER_28_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_217_ VGND _217_/Y VPWR _217_/A VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[8\].id.delayenb0 _360_/X VGND ringosc.dstage\[8\].id.delayen0/Z VPWR
+ ringosc.dstage\[8\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
X_396_ _331_/X _396_/Q VGND _349_/A VPWR VPWR VGND _396_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_250_ VGND _267_/A _239_/A VPWR _269_/B _249_/Y _247_/A _269_/A VPWR VGND sky130_fd_sc_hd__o32a_1
X_181_ VGND _208_/B VPWR _399_/Q VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_379_ _321_/X _379_/A1 _379_/S VGND VGND VPWR VPWR _379_/X sky130_fd_sc_hd__mux2_1
X_302_ _294_/A _297_/Y _299_/A VGND VGND VPWR VPWR _302_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_233_ _397_/Q _233_/B _398_/Q _396_/Q VGND VGND VPWR VPWR _233_/Y sky130_fd_sc_hd__nand4_2
XFILLER_10_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_216_ _176_/Y _177_/Y _218_/A _218_/B _214_/X VGND VGND VPWR VPWR _217_/A sky130_fd_sc_hd__o221a_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.iss.delayint0 ringosc.iss.delayen1/Z VGND VGND VPWR VPWR ringosc.iss.delayen0/A
+ sky130_fd_sc_hd__clkinv_1
XFILLER_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[8\].id.delayenb1 _361_/X VGND ringosc.dstage\[8\].id.delayen1/Z VPWR
+ ringosc.dstage\[8\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
X_395_ _332_/X _395_/Q VGND _349_/A VPWR VPWR VGND _395_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_4_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_180_ VGND _279_/B VPWR _384_/Q VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_378_ _300_/Y _378_/A1 _379_/S VGND VGND VPWR VPWR _378_/X sky130_fd_sc_hd__mux2_1
X_301_ _249_/Y _297_/Y _299_/A VGND VGND VPWR VPWR _301_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_232_ input2/X _227_/X _231_/X VGND VGND VPWR VPWR _232_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[6\].id.delayen0 ringosc.dstage\[6\].id.delayen0/A _364_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
X_215_ _214_/A _214_/B _214_/X VGND VGND VPWR VPWR _218_/B sky130_fd_sc_hd__a21bo_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_394_ _333_/X _394_/Q VGND _349_/A VPWR VPWR VGND _394_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_377_ _308_/X _377_/A1 _377_/S VGND VGND VPWR VPWR _377_/X sky130_fd_sc_hd__mux2_2
Xringosc.dstage\[8\].id.delaybuf0 ringosc.dstage\[7\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[4\].id.delayenb0 _368_/X VGND ringosc.dstage\[4\].id.delayen0/Z VPWR
+ ringosc.dstage\[4\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_300_ _311_/C _294_/A _297_/Y VGND VGND VPWR VPWR _300_/Y sky130_fd_sc_hd__o21ai_1
X_231_ _229_/A _229_/B input2/X _227_/X _230_/A VGND VGND VPWR VPWR _231_/X sky130_fd_sc_hd__o221a_1
Xinput1 dco VGND VGND VPWR VPWR _379_/S sky130_fd_sc_hd__buf_8
Xringosc.dstage\[10\].id.delayen0 ringosc.dstage\[10\].id.delayen0/A _356_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[6\].id.delayen1 ringosc.dstage\[6\].id.delayen1/A _365_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
X_214_ _214_/A _214_/B VGND VGND VPWR VPWR _214_/X sky130_fd_sc_hd__or2_1
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_393_ _334_/X _393_/Q VGND _349_/A VPWR VPWR VGND _393_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_376_ _292_/X input7/X _379_/S VGND VGND VPWR VPWR _376_/X sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[8\].id.delaybuf1 ringosc.dstage\[8\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[4\].id.delayenb1 _369_/X VGND ringosc.dstage\[4\].id.delayen1/Z VPWR
+ ringosc.dstage\[4\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_230_ VGND _230_/Y VPWR _230_/A VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_1_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_359_ _312_/X _359_/A1 _379_/S VGND VGND VPWR VPWR _359_/X sky130_fd_sc_hd__mux2_1
Xinput2 VGND input2/X VPWR div[0] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[10\].id.delayen1 ringosc.dstage\[10\].id.delayen1/A _357_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_213_ _387_/Q _402_/Q _206_/Y _212_/X VGND VGND VPWR VPWR _214_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_392_ _335_/X _392_/Q VGND _349_/A VPWR VPWR VGND _392_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_375_ _316_/X _375_/A1 _379_/S VGND VGND VPWR VPWR _375_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_358_ _301_/Y _358_/A1 _379_/S VGND VGND VPWR VPWR _358_/X sky130_fd_sc_hd__mux2_1
X_289_ _387_/Q _284_/B _388_/Q _279_/B _233_/B VGND VGND VPWR VPWR _384_/D sky130_fd_sc_hd__a311o_1
XFILLER_36_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput3 VGND _229_/A VPWR div[1] VPWR VGND sky130_fd_sc_hd__buf_1
Xringosc.dstage\[4\].id.delaybuf0 ringosc.dstage\[3\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[0\].id.delayenb0 _376_/X VGND ringosc.dstage\[0\].id.delayen0/Z VPWR
+ ringosc.dstage\[0\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_212_ _386_/Q _401_/Q _207_/Y _211_/Y VGND VGND VPWR VPWR _212_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_35_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[7\].id.delayint0 ringosc.dstage\[7\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_18_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xirb VGND irb/Y VPWR irb/A VPWR VGND sky130_fd_sc_hd__inv_4
XFILLER_12_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_391_ _336_/X _391_/Q VGND _349_/A VPWR VPWR VGND _391_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_374_ _299_/Y _374_/A1 _379_/S VGND VGND VPWR VPWR _374_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_357_ _347_/X _357_/A1 _379_/S VGND VGND VPWR VPWR _357_/X sky130_fd_sc_hd__mux2_1
X_288_ _288_/A _288_/B VGND VGND VPWR VPWR _385_/D sky130_fd_sc_hd__or2_1
Xinput4 VGND _190_/A VPWR div[2] VPWR VGND sky130_fd_sc_hd__buf_1
Xringosc.dstage\[3\].id.delayen0 ringosc.dstage\[3\].id.delayen0/A _370_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XFILLER_36_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[4\].id.delaybuf1 ringosc.dstage\[4\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[0\].id.delayenb1 _377_/X VGND ringosc.dstage\[0\].id.delayen1/Z VPWR
+ ringosc.dstage\[0\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_211_ VGND _211_/Y VPWR _211_/A VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.iss.delayenb0 ringosc.iss.ctrlen0/X VGND ringosc.ibufp00/A VPWR ringosc.iss.delayenb1/A
+ VPWR VGND sky130_fd_sc_hd__einvn_4
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_390_ _337_/X _390_/Q VGND _349_/A VPWR VPWR VGND _390_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_373_ _317_/X _373_/A1 _379_/S VGND VGND VPWR VPWR _373_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_356_ _306_/X input8/X _379_/S VGND VGND VPWR VPWR _356_/X sky130_fd_sc_hd__mux2_1
X_287_ _279_/A _279_/B _385_/Q _384_/Q _284_/D VGND VGND VPWR VPWR _288_/B sky130_fd_sc_hd__o221a_1
Xinput5 VGND _189_/A VPWR div[3] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_36_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[3\].id.delayen1 ringosc.dstage\[3\].id.delayen1/A _371_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_210_ VGND _211_/A _208_/Y VPWR _209_/X _385_/Q _400_/Q VPWR VGND sky130_fd_sc_hd__a22o_1
XFILLER_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_339_ _348_/A VGND VGND VPWR VPWR _339_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.iss.delayenb1 _379_/X VGND ringosc.iss.delayen1/Z VPWR ringosc.iss.delayenb1/A
+ VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_21_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[0\].id.delaybuf0 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.dstage\[0\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[3\].id.delayint0 ringosc.dstage\[3\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_14_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput30 ext_trim[7] VGND VGND VPWR VPWR _362_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_372_ _297_/A _372_/A1 _377_/S VGND VGND VPWR VPWR _372_/X sky130_fd_sc_hd__mux2_2
XFILLER_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_355_ _315_/X _355_/A1 _379_/S VGND VGND VPWR VPWR _355_/X sky130_fd_sc_hd__mux2_1
X_286_ _284_/D _280_/A _285_/Y _288_/A VGND VGND VPWR VPWR _386_/D sky130_fd_sc_hd__a31o_1
XFILLER_36_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput6 VGND _218_/A VPWR div[4] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_19_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xidiv16 idiv8/D idiv16/D irb/Y VGND VGND VPWR VPWR idiv16/Q idiv16/D sky130_fd_sc_hd__dfrbp_1
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_338_ _348_/A VGND VGND VPWR VPWR _338_/X sky130_fd_sc_hd__clkbuf_1
X_269_ _269_/A _269_/B VGND VGND VPWR VPWR _269_/X sky130_fd_sc_hd__or2_1
XFILLER_2_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[0\].id.delaybuf1 ringosc.dstage\[0\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput31 ext_trim[8] VGND VGND VPWR VPWR _360_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput20 ext_trim[21] VGND VGND VPWR VPWR _361_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.iss.delaybuf0 ringosc.iss.delayenb1/A VGND VGND VPWR VPWR ringosc.iss.delayen1/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_371_ _318_/X _371_/A1 _379_/S VGND VGND VPWR VPWR _371_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_354_ _307_/X input9/X _377_/S VGND VGND VPWR VPWR _354_/X sky130_fd_sc_hd__mux2_2
X_285_ _279_/A _279_/B _279_/C VGND VGND VPWR VPWR _285_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_36_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput7 VGND input7/X VPWR ext_trim[0] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_337_ _348_/A VGND VGND VPWR VPWR _337_/X sky130_fd_sc_hd__clkbuf_1
X_199_ VGND _401_/D _386_/Q VPWR _233_/B _401_/Q _284_/D VPWR VGND sky130_fd_sc_hd__a22o_1
X_268_ _235_/Y _262_/X _267_/Y _393_/Q _235_/A VGND VGND VPWR VPWR _393_/D sky130_fd_sc_hd__a32o_1
XFILLER_24_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput10 VGND _378_/A1 VPWR ext_trim[12] VPWR VGND sky130_fd_sc_hd__buf_1
Xinput32 ext_trim[9] VGND VGND VPWR VPWR _358_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput21 ext_trim[22] VGND VGND VPWR VPWR _359_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_370_ _291_/X _370_/A1 _379_/S VGND VGND VPWR VPWR _370_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[0\].id.delayen0 ringosc.dstage\[0\].id.delayen0/A _376_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
X_353_ _352_/X _349_/A _353_/S VGND VGND VPWR VPWR _353_/X sky130_fd_sc_hd__mux2_1
X_284_ _387_/Q _284_/B _388_/Q _284_/D VGND VGND VPWR VPWR _288_/A sky130_fd_sc_hd__and4_1
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 ext_trim[10] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_336_ _348_/A VGND VGND VPWR VPWR _336_/X sky130_fd_sc_hd__clkbuf_1
X_267_ _267_/A _267_/B VGND VGND VPWR VPWR _267_/Y sky130_fd_sc_hd__nand2_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[7\].id.delayenb0 _362_/X VGND ringosc.dstage\[7\].id.delayen0/Z VPWR
+ ringosc.dstage\[7\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
X_198_ VGND _402_/D _387_/Q VPWR _233_/B _402_/Q _284_/D VPWR VGND sky130_fd_sc_hd__a22o_1
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput11 ext_trim[13] VGND VGND VPWR VPWR _377_/A1 sky130_fd_sc_hd__clkbuf_1
X_319_ VGND _319_/X _310_/Y VPWR _306_/B _315_/C VPWR VGND sky130_fd_sc_hd__o21a_1
Xinput33 VGND _196_/A VPWR extclk_sel VPWR VGND sky130_fd_sc_hd__buf_1
Xinput22 VGND _357_/A1 VPWR ext_trim[23] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[0\].id.delayen1 ringosc.dstage\[0\].id.delayen1/A _377_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
X_352_ _351_/X idiv2/D _352_/S VGND VGND VPWR VPWR _352_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_283_ _387_/Q _284_/B _388_/Q _281_/Y _284_/D VGND VGND VPWR VPWR _387_/D sky130_fd_sc_hd__o221a_1
Xinput9 VGND input9/X VPWR ext_trim[11] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_197_ _377_/S _197_/B VGND VGND VPWR VPWR _348_/A sky130_fd_sc_hd__nor2_8
Xringosc.dstage\[7\].id.delayenb1 _363_/X VGND ringosc.dstage\[7\].id.delayen1/Z VPWR
+ ringosc.dstage\[7\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
X_335_ _348_/A VGND VGND VPWR VPWR _335_/X sky130_fd_sc_hd__clkbuf_1
X_266_ _309_/A _235_/Y _265_/X VGND VGND VPWR VPWR _394_/D sky130_fd_sc_hd__o21ai_1
XFILLER_32_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput23 ext_trim[24] VGND VGND VPWR VPWR _355_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput12 ext_trim[14] VGND VGND VPWR VPWR _375_/A1 sky130_fd_sc_hd__clkbuf_1
X_249_ VGND _249_/Y VPWR _290_/A VPWR VGND sky130_fd_sc_hd__inv_2
X_318_ _380_/X _318_/B VGND VGND VPWR VPWR _318_/X sky130_fd_sc_hd__and2_1
Xinput34 osc VGND VGND VPWR VPWR _381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[8\].id.delayen0 VGND ringosc.dstage\[8\].id.delayen0/Z VPWR _360_/X
+ ringosc.dstage\[8\].id.delayen0/A VPWR VGND sky130_fd_sc_hd__einvp_2
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_351_ _350_/X idiv4/D _351_/S VGND VGND VPWR VPWR _351_/X sky130_fd_sc_hd__mux2_1
X_282_ VGND _388_/D _233_/B VPWR _176_/Y _281_/Y VPWR VGND sky130_fd_sc_hd__a21oi_1
XFILLER_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_403_ _348_/X _403_/Q VGND _349_/A VPWR VPWR VGND _403_/D sky130_fd_sc_hd__dfrtp_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ _348_/A VGND VGND VPWR VPWR _334_/X sky130_fd_sc_hd__clkbuf_1
X_196_ _196_/A irb/A VGND VGND VPWR VPWR _197_/B sky130_fd_sc_hd__or2_4
X_265_ _253_/Y _264_/A _253_/A _264_/Y _235_/A VGND VGND VPWR VPWR _265_/X sky130_fd_sc_hd__a221o_1
XFILLER_2_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_317_ VGND _317_/X _310_/Y VPWR _290_/A _315_/C VPWR VGND sky130_fd_sc_hd__o21a_1
Xinput13 ext_trim[15] VGND VGND VPWR VPWR _373_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput35 reset VGND VGND VPWR VPWR irb/A sky130_fd_sc_hd__clkbuf_2
X_248_ _392_/Q _391_/Q VGND VGND VPWR VPWR _290_/A sky130_fd_sc_hd__or2_2
X_179_ VGND _279_/A VPWR _385_/Q VPWR VGND sky130_fd_sc_hd__inv_2
Xinput24 VGND _379_/A1 VPWR ext_trim[25] VPWR VGND sky130_fd_sc_hd__buf_1
Xringosc.dstage\[7\].id.delaybuf0 ringosc.dstage\[6\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[3\].id.delayenb0 _370_/X VGND ringosc.dstage\[3\].id.delayen0/Z VPWR
+ ringosc.dstage\[3\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[11\].id.delayint0 ringosc.dstage\[11\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_7_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[8\].id.delayen1 ringosc.dstage\[8\].id.delayen1/A _361_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[8\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_350_ idiv16/D idiv8/D _350_/S VGND VGND VPWR VPWR _350_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_281_ _387_/Q _284_/B VGND VGND VPWR VPWR _281_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_402_ _348_/A _402_/Q VGND _349_/A VPWR VPWR VGND _402_/D sky130_fd_sc_hd__dfrtp_1
X_333_ _348_/A VGND VGND VPWR VPWR _333_/X sky130_fd_sc_hd__clkbuf_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_264_ VGND _264_/Y VPWR _264_/A VPWR VGND sky130_fd_sc_hd__inv_2
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_195_ VGND _403_/D _388_/Q VPWR _233_/B _403_/Q _284_/D VPWR VGND sky130_fd_sc_hd__a22o_1
XFILLER_37_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput25 ext_trim[2] VGND VGND VPWR VPWR _372_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput36 sel[0] VGND VGND VPWR VPWR _324_/C sky130_fd_sc_hd__clkbuf_2
X_316_ _309_/A _393_/Q _313_/A _290_/A _315_/X VGND VGND VPWR VPWR _316_/X sky130_fd_sc_hd__o41a_1
X_247_ VGND _247_/Y VPWR _247_/A VPWR VGND sky130_fd_sc_hd__inv_2
Xinput14 VGND _371_/A1 VPWR ext_trim[16] VPWR VGND sky130_fd_sc_hd__buf_1
X_178_ VGND _279_/C VPWR _386_/Q VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_37_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[7\].id.delaybuf1 ringosc.dstage\[7\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[3\].id.delayenb1 _371_/X VGND ringosc.dstage\[3\].id.delayen1/Z VPWR
+ ringosc.dstage\[3\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_280_ VGND _284_/B VPWR _280_/A VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_401_ _326_/X _401_/Q VGND _349_/A VPWR VPWR VGND _401_/D sky130_fd_sc_hd__dfrtp_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_332_ _348_/A VGND VGND VPWR VPWR _332_/X sky130_fd_sc_hd__clkbuf_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_263_ _311_/C _239_/A _262_/X VGND VGND VPWR VPWR _264_/A sky130_fd_sc_hd__o21ai_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_194_ _284_/D VGND VGND VPWR VPWR _233_/B sky130_fd_sc_hd__clkinv_4
XFILLER_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput37 sel[1] VGND VGND VPWR VPWR _323_/B sky130_fd_sc_hd__buf_2
Xinput15 ext_trim[17] VGND VGND VPWR VPWR _369_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput26 ext_trim[3] VGND VGND VPWR VPWR _370_/A1 sky130_fd_sc_hd__clkbuf_1
X_315_ VGND _315_/X VPWR _395_/Q VPWR _315_/B VGND _315_/C sky130_fd_sc_hd__and3_1
X_246_ VGND _247_/A _392_/Q VPWR _239_/A _294_/A _239_/Y VPWR VGND sky130_fd_sc_hd__o22a_1
X_177_ VGND _177_/Y VPWR _403_/Q VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_229_ _229_/A _229_/B VGND VGND VPWR VPWR _230_/A sky130_fd_sc_hd__nand2_1
Xringosc.dstage\[3\].id.delaybuf0 ringosc.dstage\[2\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[6\].id.delayint0 ringosc.dstage\[6\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.ibufp10 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.ibufp11/A sky130_fd_sc_hd__inv_1
XFILLER_5_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_400_ _327_/X _400_/Q VGND _349_/A VPWR VPWR VGND _400_/D sky130_fd_sc_hd__dfrtp_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ _348_/A VGND VGND VPWR VPWR _331_/X sky130_fd_sc_hd__clkbuf_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_262_ _267_/A _267_/B VGND VGND VPWR VPWR _262_/X sky130_fd_sc_hd__or2_1
X_193_ _383_/D _383_/Q _383_/D _383_/Q VGND VGND VPWR VPWR _284_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_314_ VGND _314_/X _395_/Q VPWR _392_/Q _315_/B VPWR VGND sky130_fd_sc_hd__o21a_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput38 sel[2] VGND VGND VPWR VPWR _325_/A sky130_fd_sc_hd__clkbuf_2
Xinput27 VGND _368_/A1 VPWR ext_trim[4] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_14_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_245_ VGND _269_/B VPWR _274_/B VPWR VGND sky130_fd_sc_hd__inv_2
X_176_ VGND _176_/Y VPWR _388_/Q VPWR VGND sky130_fd_sc_hd__inv_2
Xinput16 VGND _367_/A1 VPWR ext_trim[18] VPWR VGND sky130_fd_sc_hd__buf_1
Xringosc.dstage\[5\].id.delayen0 VGND ringosc.ibufp10/A VPWR _366_/X ringosc.dstage\[5\].id.delayen0/A
+ VPWR VGND sky130_fd_sc_hd__einvp_2
XFILLER_11_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_228_ _208_/Y _209_/X _208_/Y _209_/X VGND VGND VPWR VPWR _229_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[3\].id.delaybuf1 ringosc.dstage\[3\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.ibufp11 VGND idiv2/CLK VPWR ringosc.ibufp11/A VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.ibufp00 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.ibufp01/A sky130_fd_sc_hd__clkinv_2
XFILLER_30_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xidiv2 idiv2/CLK idiv2/D irb/Y VGND VGND VPWR VPWR idiv2/Q idiv2/D sky130_fd_sc_hd__dfrbp_2
XFILLER_35_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ _348_/A VGND VGND VPWR VPWR _330_/X sky130_fd_sc_hd__clkbuf_1
X_192_ VGND _325_/C VPWR _324_/C VPWR VGND sky130_fd_sc_hd__inv_2
X_261_ _313_/A _235_/Y _260_/X VGND VGND VPWR VPWR _395_/D sky130_fd_sc_hd__o21ai_1
XFILLER_2_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_313_ _313_/A _313_/B VGND VGND VPWR VPWR _318_/B sky130_fd_sc_hd__nand2_1
X_244_ VGND _274_/B _391_/Q VPWR _239_/Y _294_/B _239_/A VPWR VGND sky130_fd_sc_hd__o22a_1
Xinput17 ext_trim[19] VGND VGND VPWR VPWR _365_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput28 VGND _366_/A1 VPWR ext_trim[5] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_37_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[5\].id.delayen1 ringosc.dstage\[5\].id.delayen1/A _367_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[5\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_3_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_227_ _279_/B _208_/B _208_/Y VGND VGND VPWR VPWR _227_/X sky130_fd_sc_hd__a21o_1
XFILLER_6_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[2\].id.delayint0 ringosc.dstage\[2\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.ibufp01 ringosc.ibufp01/A VGND VGND VPWR VPWR _349_/A sky130_fd_sc_hd__clkinv_8
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ _257_/Y _259_/A _257_/A _259_/Y _235_/A VGND VGND VPWR VPWR _260_/X sky130_fd_sc_hd__a221o_1
XFILLER_25_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_191_ VGND _325_/B VPWR _323_/B VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_389_ _338_/X _389_/Q VGND _349_/A VPWR VPWR VGND _389_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_36_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_312_ VGND _312_/X _310_/Y VPWR _392_/Q _315_/C VPWR VGND sky130_fd_sc_hd__o21a_1
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_243_ VGND _269_/A VPWR _274_/A VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_36_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput18 VGND _374_/A1 VPWR ext_trim[1] VPWR VGND sky130_fd_sc_hd__buf_1
Xinput29 ext_trim[6] VGND VGND VPWR VPWR _364_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[11\].id.delayenb0 _354_/X VGND ringosc.iss.delayenb1/A VPWR ringosc.dstage\[11\].id.delayenb1/A
+ VPWR VGND sky130_fd_sc_hd__einvn_4
XFILLER_6_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_226_ _237_/A _237_/B _190_/A _225_/A _237_/C VGND VGND VPWR VPWR _226_/Y sky130_fd_sc_hd__a221oi_2
XFILLER_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_209_ _385_/Q _400_/Q _385_/Q _400_/Q VGND VGND VPWR VPWR _209_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xidiv4 idiv2/D idiv4/D irb/Y VGND VGND VPWR VPWR idiv4/Q idiv4/D sky130_fd_sc_hd__dfrbp_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_190_ VGND _237_/A VPWR _190_/A VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_388_ _339_/X _388_/Q VGND _349_/A VPWR VPWR VGND _388_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_311_ VGND _315_/C VPWR _313_/A VPWR _394_/Q VGND _311_/C sky130_fd_sc_hd__or3_4
X_242_ _187_/Y _239_/A _241_/Y VGND VGND VPWR VPWR _274_/A sky130_fd_sc_hd__o21ai_1
Xinput19 ext_trim[20] VGND VGND VPWR VPWR _363_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[11\].id.delayenb1 _355_/X VGND ringosc.dstage\[11\].id.delayen1/Z
+ VPWR ringosc.dstage\[11\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_6_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_225_ VGND _237_/B VPWR _225_/A VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_33_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_208_ VGND _208_/Y VPWR _279_/B VPWR _208_/B VGND sky130_fd_sc_hd__nor2_2
XFILLER_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_387_ _340_/X _387_/Q VGND _349_/A VPWR VPWR VGND _387_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_310_ VGND _310_/Y VPWR _313_/A VPWR _310_/B VGND sky130_fd_sc_hd__nor2_2
XFILLER_36_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[2\].id.delayen0 ringosc.dstage\[2\].id.delayen0/A _372_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
X_241_ _389_/Q _276_/B VGND VGND VPWR VPWR _241_/Y sky130_fd_sc_hd__nand2_1
Xringosc.iss.const1 ringosc.iss.const1/HI VGND VPWR VPWR VGND sky130_fd_sc_hd__conb_1
XFILLER_37_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_224_ _211_/A _223_/Y _211_/A _223_/Y VGND VGND VPWR VPWR _225_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[11\].id.delaybuf0 ringosc.dstage\[10\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_207_ VGND _207_/Y VPWR _386_/Q VPWR _401_/Q VGND sky130_fd_sc_hd__nor2_1
Xringosc.dstage\[6\].id.delayenb0 _364_/X VGND ringosc.dstage\[6\].id.delayen0/Z VPWR
+ ringosc.dstage\[6\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_9_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_386_ _341_/X _386_/Q VGND _349_/A VPWR VPWR VGND _386_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_32_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[2\].id.delayen1 ringosc.dstage\[2\].id.delayen1/A _373_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
X_240_ VGND _276_/B _390_/Q VPWR _239_/Y _187_/Y _239_/A VPWR VGND sky130_fd_sc_hd__o22a_1
X_369_ _319_/X _369_/A1 _379_/S VGND VGND VPWR VPWR _369_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_223_ VGND _223_/Y _207_/Y VPWR _386_/Q _401_/Q VPWR VGND sky130_fd_sc_hd__a21oi_1
XFILLER_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[11\].id.delaybuf1 ringosc.dstage\[11\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_206_ VGND _206_/Y VPWR _387_/Q VPWR _402_/Q VGND sky130_fd_sc_hd__nor2_1
Xringosc.dstage\[6\].id.delayenb1 _365_/X VGND ringosc.dstage\[6\].id.delayen1/Z VPWR
+ ringosc.dstage\[6\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.iss.delayen0 VGND ringosc.ibufp00/A VPWR _378_/X ringosc.iss.delayen0/A VPWR
+ VGND sky130_fd_sc_hd__einvp_4
X_385_ _342_/X _385_/Q VGND _349_/A VPWR VPWR VGND _385_/D sky130_fd_sc_hd__dfrtp_2
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_368_ _302_/Y _368_/A1 _379_/S VGND VGND VPWR VPWR _368_/X sky130_fd_sc_hd__mux2_1
X_299_ VGND _299_/Y VPWR _299_/A VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_222_ _221_/A _221_/B _221_/X VGND VGND VPWR VPWR _237_/C sky130_fd_sc_hd__a21bo_1
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_205_ VGND _214_/A _176_/Y VPWR _177_/Y _388_/Q _403_/Q VPWR VGND sky130_fd_sc_hd__a22o_1
XFILLER_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[6\].id.delaybuf0 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.dstage\[6\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[2\].id.delayenb0 _372_/X VGND ringosc.dstage\[2\].id.delayen0/Z VPWR
+ ringosc.dstage\[2\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[10\].id.delayint0 ringosc.dstage\[10\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[9\].id.delayint0 ringosc.dstage\[9\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xidiv8 idiv4/D idiv8/D irb/Y VGND VGND VPWR VPWR idiv8/Q idiv8/D sky130_fd_sc_hd__dfrbp_2
XFILLER_35_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.iss.delayen1 ringosc.iss.delayen1/A _379_/X VGND VGND VPWR VPWR ringosc.iss.delayen1/Z
+ sky130_fd_sc_hd__einvp_1
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_384_ _343_/X _384_/Q VGND _349_/A VPWR VPWR VGND _384_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_367_ _310_/Y _367_/A1 _377_/S VGND VGND VPWR VPWR _367_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_298_ _394_/Q _311_/C _313_/A _297_/Y VGND VGND VPWR VPWR _299_/A sky130_fd_sc_hd__a31o_1
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_221_ _221_/A _221_/B VGND VGND VPWR VPWR _221_/X sky130_fd_sc_hd__or2_1
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_204_ _396_/Q _233_/B VGND VGND VPWR VPWR _396_/D sky130_fd_sc_hd__or2_1
XFILLER_24_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[6\].id.delaybuf1 ringosc.dstage\[6\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[2\].id.delayenb1 _373_/X VGND ringosc.dstage\[2\].id.delayen1/Z VPWR
+ ringosc.dstage\[2\].id.delayenb1/A VPWR VGND sky130_fd_sc_hd__einvn_2
XFILLER_29_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_383_ _344_/X _383_/Q VGND _349_/A VPWR VPWR VGND _383_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_15_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_366_ _304_/X _366_/A1 _377_/S VGND VGND VPWR VPWR _366_/X sky130_fd_sc_hd__mux2_2
XFILLER_9_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_297_ VGND _297_/Y VPWR _297_/A VPWR VGND sky130_fd_sc_hd__inv_2
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_220_ _212_/X _219_/X _212_/X _219_/X VGND VGND VPWR VPWR _221_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_349_ _349_/A VGND VGND VPWR VPWR _349_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_203_ VGND _397_/D _396_/Q VPWR _233_/B _397_/Q _284_/D VPWR VGND sky130_fd_sc_hd__a22o_1
Xringosc.iss.ctrlen0 _197_/B _378_/X VGND VGND VPWR VPWR ringosc.iss.ctrlen0/X sky130_fd_sc_hd__or2_2
XFILLER_29_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[2\].id.delaybuf0 ringosc.dstage\[1\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_382_ _345_/X _383_/D VGND _349_/A VPWR VPWR VGND _382_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_15_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[5\].id.delayint0 ringosc.dstage\[5\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_365_ _318_/B _365_/A1 _379_/S VGND VGND VPWR VPWR _365_/X sky130_fd_sc_hd__mux2_2
X_296_ _395_/Q _394_/Q VGND VGND VPWR VPWR _297_/A sky130_fd_sc_hd__or2_2
XFILLER_9_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_279_ _279_/A _279_/B _279_/C VGND VGND VPWR VPWR _280_/A sky130_fd_sc_hd__or3_1
X_348_ _348_/A VGND VGND VPWR VPWR _348_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_202_ VGND _398_/D _398_/Q VPWR _284_/D _397_/Q _233_/B VPWR VGND sky130_fd_sc_hd__a22o_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[7\].id.delayen0 VGND ringosc.dstage\[7\].id.delayen0/Z VPWR _362_/X
+ ringosc.dstage\[7\].id.delayen0/A VPWR VGND sky130_fd_sc_hd__einvp_2
XFILLER_18_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[2\].id.delaybuf1 ringosc.dstage\[2\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_381_ _346_/X _382_/D VGND _349_/A VPWR VPWR VGND _381_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_31_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput40 idiv2/D VGND VGND VPWR VPWR clockd[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_295_ VGND _306_/B VPWR _309_/C VPWR VGND sky130_fd_sc_hd__inv_2
X_364_ _293_/X _364_/A1 _377_/S VGND VGND VPWR VPWR _364_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_347_ _395_/Q VGND VGND VPWR VPWR _347_/X sky130_fd_sc_hd__clkbuf_1
X_278_ VGND _389_/D _188_/Y VPWR _235_/A _389_/Q _235_/Y VPWR VGND sky130_fd_sc_hd__o22a_1
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_201_ VGND _399_/D _384_/Q VPWR _233_/B _399_/Q _284_/D VPWR VGND sky130_fd_sc_hd__a22o_1
Xringosc.dstage\[11\].id.delayen0 VGND ringosc.iss.delayenb1/A VPWR _354_/X ringosc.dstage\[11\].id.delayen0/A
+ VPWR VGND sky130_fd_sc_hd__einvp_4
XFILLER_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[7\].id.delayen1 ringosc.dstage\[7\].id.delayen1/A _363_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[7\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_380_ _313_/B _292_/B _395_/Q VGND VGND VPWR VPWR _380_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput41 idiv4/D VGND VGND VPWR VPWR clockd[1] sky130_fd_sc_hd__clkbuf_2
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

