magic
tech sky130A
magscale 1 2
timestamp 1623891339
<< obsli1 >>
rect 1104 2159 16100 16881
<< obsm1 >>
rect 474 2128 16638 16912
<< metal2 >>
rect 5078 18590 5134 19390
rect 11058 18590 11114 19390
rect 16578 18590 16634 19390
rect 478 0 534 800
rect 5998 0 6054 800
rect 11978 0 12034 800
<< obsm2 >>
rect 480 18534 5022 18590
rect 5190 18534 11002 18590
rect 11170 18534 16522 18590
rect 480 856 16632 18534
rect 590 800 5942 856
rect 6110 800 11922 856
rect 12090 800 16632 856
<< metal3 >>
rect 0 17688 800 17808
rect 16446 10208 17246 10328
rect 0 8848 800 8968
rect 16446 1368 17246 1488
<< obsm3 >>
rect 880 17608 16446 17781
rect 800 10408 16446 17608
rect 800 10128 16366 10408
rect 800 9048 16446 10128
rect 880 8768 16446 9048
rect 800 1568 16446 8768
rect 800 1395 16366 1568
<< metal4 >>
rect 3443 2128 3763 16912
rect 5943 2128 6263 16912
rect 8442 2128 8762 16912
rect 10941 2128 11261 16912
rect 13441 2128 13761 16912
<< obsm4 >>
rect 6343 2128 8362 16912
rect 8842 2128 10861 16912
rect 11341 2128 13361 16912
<< metal5 >>
rect 1104 14208 16100 14528
rect 1104 11760 16100 12080
rect 1104 9312 16100 9632
rect 1104 6864 16100 7184
rect 1104 4416 16100 4736
<< labels >>
rlabel metal2 s 5998 0 6054 800 6 clockp[0]
port 1 nsew signal output
rlabel metal2 s 11058 18590 11114 19390 6 clockp[1]
port 2 nsew signal output
rlabel metal2 s 5078 18590 5134 19390 6 div[0]
port 3 nsew signal input
rlabel metal2 s 478 0 534 800 6 div[1]
port 4 nsew signal input
rlabel metal2 s 16578 18590 16634 19390 6 div[2]
port 5 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 div[3]
port 6 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 div[4]
port 7 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 enable
port 8 nsew signal input
rlabel metal3 s 16446 1368 17246 1488 6 osc
port 9 nsew signal input
rlabel metal3 s 16446 10208 17246 10328 6 resetb
port 10 nsew signal input
rlabel metal4 s 13441 2128 13761 16912 6 VPWR
port 11 nsew power bidirectional
rlabel metal4 s 8442 2128 8762 16912 6 VPWR
port 12 nsew power bidirectional
rlabel metal4 s 3443 2128 3763 16912 6 VPWR
port 13 nsew power bidirectional
rlabel metal5 s 1104 14208 16100 14528 6 VPWR
port 14 nsew power bidirectional
rlabel metal5 s 1104 9312 16100 9632 6 VPWR
port 15 nsew power bidirectional
rlabel metal5 s 1104 4416 16100 4736 6 VPWR
port 16 nsew power bidirectional
rlabel metal4 s 10941 2128 11261 16912 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 5943 2128 6263 16912 6 VGND
port 18 nsew ground bidirectional
rlabel metal5 s 1104 11760 16100 12080 6 VGND
port 19 nsew ground bidirectional
rlabel metal5 s 1104 6864 16100 7184 6 VGND
port 20 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 17246 19390
string LEFview TRUE
string GDS_FILE /openLANE_flow/designs/digital_pll/runs/atork_run_2_pwr_gnd/results/magic/digital_pll.gds
string GDS_END 1159804
string GDS_START 486718
<< end >>

