magic
tech sky130A
magscale 1 2
timestamp 1619506813
<< locali >>
rect 6285 16983 6319 17085
rect 16773 17051 16807 17289
rect 14197 16031 14231 16201
rect 5641 10591 5675 10761
rect 14197 5559 14231 5865
<< viali >>
rect 1501 20009 1535 20043
rect 7757 19941 7791 19975
rect 18245 19941 18279 19975
rect 1593 19873 1627 19907
rect 2329 19873 2363 19907
rect 3157 19873 3191 19907
rect 4261 19873 4295 19907
rect 5549 19873 5583 19907
rect 6929 19873 6963 19907
rect 7573 19873 7607 19907
rect 7849 19873 7883 19907
rect 7987 19873 8021 19907
rect 9873 19873 9907 19907
rect 10517 19873 10551 19907
rect 12449 19873 12483 19907
rect 13093 19873 13127 19907
rect 15117 19873 15151 19907
rect 15853 19873 15887 19907
rect 16681 19873 16715 19907
rect 7113 19737 7147 19771
rect 9689 19737 9723 19771
rect 18061 19737 18095 19771
rect 2513 19669 2547 19703
rect 2973 19669 3007 19703
rect 4445 19669 4479 19703
rect 5733 19669 5767 19703
rect 8125 19669 8159 19703
rect 10333 19669 10367 19703
rect 12265 19669 12299 19703
rect 12909 19669 12943 19703
rect 14933 19669 14967 19703
rect 15669 19669 15703 19703
rect 16497 19669 16531 19703
rect 1685 19465 1719 19499
rect 2697 19329 2731 19363
rect 7764 19329 7798 19363
rect 8033 19329 8067 19363
rect 1869 19261 1903 19295
rect 2421 19261 2455 19295
rect 5733 19261 5767 19295
rect 7113 19261 7147 19295
rect 10425 19261 10459 19295
rect 12817 19261 12851 19295
rect 15301 19261 15335 19295
rect 17509 19261 17543 19295
rect 18153 19261 18187 19295
rect 7297 19193 7331 19227
rect 13093 19193 13127 19227
rect 4169 19125 4203 19159
rect 5917 19125 5951 19159
rect 6929 19125 6963 19159
rect 9505 19125 9539 19159
rect 10609 19125 10643 19159
rect 14565 19125 14599 19159
rect 15485 19125 15519 19159
rect 17325 19125 17359 19159
rect 17969 19125 18003 19159
rect 3341 18921 3375 18955
rect 6745 18921 6779 18955
rect 13829 18921 13863 18955
rect 5273 18853 5307 18887
rect 12265 18853 12299 18887
rect 13001 18853 13035 18887
rect 15025 18853 15059 18887
rect 3157 18785 3191 18819
rect 4445 18785 4479 18819
rect 7849 18785 7883 18819
rect 7941 18785 7975 18819
rect 8033 18785 8067 18819
rect 8217 18785 8251 18819
rect 9689 18785 9723 18819
rect 12081 18785 12115 18819
rect 12173 18785 12207 18819
rect 12449 18785 12483 18819
rect 12909 18785 12943 18819
rect 13185 18785 13219 18819
rect 13645 18785 13679 18819
rect 17141 18785 17175 18819
rect 17693 18785 17727 18819
rect 17877 18785 17911 18819
rect 4997 18717 5031 18751
rect 9965 18717 9999 18751
rect 14749 18717 14783 18751
rect 16957 18717 16991 18751
rect 11897 18649 11931 18683
rect 13185 18649 13219 18683
rect 4353 18581 4387 18615
rect 7665 18581 7699 18615
rect 11437 18581 11471 18615
rect 16497 18581 16531 18615
rect 18153 18581 18187 18615
rect 3709 18377 3743 18411
rect 9045 18377 9079 18411
rect 16405 18377 16439 18411
rect 11069 18309 11103 18343
rect 18337 18309 18371 18343
rect 4169 18241 4203 18275
rect 14933 18241 14967 18275
rect 3893 18173 3927 18207
rect 3985 18173 4019 18207
rect 4261 18173 4295 18207
rect 4905 18173 4939 18207
rect 7021 18173 7055 18207
rect 7757 18173 7791 18207
rect 7941 18173 7975 18207
rect 8309 18173 8343 18207
rect 8493 18173 8527 18207
rect 8585 18173 8619 18207
rect 9229 18173 9263 18207
rect 11161 18173 11195 18207
rect 12265 18173 12299 18207
rect 12357 18173 12391 18207
rect 13369 18173 13403 18207
rect 13737 18173 13771 18207
rect 14657 18173 14691 18207
rect 13461 18105 13495 18139
rect 13553 18105 13587 18139
rect 18153 18105 18187 18139
rect 4813 18037 4847 18071
rect 6837 18037 6871 18071
rect 12081 18037 12115 18071
rect 12725 18037 12759 18071
rect 13185 18037 13219 18071
rect 7389 17833 7423 17867
rect 12909 17833 12943 17867
rect 17509 17833 17543 17867
rect 17969 17833 18003 17867
rect 12725 17765 12759 17799
rect 16037 17765 16071 17799
rect 1409 17697 1443 17731
rect 2789 17697 2823 17731
rect 4445 17697 4479 17731
rect 4629 17697 4663 17731
rect 5641 17697 5675 17731
rect 9781 17697 9815 17731
rect 10701 17697 10735 17731
rect 10885 17697 10919 17731
rect 11529 17697 11563 17731
rect 11805 17697 11839 17731
rect 11897 17697 11931 17731
rect 12081 17697 12115 17731
rect 12541 17697 12575 17731
rect 13553 17697 13587 17731
rect 14933 17697 14967 17731
rect 18153 17697 18187 17731
rect 5917 17629 5951 17663
rect 11345 17629 11379 17663
rect 11713 17629 11747 17663
rect 15761 17629 15795 17663
rect 1593 17561 1627 17595
rect 13461 17561 13495 17595
rect 2605 17493 2639 17527
rect 4261 17493 4295 17527
rect 9873 17493 9907 17527
rect 10793 17493 10827 17527
rect 14749 17493 14783 17527
rect 5457 17289 5491 17323
rect 16037 17289 16071 17323
rect 16773 17289 16807 17323
rect 18061 17289 18095 17323
rect 3341 17221 3375 17255
rect 1869 17153 1903 17187
rect 3801 17153 3835 17187
rect 4997 17153 5031 17187
rect 9689 17153 9723 17187
rect 9873 17153 9907 17187
rect 9965 17153 9999 17187
rect 10057 17153 10091 17187
rect 10517 17153 10551 17187
rect 12642 17153 12676 17187
rect 15301 17153 15335 17187
rect 1593 17085 1627 17119
rect 3985 17085 4019 17119
rect 4445 17085 4479 17119
rect 4905 17085 4939 17119
rect 5181 17085 5215 17119
rect 5273 17085 5307 17119
rect 6285 17085 6319 17119
rect 6837 17085 6871 17119
rect 7021 17085 7055 17119
rect 7481 17085 7515 17119
rect 9597 17085 9631 17119
rect 10701 17085 10735 17119
rect 10793 17085 10827 17119
rect 12357 17085 12391 17119
rect 12541 17085 12575 17119
rect 12725 17085 12759 17119
rect 12909 17085 12943 17119
rect 13553 17085 13587 17119
rect 15853 17085 15887 17119
rect 16313 17085 16347 17119
rect 4077 17017 4111 17051
rect 4169 17017 4203 17051
rect 4307 17017 4341 17051
rect 17601 17153 17635 17187
rect 17693 17153 17727 17187
rect 17325 17085 17359 17119
rect 17509 17085 17543 17119
rect 17831 17085 17865 17119
rect 9413 17017 9447 17051
rect 13093 17017 13127 17051
rect 13829 17017 13863 17051
rect 16773 17017 16807 17051
rect 6285 16949 6319 16983
rect 6837 16949 6871 16983
rect 7665 16949 7699 16983
rect 10517 16949 10551 16983
rect 16221 16949 16255 16983
rect 13369 16745 13403 16779
rect 15393 16745 15427 16779
rect 16037 16745 16071 16779
rect 5549 16677 5583 16711
rect 9505 16677 9539 16711
rect 4997 16609 5031 16643
rect 5457 16609 5491 16643
rect 9965 16609 9999 16643
rect 10241 16609 10275 16643
rect 10333 16609 10367 16643
rect 10517 16609 10551 16643
rect 10793 16609 10827 16643
rect 12081 16609 12115 16643
rect 12265 16609 12299 16643
rect 13369 16609 13403 16643
rect 13553 16609 13587 16643
rect 15485 16609 15519 16643
rect 15945 16609 15979 16643
rect 16129 16609 16163 16643
rect 4721 16541 4755 16575
rect 6561 16541 6595 16575
rect 6837 16541 6871 16575
rect 16589 16541 16623 16575
rect 16865 16541 16899 16575
rect 4813 16473 4847 16507
rect 4905 16405 4939 16439
rect 8309 16405 8343 16439
rect 12265 16405 12299 16439
rect 18337 16405 18371 16439
rect 5825 16201 5859 16235
rect 6929 16201 6963 16235
rect 14197 16201 14231 16235
rect 17325 16201 17359 16235
rect 10793 16133 10827 16167
rect 1869 16065 1903 16099
rect 3617 16065 3651 16099
rect 9505 16065 9539 16099
rect 10149 16065 10183 16099
rect 4813 15997 4847 16031
rect 5733 15997 5767 16031
rect 7113 15997 7147 16031
rect 7297 15997 7331 16031
rect 7573 15997 7607 16031
rect 8585 15997 8619 16031
rect 8677 15997 8711 16031
rect 9413 15997 9447 16031
rect 9781 15997 9815 16031
rect 9965 15997 9999 16031
rect 10241 15997 10275 16031
rect 10885 15997 10919 16031
rect 12081 15997 12115 16031
rect 12265 15997 12299 16031
rect 12449 15997 12483 16031
rect 14197 15997 14231 16031
rect 14289 15997 14323 16031
rect 14381 15997 14415 16031
rect 14565 15997 14599 16031
rect 14781 15997 14815 16031
rect 15393 15997 15427 16031
rect 16221 15997 16255 16031
rect 17509 15997 17543 16031
rect 17785 15997 17819 16031
rect 2145 15929 2179 15963
rect 4997 15929 5031 15963
rect 7205 15929 7239 15963
rect 7435 15929 7469 15963
rect 12357 15929 12391 15963
rect 14657 15929 14691 15963
rect 4629 15861 4663 15895
rect 12633 15861 12667 15895
rect 14933 15861 14967 15895
rect 15577 15861 15611 15895
rect 16405 15861 16439 15895
rect 17693 15861 17727 15895
rect 2973 15657 3007 15691
rect 4261 15657 4295 15691
rect 7573 15657 7607 15691
rect 10057 15657 10091 15691
rect 11345 15657 11379 15691
rect 16957 15657 16991 15691
rect 4537 15589 4571 15623
rect 5365 15589 5399 15623
rect 5549 15589 5583 15623
rect 6285 15589 6319 15623
rect 13461 15589 13495 15623
rect 15025 15589 15059 15623
rect 17233 15589 17267 15623
rect 1409 15521 1443 15555
rect 2789 15521 2823 15555
rect 4445 15521 4479 15555
rect 4629 15521 4663 15555
rect 4747 15521 4781 15555
rect 4905 15521 4939 15555
rect 5733 15521 5767 15555
rect 6193 15521 6227 15555
rect 7481 15521 7515 15555
rect 7665 15521 7699 15555
rect 9689 15521 9723 15555
rect 11404 15521 11438 15555
rect 17141 15521 17175 15555
rect 17325 15521 17359 15555
rect 17509 15521 17543 15555
rect 18153 15521 18187 15555
rect 9781 15453 9815 15487
rect 10885 15453 10919 15487
rect 13737 15453 13771 15487
rect 14749 15453 14783 15487
rect 11529 15385 11563 15419
rect 1593 15317 1627 15351
rect 9689 15317 9723 15351
rect 10977 15317 11011 15351
rect 11989 15317 12023 15351
rect 16497 15317 16531 15351
rect 18061 15317 18095 15351
rect 4721 15113 4755 15147
rect 5181 15113 5215 15147
rect 5825 15113 5859 15147
rect 7849 15113 7883 15147
rect 9689 15113 9723 15147
rect 18153 15113 18187 15147
rect 14473 15045 14507 15079
rect 17601 15045 17635 15079
rect 9873 14977 9907 15011
rect 10333 14977 10367 15011
rect 10793 14977 10827 15011
rect 4905 14909 4939 14943
rect 4997 14909 5031 14943
rect 5273 14909 5307 14943
rect 5733 14909 5767 14943
rect 7297 14909 7331 14943
rect 7665 14909 7699 14943
rect 8309 14909 8343 14943
rect 9965 14909 9999 14943
rect 11161 14909 11195 14943
rect 12265 14909 12299 14943
rect 12541 14909 12575 14943
rect 14657 14909 14691 14943
rect 14749 14909 14783 14943
rect 17417 14909 17451 14943
rect 17601 14909 17635 14943
rect 18337 14909 18371 14943
rect 7481 14841 7515 14875
rect 7573 14841 7607 14875
rect 8493 14841 8527 14875
rect 10977 14841 11011 14875
rect 12449 14841 12483 14875
rect 14841 14841 14875 14875
rect 8677 14773 8711 14807
rect 12081 14773 12115 14807
rect 15025 14773 15059 14807
rect 5825 14569 5859 14603
rect 10977 14569 11011 14603
rect 11161 14569 11195 14603
rect 14933 14569 14967 14603
rect 16221 14569 16255 14603
rect 17049 14569 17083 14603
rect 17233 14569 17267 14603
rect 18153 14569 18187 14603
rect 1501 14433 1535 14467
rect 2053 14433 2087 14467
rect 3065 14433 3099 14467
rect 4721 14433 4755 14467
rect 5181 14433 5215 14467
rect 5457 14433 5491 14467
rect 5641 14433 5675 14467
rect 6929 14433 6963 14467
rect 7665 14433 7699 14467
rect 7941 14433 7975 14467
rect 8125 14433 8159 14467
rect 9505 14433 9539 14467
rect 11158 14433 11192 14467
rect 11529 14433 11563 14467
rect 13369 14433 13403 14467
rect 15025 14433 15059 14467
rect 16129 14433 16163 14467
rect 16773 14433 16807 14467
rect 16957 14433 16991 14467
rect 17325 14433 17359 14467
rect 18337 14433 18371 14467
rect 4445 14365 4479 14399
rect 4629 14365 4663 14399
rect 5365 14365 5399 14399
rect 7021 14365 7055 14399
rect 7205 14365 7239 14399
rect 7849 14365 7883 14399
rect 8309 14365 8343 14399
rect 11621 14365 11655 14399
rect 2053 14297 2087 14331
rect 5549 14297 5583 14331
rect 8033 14297 8067 14331
rect 2973 14229 3007 14263
rect 4537 14229 4571 14263
rect 7113 14229 7147 14263
rect 9597 14229 9631 14263
rect 13277 14229 13311 14263
rect 3065 14025 3099 14059
rect 10241 14025 10275 14059
rect 12633 14025 12667 14059
rect 1593 13957 1627 13991
rect 9597 13957 9631 13991
rect 13737 13957 13771 13991
rect 17877 13957 17911 13991
rect 2605 13889 2639 13923
rect 4169 13889 4203 13923
rect 10057 13889 10091 13923
rect 13185 13889 13219 13923
rect 13277 13889 13311 13923
rect 14749 13889 14783 13923
rect 15117 13889 15151 13923
rect 1409 13821 1443 13855
rect 2053 13821 2087 13855
rect 2513 13821 2547 13855
rect 3065 13821 3099 13855
rect 3433 13821 3467 13855
rect 4261 13821 4295 13855
rect 4859 13821 4893 13855
rect 5217 13821 5251 13855
rect 5365 13821 5399 13855
rect 7159 13821 7193 13855
rect 7572 13821 7606 13855
rect 7665 13821 7699 13855
rect 8125 13821 8159 13855
rect 8953 13821 8987 13855
rect 9101 13821 9135 13855
rect 9321 13821 9355 13855
rect 9459 13821 9493 13855
rect 10333 13821 10367 13855
rect 12817 13821 12851 13855
rect 12909 13821 12943 13855
rect 14013 13821 14047 13855
rect 14933 13821 14967 13855
rect 15025 13821 15059 13855
rect 15209 13821 15243 13855
rect 16129 13821 16163 13855
rect 16313 13821 16347 13855
rect 17325 13821 17359 13855
rect 17509 13821 17543 13855
rect 17693 13821 17727 13855
rect 4997 13753 5031 13787
rect 5089 13753 5123 13787
rect 7297 13753 7331 13787
rect 7389 13753 7423 13787
rect 9229 13753 9263 13787
rect 13737 13753 13771 13787
rect 15945 13753 15979 13787
rect 17601 13753 17635 13787
rect 4721 13685 4755 13719
rect 7021 13685 7055 13719
rect 8217 13685 8251 13719
rect 10057 13685 10091 13719
rect 13921 13685 13955 13719
rect 1501 13481 1535 13515
rect 1961 13481 1995 13515
rect 5641 13481 5675 13515
rect 7849 13481 7883 13515
rect 9597 13481 9631 13515
rect 12541 13481 12575 13515
rect 12725 13481 12759 13515
rect 13737 13481 13771 13515
rect 14749 13481 14783 13515
rect 15577 13481 15611 13515
rect 17509 13481 17543 13515
rect 17693 13481 17727 13515
rect 2789 13413 2823 13447
rect 10425 13413 10459 13447
rect 16865 13413 16899 13447
rect 1869 13345 1903 13379
rect 2697 13345 2731 13379
rect 3249 13345 3283 13379
rect 5089 13345 5123 13379
rect 5549 13345 5583 13379
rect 7297 13345 7331 13379
rect 7757 13345 7791 13379
rect 9505 13345 9539 13379
rect 12722 13345 12756 13379
rect 13093 13345 13127 13379
rect 13645 13345 13679 13379
rect 13829 13345 13863 13379
rect 15117 13345 15151 13379
rect 15761 13345 15795 13379
rect 15945 13345 15979 13379
rect 16129 13345 16163 13379
rect 16313 13345 16347 13379
rect 16957 13345 16991 13379
rect 17690 13345 17724 13379
rect 18153 13345 18187 13379
rect 2053 13277 2087 13311
rect 4813 13277 4847 13311
rect 7021 13277 7055 13311
rect 7205 13277 7239 13311
rect 10149 13277 10183 13311
rect 13185 13277 13219 13311
rect 15025 13277 15059 13311
rect 16037 13277 16071 13311
rect 7113 13209 7147 13243
rect 4905 13141 4939 13175
rect 4997 13141 5031 13175
rect 11897 13141 11931 13175
rect 15117 13141 15151 13175
rect 18061 13141 18095 13175
rect 3157 12937 3191 12971
rect 5181 12937 5215 12971
rect 5641 12937 5675 12971
rect 7573 12937 7607 12971
rect 8033 12937 8067 12971
rect 14933 12937 14967 12971
rect 15025 12937 15059 12971
rect 8953 12869 8987 12903
rect 11069 12869 11103 12903
rect 9413 12801 9447 12835
rect 14841 12801 14875 12835
rect 15669 12801 15703 12835
rect 3341 12733 3375 12767
rect 5365 12733 5399 12767
rect 5457 12733 5491 12767
rect 5733 12733 5767 12767
rect 7481 12733 7515 12767
rect 7757 12733 7791 12767
rect 7849 12733 7883 12767
rect 10977 12733 11011 12767
rect 12725 12733 12759 12767
rect 12817 12733 12851 12767
rect 13093 12733 13127 12767
rect 15117 12733 15151 12767
rect 15761 12733 15795 12767
rect 17509 12733 17543 12767
rect 17877 12733 17911 12767
rect 9505 12665 9539 12699
rect 12909 12665 12943 12699
rect 17601 12665 17635 12699
rect 17693 12665 17727 12699
rect 9413 12597 9447 12631
rect 12541 12597 12575 12631
rect 17325 12597 17359 12631
rect 11345 12393 11379 12427
rect 13829 12393 13863 12427
rect 18337 12393 18371 12427
rect 2237 12325 2271 12359
rect 3157 12325 3191 12359
rect 4537 12325 4571 12359
rect 12357 12325 12391 12359
rect 16865 12325 16899 12359
rect 1777 12257 1811 12291
rect 2329 12257 2363 12291
rect 2973 12257 3007 12291
rect 6561 12257 6595 12291
rect 7481 12257 7515 12291
rect 8493 12257 8527 12291
rect 9689 12257 9723 12291
rect 9781 12257 9815 12291
rect 10057 12257 10091 12291
rect 10517 12257 10551 12291
rect 11161 12257 11195 12291
rect 15117 12257 15151 12291
rect 16589 12257 16623 12291
rect 4261 12189 4295 12223
rect 6653 12189 6687 12223
rect 9965 12189 9999 12223
rect 12081 12189 12115 12223
rect 9505 12121 9539 12155
rect 6009 12053 6043 12087
rect 7665 12053 7699 12087
rect 8401 12053 8435 12087
rect 10609 12053 10643 12087
rect 15301 12053 15335 12087
rect 2237 11849 2271 11883
rect 3065 11849 3099 11883
rect 4537 11849 4571 11883
rect 5549 11849 5583 11883
rect 7100 11849 7134 11883
rect 8585 11849 8619 11883
rect 9873 11849 9907 11883
rect 13369 11849 13403 11883
rect 17969 11849 18003 11883
rect 9505 11781 9539 11815
rect 1593 11713 1627 11747
rect 1777 11713 1811 11747
rect 2697 11713 2731 11747
rect 4813 11713 4847 11747
rect 6837 11713 6871 11747
rect 9413 11713 9447 11747
rect 14473 11713 14507 11747
rect 16221 11713 16255 11747
rect 3065 11645 3099 11679
rect 4721 11645 4755 11679
rect 4905 11645 4939 11679
rect 4997 11645 5031 11679
rect 5733 11645 5767 11679
rect 9137 11645 9171 11679
rect 9321 11645 9355 11679
rect 9597 11645 9631 11679
rect 10609 11645 10643 11679
rect 10793 11645 10827 11679
rect 13553 11645 13587 11679
rect 14197 11645 14231 11679
rect 17509 11645 17543 11679
rect 18153 11645 18187 11679
rect 1869 11577 1903 11611
rect 10793 11509 10827 11543
rect 17325 11509 17359 11543
rect 1501 11305 1535 11339
rect 2881 11305 2915 11339
rect 4261 11305 4295 11339
rect 5181 11305 5215 11339
rect 7665 11305 7699 11339
rect 8585 11305 8619 11339
rect 10241 11305 10275 11339
rect 11345 11305 11379 11339
rect 11805 11305 11839 11339
rect 17877 11305 17911 11339
rect 6101 11237 6135 11271
rect 6285 11237 6319 11271
rect 10149 11237 10183 11271
rect 12449 11237 12483 11271
rect 16405 11237 16439 11271
rect 1593 11169 1627 11203
rect 2789 11169 2823 11203
rect 4629 11169 4663 11203
rect 5273 11169 5307 11203
rect 6929 11169 6963 11203
rect 7573 11169 7607 11203
rect 8217 11169 8251 11203
rect 8309 11169 8343 11203
rect 11437 11169 11471 11203
rect 12633 11169 12667 11203
rect 4537 11101 4571 11135
rect 6469 11101 6503 11135
rect 9965 11101 9999 11135
rect 11253 11101 11287 11135
rect 16129 11101 16163 11135
rect 7021 11033 7055 11067
rect 10609 11033 10643 11067
rect 4629 10965 4663 10999
rect 8309 10965 8343 10999
rect 12817 10965 12851 10999
rect 4905 10761 4939 10795
rect 5641 10761 5675 10795
rect 5825 10761 5859 10795
rect 9689 10761 9723 10795
rect 11069 10761 11103 10795
rect 12081 10761 12115 10795
rect 2789 10693 2823 10727
rect 3249 10693 3283 10727
rect 18153 10693 18187 10727
rect 8401 10625 8435 10659
rect 9781 10625 9815 10659
rect 12449 10625 12483 10659
rect 13553 10625 13587 10659
rect 2421 10557 2455 10591
rect 3433 10557 3467 10591
rect 4629 10557 4663 10591
rect 5641 10557 5675 10591
rect 5733 10557 5767 10591
rect 7021 10557 7055 10591
rect 8309 10557 8343 10591
rect 8585 10557 8619 10591
rect 9505 10557 9539 10591
rect 9873 10557 9907 10591
rect 9965 10557 9999 10591
rect 10241 10557 10275 10591
rect 12265 10557 12299 10591
rect 13369 10557 13403 10591
rect 13461 10557 13495 10591
rect 14841 10557 14875 10591
rect 15393 10557 15427 10591
rect 18337 10557 18371 10591
rect 4813 10489 4847 10523
rect 6837 10489 6871 10523
rect 9045 10489 9079 10523
rect 10701 10489 10735 10523
rect 10885 10489 10919 10523
rect 15301 10489 15335 10523
rect 2789 10421 2823 10455
rect 7113 10421 7147 10455
rect 13001 10421 13035 10455
rect 10867 10217 10901 10251
rect 11345 10217 11379 10251
rect 17049 10217 17083 10251
rect 4813 10149 4847 10183
rect 11161 10149 11195 10183
rect 13461 10149 13495 10183
rect 15485 10149 15519 10183
rect 2237 10081 2271 10115
rect 2789 10081 2823 10115
rect 4905 10081 4939 10115
rect 5917 10081 5951 10115
rect 6745 10081 6779 10115
rect 6837 10081 6871 10115
rect 7297 10081 7331 10115
rect 8309 10081 8343 10115
rect 8401 10081 8435 10115
rect 9597 10081 9631 10115
rect 9781 10081 9815 10115
rect 12265 10081 12299 10115
rect 13277 10081 13311 10115
rect 13553 10081 13587 10115
rect 15577 10081 15611 10115
rect 17141 10081 17175 10115
rect 4813 10013 4847 10047
rect 5641 10013 5675 10047
rect 5733 10013 5767 10047
rect 5825 10013 5859 10047
rect 6561 10013 6595 10047
rect 7389 10013 7423 10047
rect 7573 10013 7607 10047
rect 8125 10013 8159 10047
rect 9505 10013 9539 10047
rect 11437 10013 11471 10047
rect 12983 10013 13017 10047
rect 15669 10013 15703 10047
rect 16865 10013 16899 10047
rect 2789 9945 2823 9979
rect 5457 9945 5491 9979
rect 9965 9945 9999 9979
rect 12449 9945 12483 9979
rect 15117 9945 15151 9979
rect 4353 9877 4387 9911
rect 6653 9877 6687 9911
rect 7481 9877 7515 9911
rect 17509 9877 17543 9911
rect 7665 9673 7699 9707
rect 5457 9605 5491 9639
rect 15393 9605 15427 9639
rect 15853 9605 15887 9639
rect 18153 9605 18187 9639
rect 1685 9537 1719 9571
rect 4629 9537 4663 9571
rect 7389 9537 7423 9571
rect 13277 9537 13311 9571
rect 15025 9537 15059 9571
rect 2881 9469 2915 9503
rect 4721 9469 4755 9503
rect 4813 9469 4847 9503
rect 4905 9469 4939 9503
rect 5641 9469 5675 9503
rect 5825 9469 5859 9503
rect 7205 9469 7239 9503
rect 7297 9469 7331 9503
rect 7481 9469 7515 9503
rect 8677 9469 8711 9503
rect 8861 9469 8895 9503
rect 8953 9469 8987 9503
rect 9413 9469 9447 9503
rect 12909 9469 12943 9503
rect 16037 9469 16071 9503
rect 18337 9469 18371 9503
rect 1777 9401 1811 9435
rect 2697 9401 2731 9435
rect 1869 9333 1903 9367
rect 2237 9333 2271 9367
rect 4445 9333 4479 9367
rect 8493 9333 8527 9367
rect 9505 9333 9539 9367
rect 12909 9333 12943 9367
rect 15393 9333 15427 9367
rect 2881 9129 2915 9163
rect 9710 9129 9744 9163
rect 11253 9129 11287 9163
rect 15577 9129 15611 9163
rect 17601 9129 17635 9163
rect 9505 9061 9539 9095
rect 12633 9061 12667 9095
rect 14841 9061 14875 9095
rect 15025 9061 15059 9095
rect 1593 8993 1627 9027
rect 3065 8993 3099 9027
rect 5170 8993 5204 9027
rect 5917 8993 5951 9027
rect 6561 8993 6595 9027
rect 7297 8993 7331 9027
rect 8309 8993 8343 9027
rect 11345 8993 11379 9027
rect 12541 8993 12575 9027
rect 13093 8993 13127 9027
rect 16497 8993 16531 9027
rect 17233 8993 17267 9027
rect 18245 8993 18279 9027
rect 3341 8925 3375 8959
rect 5089 8925 5123 8959
rect 5273 8925 5307 8959
rect 5365 8925 5399 8959
rect 6009 8925 6043 8959
rect 6653 8925 6687 8959
rect 6837 8925 6871 8959
rect 7389 8925 7423 8959
rect 8585 8925 8619 8959
rect 11161 8925 11195 8959
rect 1409 8857 1443 8891
rect 6745 8857 6779 8891
rect 8493 8857 8527 8891
rect 17601 8857 17635 8891
rect 18061 8857 18095 8891
rect 3249 8789 3283 8823
rect 4905 8789 4939 8823
rect 8125 8789 8159 8823
rect 9689 8789 9723 8823
rect 9873 8789 9907 8823
rect 11713 8789 11747 8823
rect 15669 8789 15703 8823
rect 16589 8789 16623 8823
rect 2237 8585 2271 8619
rect 2697 8585 2731 8619
rect 5181 8585 5215 8619
rect 9413 8585 9447 8619
rect 11161 8585 11195 8619
rect 12081 8585 12115 8619
rect 13001 8585 13035 8619
rect 4445 8517 4479 8551
rect 9781 8517 9815 8551
rect 15853 8517 15887 8551
rect 3065 8449 3099 8483
rect 4077 8449 4111 8483
rect 5641 8449 5675 8483
rect 5825 8449 5859 8483
rect 8769 8449 8803 8483
rect 15485 8449 15519 8483
rect 17693 8449 17727 8483
rect 1685 8381 1719 8415
rect 2237 8381 2271 8415
rect 2697 8381 2731 8415
rect 7113 8381 7147 8415
rect 9321 8381 9355 8415
rect 9597 8381 9631 8415
rect 10609 8381 10643 8415
rect 11161 8381 11195 8415
rect 12081 8381 12115 8415
rect 12449 8381 12483 8415
rect 12909 8381 12943 8415
rect 14473 8381 14507 8415
rect 15025 8381 15059 8415
rect 17325 8381 17359 8415
rect 17877 8381 17911 8415
rect 3893 8313 3927 8347
rect 3985 8313 4019 8347
rect 5549 8313 5583 8347
rect 8585 8313 8619 8347
rect 14933 8313 14967 8347
rect 6929 8245 6963 8279
rect 8125 8245 8159 8279
rect 8493 8245 8527 8279
rect 15853 8245 15887 8279
rect 2697 8041 2731 8075
rect 11989 8041 12023 8075
rect 13277 8041 13311 8075
rect 17601 8041 17635 8075
rect 3157 7973 3191 8007
rect 4445 7973 4479 8007
rect 4629 7973 4663 8007
rect 7481 7973 7515 8007
rect 11161 7973 11195 8007
rect 2513 7905 2547 7939
rect 7297 7905 7331 7939
rect 9505 7905 9539 7939
rect 9689 7905 9723 7939
rect 10977 7905 11011 7939
rect 11805 7905 11839 7939
rect 12909 7905 12943 7939
rect 16773 7905 16807 7939
rect 17417 7905 17451 7939
rect 4353 7837 4387 7871
rect 16405 7837 16439 7871
rect 4905 7769 4939 7803
rect 13277 7769 13311 7803
rect 3249 7701 3283 7735
rect 9505 7701 9539 7735
rect 9873 7701 9907 7735
rect 11345 7701 11379 7735
rect 16773 7701 16807 7735
rect 13369 7497 13403 7531
rect 16313 7497 16347 7531
rect 11069 7429 11103 7463
rect 5457 7361 5491 7395
rect 1777 7293 1811 7327
rect 2329 7293 2363 7327
rect 3985 7293 4019 7327
rect 4261 7293 4295 7327
rect 5733 7293 5767 7327
rect 7021 7293 7055 7327
rect 7573 7293 7607 7327
rect 12817 7293 12851 7327
rect 13369 7293 13403 7327
rect 15761 7293 15795 7327
rect 16313 7293 16347 7327
rect 2237 7225 2271 7259
rect 4169 7225 4203 7259
rect 5917 7225 5951 7259
rect 10885 7225 10919 7259
rect 3801 7157 3835 7191
rect 7941 7157 7975 7191
rect 8677 7157 8711 7191
rect 8769 7157 8803 7191
rect 2145 6953 2179 6987
rect 12081 6953 12115 6987
rect 13185 6953 13219 6987
rect 13645 6953 13679 6987
rect 4721 6885 4755 6919
rect 4813 6885 4847 6919
rect 4997 6885 5031 6919
rect 15117 6885 15151 6919
rect 16497 6885 16531 6919
rect 3341 6817 3375 6851
rect 6193 6817 6227 6851
rect 6653 6817 6687 6851
rect 7573 6817 7607 6851
rect 8033 6817 8067 6851
rect 8585 6817 8619 6851
rect 9965 6817 9999 6851
rect 10609 6817 10643 6851
rect 10885 6817 10919 6851
rect 13829 6817 13863 6851
rect 15209 6817 15243 6851
rect 18337 6817 18371 6851
rect 2237 6749 2271 6783
rect 2421 6749 2455 6783
rect 2973 6749 3007 6783
rect 6929 6749 6963 6783
rect 11805 6749 11839 6783
rect 11989 6749 12023 6783
rect 15301 6749 15335 6783
rect 1777 6681 1811 6715
rect 5273 6681 5307 6715
rect 18153 6681 18187 6715
rect 3341 6613 3375 6647
rect 8585 6613 8619 6647
rect 12449 6613 12483 6647
rect 13093 6613 13127 6647
rect 14749 6613 14783 6647
rect 16405 6613 16439 6647
rect 1593 6409 1627 6443
rect 12725 6341 12759 6375
rect 4077 6273 4111 6307
rect 10885 6273 10919 6307
rect 14657 6273 14691 6307
rect 1409 6205 1443 6239
rect 7021 6205 7055 6239
rect 7941 6205 7975 6239
rect 8401 6205 8435 6239
rect 9137 6205 9171 6239
rect 9321 6205 9355 6239
rect 10241 6205 10275 6239
rect 10977 6205 11011 6239
rect 12357 6205 12391 6239
rect 14841 6205 14875 6239
rect 15025 6205 15059 6239
rect 15301 6205 15335 6239
rect 15853 6205 15887 6239
rect 16037 6205 16071 6239
rect 16221 6205 16255 6239
rect 4537 6137 4571 6171
rect 4629 6137 4663 6171
rect 5089 6137 5123 6171
rect 7665 6137 7699 6171
rect 5273 6069 5307 6103
rect 12725 6069 12759 6103
rect 15853 6069 15887 6103
rect 5641 5865 5675 5899
rect 6653 5865 6687 5899
rect 7021 5865 7055 5899
rect 8585 5865 8619 5899
rect 10793 5865 10827 5899
rect 14197 5865 14231 5899
rect 15025 5865 15059 5899
rect 15485 5865 15519 5899
rect 17141 5865 17175 5899
rect 3065 5797 3099 5831
rect 4905 5797 4939 5831
rect 12541 5797 12575 5831
rect 3249 5729 3283 5763
rect 4261 5729 4295 5763
rect 5181 5729 5215 5763
rect 6009 5729 6043 5763
rect 7113 5729 7147 5763
rect 8217 5729 8251 5763
rect 9689 5729 9723 5763
rect 10701 5729 10735 5763
rect 12081 5729 12115 5763
rect 12633 5729 12667 5763
rect 5641 5661 5675 5695
rect 7297 5661 7331 5695
rect 8585 5593 8619 5627
rect 9505 5593 9539 5627
rect 15117 5729 15151 5763
rect 16129 5729 16163 5763
rect 16313 5729 16347 5763
rect 16497 5729 16531 5763
rect 17049 5729 17083 5763
rect 14933 5661 14967 5695
rect 15945 5661 15979 5695
rect 14197 5525 14231 5559
rect 15025 5321 15059 5355
rect 16313 5321 16347 5355
rect 7205 5253 7239 5287
rect 10517 5253 10551 5287
rect 10977 5253 11011 5287
rect 5273 5185 5307 5219
rect 15669 5185 15703 5219
rect 17785 5185 17819 5219
rect 2754 5117 2788 5151
rect 3341 5117 3375 5151
rect 4905 5117 4939 5151
rect 5457 5117 5491 5151
rect 6837 5117 6871 5151
rect 7021 5117 7055 5151
rect 10149 5117 10183 5151
rect 11161 5117 11195 5151
rect 12633 5117 12667 5151
rect 13369 5117 13403 5151
rect 16405 5117 16439 5151
rect 17325 5117 17359 5151
rect 17601 5117 17635 5151
rect 12449 5049 12483 5083
rect 15393 5049 15427 5083
rect 2651 4981 2685 5015
rect 3433 4981 3467 5015
rect 10517 4981 10551 5015
rect 13185 4981 13219 5015
rect 15485 4981 15519 5015
rect 17417 4981 17451 5015
rect 1501 4777 1535 4811
rect 5641 4777 5675 4811
rect 13277 4777 13311 4811
rect 16037 4777 16071 4811
rect 18153 4777 18187 4811
rect 10517 4709 10551 4743
rect 1593 4641 1627 4675
rect 2421 4641 2455 4675
rect 5825 4641 5859 4675
rect 6285 4641 6319 4675
rect 6469 4641 6503 4675
rect 10057 4641 10091 4675
rect 10609 4641 10643 4675
rect 12449 4641 12483 4675
rect 16405 4641 16439 4675
rect 18337 4641 18371 4675
rect 7297 4573 7331 4607
rect 7665 4573 7699 4607
rect 11621 4573 11655 4607
rect 12909 4573 12943 4607
rect 16497 4573 16531 4607
rect 16681 4573 16715 4607
rect 13277 4505 13311 4539
rect 2329 4437 2363 4471
rect 7297 4437 7331 4471
rect 7665 4233 7699 4267
rect 9873 4233 9907 4267
rect 12817 4233 12851 4267
rect 7113 4097 7147 4131
rect 8493 4097 8527 4131
rect 10517 4097 10551 4131
rect 12265 4097 12299 4131
rect 12357 4097 12391 4131
rect 13645 4097 13679 4131
rect 7297 4029 7331 4063
rect 8125 4029 8159 4063
rect 8677 4029 8711 4063
rect 9229 4029 9263 4063
rect 12449 4029 12483 4063
rect 13277 4029 13311 4063
rect 13829 4029 13863 4063
rect 15025 4029 15059 4063
rect 7205 3961 7239 3995
rect 10333 3961 10367 3995
rect 14289 3961 14323 3995
rect 14473 3961 14507 3995
rect 9413 3893 9447 3927
rect 10241 3893 10275 3927
rect 15117 3893 15151 3927
rect 7481 3689 7515 3723
rect 8309 3689 8343 3723
rect 10977 3689 11011 3723
rect 11529 3689 11563 3723
rect 13277 3689 13311 3723
rect 7297 3621 7331 3655
rect 11621 3621 11655 3655
rect 1409 3553 1443 3587
rect 4353 3553 4387 3587
rect 6377 3553 6411 3587
rect 9689 3553 9723 3587
rect 12633 3553 12667 3587
rect 13461 3553 13495 3587
rect 15117 3553 15151 3587
rect 17601 3553 17635 3587
rect 18337 3553 18371 3587
rect 6101 3485 6135 3519
rect 7941 3485 7975 3519
rect 10609 3485 10643 3519
rect 12265 3485 12299 3519
rect 14749 3485 14783 3519
rect 15577 3485 15611 3519
rect 15853 3485 15887 3519
rect 8309 3417 8343 3451
rect 9505 3417 9539 3451
rect 10977 3417 11011 3451
rect 1593 3349 1627 3383
rect 12265 3349 12299 3383
rect 15117 3349 15151 3383
rect 18153 3349 18187 3383
rect 8401 3145 8435 3179
rect 10517 3145 10551 3179
rect 11069 3145 11103 3179
rect 12081 3145 12115 3179
rect 13369 3145 13403 3179
rect 17325 3145 17359 3179
rect 18153 3145 18187 3179
rect 9505 3077 9539 3111
rect 3065 3009 3099 3043
rect 3341 3009 3375 3043
rect 16405 3009 16439 3043
rect 1409 2941 1443 2975
rect 5089 2941 5123 2975
rect 6929 2941 6963 2975
rect 7849 2941 7883 2975
rect 8401 2941 8435 2975
rect 9965 2941 9999 2975
rect 10517 2941 10551 2975
rect 12081 2941 12115 2975
rect 12633 2941 12667 2975
rect 13369 2941 13403 2975
rect 13921 2941 13955 2975
rect 17509 2941 17543 2975
rect 18337 2941 18371 2975
rect 9321 2873 9355 2907
rect 11161 2873 11195 2907
rect 16129 2873 16163 2907
rect 1593 2805 1627 2839
rect 7113 2805 7147 2839
rect 14381 2805 14415 2839
rect 3341 2601 3375 2635
rect 4813 2601 4847 2635
rect 5825 2601 5859 2635
rect 7665 2601 7699 2635
rect 8125 2601 8159 2635
rect 9965 2601 9999 2635
rect 10333 2601 10367 2635
rect 10885 2601 10919 2635
rect 12633 2601 12667 2635
rect 14933 2601 14967 2635
rect 15393 2601 15427 2635
rect 2053 2533 2087 2567
rect 16221 2533 16255 2567
rect 18153 2533 18187 2567
rect 3157 2465 3191 2499
rect 4629 2465 4663 2499
rect 6009 2465 6043 2499
rect 7021 2465 7055 2499
rect 8033 2465 8067 2499
rect 10793 2465 10827 2499
rect 12817 2465 12851 2499
rect 13921 2465 13955 2499
rect 15301 2465 15335 2499
rect 8309 2397 8343 2431
rect 9689 2397 9723 2431
rect 9873 2397 9907 2431
rect 13645 2397 13679 2431
rect 15485 2397 15519 2431
rect 16405 2397 16439 2431
rect 1869 2329 1903 2363
rect 7205 2329 7239 2363
rect 17969 2329 18003 2363
<< metal1 >>
rect 1104 20154 19044 20176
rect 1104 20102 6962 20154
rect 7014 20102 7026 20154
rect 7078 20102 7090 20154
rect 7142 20102 7154 20154
rect 7206 20102 12942 20154
rect 12994 20102 13006 20154
rect 13058 20102 13070 20154
rect 13122 20102 13134 20154
rect 13186 20102 19044 20154
rect 1104 20080 19044 20102
rect 1486 20040 1492 20052
rect 1447 20012 1492 20040
rect 1486 20000 1492 20012
rect 1544 20000 1550 20052
rect 7098 19932 7104 19984
rect 7156 19972 7162 19984
rect 7745 19975 7803 19981
rect 7745 19972 7757 19975
rect 7156 19944 7757 19972
rect 7156 19932 7162 19944
rect 7745 19941 7757 19944
rect 7791 19941 7803 19975
rect 7745 19935 7803 19941
rect 8294 19932 8300 19984
rect 8352 19972 8358 19984
rect 18233 19975 18291 19981
rect 8352 19944 10548 19972
rect 8352 19932 8358 19944
rect 1578 19904 1584 19916
rect 1539 19876 1584 19904
rect 1578 19864 1584 19876
rect 1636 19864 1642 19916
rect 2314 19904 2320 19916
rect 2275 19876 2320 19904
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 2958 19864 2964 19916
rect 3016 19904 3022 19916
rect 3145 19907 3203 19913
rect 3145 19904 3157 19907
rect 3016 19876 3157 19904
rect 3016 19864 3022 19876
rect 3145 19873 3157 19876
rect 3191 19873 3203 19907
rect 3145 19867 3203 19873
rect 3694 19864 3700 19916
rect 3752 19904 3758 19916
rect 4249 19907 4307 19913
rect 4249 19904 4261 19907
rect 3752 19876 4261 19904
rect 3752 19864 3758 19876
rect 4249 19873 4261 19876
rect 4295 19873 4307 19907
rect 5534 19904 5540 19916
rect 5495 19876 5540 19904
rect 4249 19867 4307 19873
rect 5534 19864 5540 19876
rect 5592 19864 5598 19916
rect 6914 19904 6920 19916
rect 6875 19876 6920 19904
rect 6914 19864 6920 19876
rect 6972 19864 6978 19916
rect 7374 19864 7380 19916
rect 7432 19904 7438 19916
rect 7561 19907 7619 19913
rect 7561 19904 7573 19907
rect 7432 19876 7573 19904
rect 7432 19864 7438 19876
rect 7561 19873 7573 19876
rect 7607 19873 7619 19907
rect 7834 19904 7840 19916
rect 7795 19876 7840 19904
rect 7561 19867 7619 19873
rect 7834 19864 7840 19876
rect 7892 19864 7898 19916
rect 7975 19907 8033 19913
rect 7975 19873 7987 19907
rect 8021 19904 8033 19907
rect 8202 19904 8208 19916
rect 8021 19876 8208 19904
rect 8021 19873 8033 19876
rect 7975 19867 8033 19873
rect 8202 19864 8208 19876
rect 8260 19864 8266 19916
rect 9674 19864 9680 19916
rect 9732 19904 9738 19916
rect 10520 19913 10548 19944
rect 18233 19941 18245 19975
rect 18279 19972 18291 19975
rect 18874 19972 18880 19984
rect 18279 19944 18880 19972
rect 18279 19941 18291 19944
rect 18233 19935 18291 19941
rect 18874 19932 18880 19944
rect 18932 19932 18938 19984
rect 9861 19907 9919 19913
rect 9861 19904 9873 19907
rect 9732 19876 9873 19904
rect 9732 19864 9738 19876
rect 9861 19873 9873 19876
rect 9907 19873 9919 19907
rect 9861 19867 9919 19873
rect 10505 19907 10563 19913
rect 10505 19873 10517 19907
rect 10551 19873 10563 19907
rect 10505 19867 10563 19873
rect 11514 19864 11520 19916
rect 11572 19904 11578 19916
rect 12437 19907 12495 19913
rect 12437 19904 12449 19907
rect 11572 19876 12449 19904
rect 11572 19864 11578 19876
rect 12437 19873 12449 19876
rect 12483 19873 12495 19907
rect 12437 19867 12495 19873
rect 12802 19864 12808 19916
rect 12860 19904 12866 19916
rect 13081 19907 13139 19913
rect 13081 19904 13093 19907
rect 12860 19876 13093 19904
rect 12860 19864 12866 19876
rect 13081 19873 13093 19876
rect 13127 19873 13139 19907
rect 13081 19867 13139 19873
rect 14274 19864 14280 19916
rect 14332 19904 14338 19916
rect 15105 19907 15163 19913
rect 15105 19904 15117 19907
rect 14332 19876 15117 19904
rect 14332 19864 14338 19876
rect 15105 19873 15117 19876
rect 15151 19873 15163 19907
rect 15105 19867 15163 19873
rect 15654 19864 15660 19916
rect 15712 19904 15718 19916
rect 15841 19907 15899 19913
rect 15841 19904 15853 19907
rect 15712 19876 15853 19904
rect 15712 19864 15718 19876
rect 15841 19873 15853 19876
rect 15887 19873 15899 19907
rect 15841 19867 15899 19873
rect 16482 19864 16488 19916
rect 16540 19904 16546 19916
rect 16669 19907 16727 19913
rect 16669 19904 16681 19907
rect 16540 19876 16681 19904
rect 16540 19864 16546 19876
rect 16669 19873 16681 19876
rect 16715 19873 16727 19907
rect 16669 19867 16727 19873
rect 7101 19771 7159 19777
rect 7101 19737 7113 19771
rect 7147 19768 7159 19771
rect 8570 19768 8576 19780
rect 7147 19740 8576 19768
rect 7147 19737 7159 19740
rect 7101 19731 7159 19737
rect 8570 19728 8576 19740
rect 8628 19728 8634 19780
rect 9677 19771 9735 19777
rect 9677 19737 9689 19771
rect 9723 19768 9735 19771
rect 10686 19768 10692 19780
rect 9723 19740 10692 19768
rect 9723 19737 9735 19740
rect 9677 19731 9735 19737
rect 10686 19728 10692 19740
rect 10744 19728 10750 19780
rect 18046 19768 18052 19780
rect 18007 19740 18052 19768
rect 18046 19728 18052 19740
rect 18104 19728 18110 19780
rect 2501 19703 2559 19709
rect 2501 19669 2513 19703
rect 2547 19700 2559 19703
rect 2682 19700 2688 19712
rect 2547 19672 2688 19700
rect 2547 19669 2559 19672
rect 2501 19663 2559 19669
rect 2682 19660 2688 19672
rect 2740 19660 2746 19712
rect 2961 19703 3019 19709
rect 2961 19669 2973 19703
rect 3007 19700 3019 19703
rect 3142 19700 3148 19712
rect 3007 19672 3148 19700
rect 3007 19669 3019 19672
rect 2961 19663 3019 19669
rect 3142 19660 3148 19672
rect 3200 19660 3206 19712
rect 4433 19703 4491 19709
rect 4433 19669 4445 19703
rect 4479 19700 4491 19703
rect 4798 19700 4804 19712
rect 4479 19672 4804 19700
rect 4479 19669 4491 19672
rect 4433 19663 4491 19669
rect 4798 19660 4804 19672
rect 4856 19660 4862 19712
rect 5626 19660 5632 19712
rect 5684 19700 5690 19712
rect 5721 19703 5779 19709
rect 5721 19700 5733 19703
rect 5684 19672 5733 19700
rect 5684 19660 5690 19672
rect 5721 19669 5733 19672
rect 5767 19669 5779 19703
rect 5721 19663 5779 19669
rect 8018 19660 8024 19712
rect 8076 19700 8082 19712
rect 8113 19703 8171 19709
rect 8113 19700 8125 19703
rect 8076 19672 8125 19700
rect 8076 19660 8082 19672
rect 8113 19669 8125 19672
rect 8159 19669 8171 19703
rect 10318 19700 10324 19712
rect 10279 19672 10324 19700
rect 8113 19663 8171 19669
rect 10318 19660 10324 19672
rect 10376 19660 10382 19712
rect 11238 19660 11244 19712
rect 11296 19700 11302 19712
rect 12253 19703 12311 19709
rect 12253 19700 12265 19703
rect 11296 19672 12265 19700
rect 11296 19660 11302 19672
rect 12253 19669 12265 19672
rect 12299 19669 12311 19703
rect 12253 19663 12311 19669
rect 12710 19660 12716 19712
rect 12768 19700 12774 19712
rect 12897 19703 12955 19709
rect 12897 19700 12909 19703
rect 12768 19672 12909 19700
rect 12768 19660 12774 19672
rect 12897 19669 12909 19672
rect 12943 19669 12955 19703
rect 12897 19663 12955 19669
rect 14366 19660 14372 19712
rect 14424 19700 14430 19712
rect 14921 19703 14979 19709
rect 14921 19700 14933 19703
rect 14424 19672 14933 19700
rect 14424 19660 14430 19672
rect 14921 19669 14933 19672
rect 14967 19669 14979 19703
rect 14921 19663 14979 19669
rect 15286 19660 15292 19712
rect 15344 19700 15350 19712
rect 15657 19703 15715 19709
rect 15657 19700 15669 19703
rect 15344 19672 15669 19700
rect 15344 19660 15350 19672
rect 15657 19669 15669 19672
rect 15703 19669 15715 19703
rect 16482 19700 16488 19712
rect 16443 19672 16488 19700
rect 15657 19663 15715 19669
rect 16482 19660 16488 19672
rect 16540 19660 16546 19712
rect 1104 19610 19044 19632
rect 1104 19558 3972 19610
rect 4024 19558 4036 19610
rect 4088 19558 4100 19610
rect 4152 19558 4164 19610
rect 4216 19558 9952 19610
rect 10004 19558 10016 19610
rect 10068 19558 10080 19610
rect 10132 19558 10144 19610
rect 10196 19558 15932 19610
rect 15984 19558 15996 19610
rect 16048 19558 16060 19610
rect 16112 19558 16124 19610
rect 16176 19558 19044 19610
rect 1104 19536 19044 19558
rect 1578 19456 1584 19508
rect 1636 19496 1642 19508
rect 1673 19499 1731 19505
rect 1673 19496 1685 19499
rect 1636 19468 1685 19496
rect 1636 19456 1642 19468
rect 1673 19465 1685 19468
rect 1719 19465 1731 19499
rect 1673 19459 1731 19465
rect 2685 19363 2743 19369
rect 2685 19329 2697 19363
rect 2731 19360 2743 19363
rect 3694 19360 3700 19372
rect 2731 19332 3700 19360
rect 2731 19329 2743 19332
rect 2685 19323 2743 19329
rect 3694 19320 3700 19332
rect 3752 19320 3758 19372
rect 7752 19363 7810 19369
rect 7752 19329 7764 19363
rect 7798 19329 7810 19363
rect 8018 19360 8024 19372
rect 7979 19332 8024 19360
rect 7752 19323 7810 19329
rect 1854 19292 1860 19304
rect 1767 19264 1860 19292
rect 1854 19252 1860 19264
rect 1912 19292 1918 19304
rect 2406 19292 2412 19304
rect 1912 19264 2412 19292
rect 1912 19252 1918 19264
rect 2406 19252 2412 19264
rect 2464 19252 2470 19304
rect 3970 19252 3976 19304
rect 4028 19292 4034 19304
rect 5721 19295 5779 19301
rect 5721 19292 5733 19295
rect 4028 19264 5733 19292
rect 4028 19252 4034 19264
rect 5721 19261 5733 19264
rect 5767 19292 5779 19295
rect 5767 19264 7052 19292
rect 5767 19261 5779 19264
rect 5721 19255 5779 19261
rect 934 19184 940 19236
rect 992 19224 998 19236
rect 2958 19224 2964 19236
rect 992 19196 2964 19224
rect 992 19184 998 19196
rect 2958 19184 2964 19196
rect 3016 19184 3022 19236
rect 3326 19184 3332 19236
rect 3384 19184 3390 19236
rect 4157 19159 4215 19165
rect 4157 19125 4169 19159
rect 4203 19156 4215 19159
rect 4522 19156 4528 19168
rect 4203 19128 4528 19156
rect 4203 19125 4215 19128
rect 4157 19119 4215 19125
rect 4522 19116 4528 19128
rect 4580 19116 4586 19168
rect 5902 19156 5908 19168
rect 5863 19128 5908 19156
rect 5902 19116 5908 19128
rect 5960 19116 5966 19168
rect 5994 19116 6000 19168
rect 6052 19156 6058 19168
rect 6917 19159 6975 19165
rect 6917 19156 6929 19159
rect 6052 19128 6929 19156
rect 6052 19116 6058 19128
rect 6917 19125 6929 19128
rect 6963 19125 6975 19159
rect 7024 19156 7052 19264
rect 7098 19252 7104 19304
rect 7156 19292 7162 19304
rect 7156 19264 7201 19292
rect 7156 19252 7162 19264
rect 7558 19252 7564 19304
rect 7616 19292 7622 19304
rect 7760 19292 7788 19323
rect 8018 19320 8024 19332
rect 8076 19320 8082 19372
rect 12636 19332 14320 19360
rect 7616 19264 7788 19292
rect 10413 19295 10471 19301
rect 7616 19252 7622 19264
rect 10413 19261 10425 19295
rect 10459 19292 10471 19295
rect 12636 19292 12664 19332
rect 12802 19292 12808 19304
rect 10459 19264 12664 19292
rect 12763 19264 12808 19292
rect 10459 19261 10471 19264
rect 10413 19255 10471 19261
rect 12802 19252 12808 19264
rect 12860 19252 12866 19304
rect 14292 19292 14320 19332
rect 14918 19292 14924 19304
rect 14292 19264 14924 19292
rect 14918 19252 14924 19264
rect 14976 19292 14982 19304
rect 15289 19295 15347 19301
rect 15289 19292 15301 19295
rect 14976 19264 15301 19292
rect 14976 19252 14982 19264
rect 15289 19261 15301 19264
rect 15335 19292 15347 19295
rect 17497 19295 17555 19301
rect 17497 19292 17509 19295
rect 15335 19264 17509 19292
rect 15335 19261 15347 19264
rect 15289 19255 15347 19261
rect 17497 19261 17509 19264
rect 17543 19261 17555 19295
rect 17497 19255 17555 19261
rect 17586 19252 17592 19304
rect 17644 19292 17650 19304
rect 18141 19295 18199 19301
rect 18141 19292 18153 19295
rect 17644 19264 18153 19292
rect 17644 19252 17650 19264
rect 18141 19261 18153 19264
rect 18187 19261 18199 19295
rect 18141 19255 18199 19261
rect 7285 19227 7343 19233
rect 7285 19193 7297 19227
rect 7331 19224 7343 19227
rect 7374 19224 7380 19236
rect 7331 19196 7380 19224
rect 7331 19193 7343 19196
rect 7285 19187 7343 19193
rect 7374 19184 7380 19196
rect 7432 19224 7438 19236
rect 7432 19196 7604 19224
rect 7432 19184 7438 19196
rect 7466 19156 7472 19168
rect 7024 19128 7472 19156
rect 6917 19119 6975 19125
rect 7466 19116 7472 19128
rect 7524 19116 7530 19168
rect 7576 19156 7604 19196
rect 9030 19184 9036 19236
rect 9088 19184 9094 19236
rect 9674 19184 9680 19236
rect 9732 19224 9738 19236
rect 12820 19224 12848 19252
rect 9732 19196 12848 19224
rect 13081 19227 13139 19233
rect 9732 19184 9738 19196
rect 13081 19193 13093 19227
rect 13127 19193 13139 19227
rect 13081 19187 13139 19193
rect 7742 19156 7748 19168
rect 7576 19128 7748 19156
rect 7742 19116 7748 19128
rect 7800 19116 7806 19168
rect 7834 19116 7840 19168
rect 7892 19156 7898 19168
rect 9493 19159 9551 19165
rect 9493 19156 9505 19159
rect 7892 19128 9505 19156
rect 7892 19116 7898 19128
rect 9493 19125 9505 19128
rect 9539 19125 9551 19159
rect 10594 19156 10600 19168
rect 10555 19128 10600 19156
rect 9493 19119 9551 19125
rect 10594 19116 10600 19128
rect 10652 19116 10658 19168
rect 13096 19156 13124 19187
rect 13814 19184 13820 19236
rect 13872 19184 13878 19236
rect 15746 19184 15752 19236
rect 15804 19224 15810 19236
rect 17770 19224 17776 19236
rect 15804 19196 17776 19224
rect 15804 19184 15810 19196
rect 17770 19184 17776 19196
rect 17828 19224 17834 19236
rect 17828 19196 18000 19224
rect 17828 19184 17834 19196
rect 13262 19156 13268 19168
rect 13096 19128 13268 19156
rect 13262 19116 13268 19128
rect 13320 19116 13326 19168
rect 13446 19116 13452 19168
rect 13504 19156 13510 19168
rect 14553 19159 14611 19165
rect 14553 19156 14565 19159
rect 13504 19128 14565 19156
rect 13504 19116 13510 19128
rect 14553 19125 14565 19128
rect 14599 19125 14611 19159
rect 15470 19156 15476 19168
rect 15431 19128 15476 19156
rect 14553 19119 14611 19125
rect 15470 19116 15476 19128
rect 15528 19116 15534 19168
rect 17310 19156 17316 19168
rect 17271 19128 17316 19156
rect 17310 19116 17316 19128
rect 17368 19116 17374 19168
rect 17972 19165 18000 19196
rect 17957 19159 18015 19165
rect 17957 19125 17969 19159
rect 18003 19125 18015 19159
rect 17957 19119 18015 19125
rect 1104 19066 19044 19088
rect 1104 19014 6962 19066
rect 7014 19014 7026 19066
rect 7078 19014 7090 19066
rect 7142 19014 7154 19066
rect 7206 19014 12942 19066
rect 12994 19014 13006 19066
rect 13058 19014 13070 19066
rect 13122 19014 13134 19066
rect 13186 19014 19044 19066
rect 1104 18992 19044 19014
rect 3326 18952 3332 18964
rect 3287 18924 3332 18952
rect 3326 18912 3332 18924
rect 3384 18912 3390 18964
rect 5994 18952 6000 18964
rect 5276 18924 6000 18952
rect 5276 18893 5304 18924
rect 5994 18912 6000 18924
rect 6052 18912 6058 18964
rect 6733 18955 6791 18961
rect 6733 18921 6745 18955
rect 6779 18952 6791 18955
rect 7282 18952 7288 18964
rect 6779 18924 7288 18952
rect 6779 18921 6791 18924
rect 6733 18915 6791 18921
rect 7282 18912 7288 18924
rect 7340 18912 7346 18964
rect 7834 18912 7840 18964
rect 7892 18952 7898 18964
rect 7892 18924 7972 18952
rect 7892 18912 7898 18924
rect 5261 18887 5319 18893
rect 5261 18853 5273 18887
rect 5307 18853 5319 18887
rect 5261 18847 5319 18853
rect 5902 18844 5908 18896
rect 5960 18844 5966 18896
rect 2774 18776 2780 18828
rect 2832 18816 2838 18828
rect 3145 18819 3203 18825
rect 3145 18816 3157 18819
rect 2832 18788 3157 18816
rect 2832 18776 2838 18788
rect 3145 18785 3157 18788
rect 3191 18816 3203 18819
rect 3970 18816 3976 18828
rect 3191 18788 3976 18816
rect 3191 18785 3203 18788
rect 3145 18779 3203 18785
rect 3970 18776 3976 18788
rect 4028 18776 4034 18828
rect 4433 18819 4491 18825
rect 4433 18785 4445 18819
rect 4479 18816 4491 18819
rect 4522 18816 4528 18828
rect 4479 18788 4528 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 4522 18776 4528 18788
rect 4580 18776 4586 18828
rect 7742 18776 7748 18828
rect 7800 18816 7806 18828
rect 7944 18825 7972 18924
rect 8202 18912 8208 18964
rect 8260 18952 8266 18964
rect 13446 18952 13452 18964
rect 8260 18924 12112 18952
rect 8260 18912 8266 18924
rect 10594 18844 10600 18896
rect 10652 18844 10658 18896
rect 7837 18819 7895 18825
rect 7837 18816 7849 18819
rect 7800 18788 7849 18816
rect 7800 18776 7806 18788
rect 7837 18785 7849 18788
rect 7883 18785 7895 18819
rect 7837 18779 7895 18785
rect 7929 18819 7987 18825
rect 7929 18785 7941 18819
rect 7975 18785 7987 18819
rect 7929 18779 7987 18785
rect 8018 18776 8024 18828
rect 8076 18816 8082 18828
rect 8202 18816 8208 18828
rect 8076 18788 8121 18816
rect 8163 18788 8208 18816
rect 8076 18776 8082 18788
rect 8202 18776 8208 18788
rect 8260 18776 8266 18828
rect 9674 18816 9680 18828
rect 9635 18788 9680 18816
rect 9646 18776 9680 18788
rect 9732 18776 9738 18828
rect 12084 18825 12112 18924
rect 12268 18924 13452 18952
rect 12268 18893 12296 18924
rect 13446 18912 13452 18924
rect 13504 18912 13510 18964
rect 13814 18952 13820 18964
rect 13775 18924 13820 18952
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 12253 18887 12311 18893
rect 12253 18853 12265 18887
rect 12299 18853 12311 18887
rect 12253 18847 12311 18853
rect 12989 18887 13047 18893
rect 12989 18853 13001 18887
rect 13035 18884 13047 18887
rect 13538 18884 13544 18896
rect 13035 18856 13544 18884
rect 13035 18853 13047 18856
rect 12989 18847 13047 18853
rect 13538 18844 13544 18856
rect 13596 18844 13602 18896
rect 14918 18884 14924 18896
rect 13648 18856 14924 18884
rect 12069 18819 12127 18825
rect 12069 18785 12081 18819
rect 12115 18785 12127 18819
rect 12069 18779 12127 18785
rect 2406 18708 2412 18760
rect 2464 18748 2470 18760
rect 4982 18748 4988 18760
rect 2464 18720 4988 18748
rect 2464 18708 2470 18720
rect 4982 18708 4988 18720
rect 5040 18708 5046 18760
rect 6546 18640 6552 18692
rect 6604 18680 6610 18692
rect 7558 18680 7564 18692
rect 6604 18652 7564 18680
rect 6604 18640 6610 18652
rect 7558 18640 7564 18652
rect 7616 18680 7622 18692
rect 9646 18680 9674 18776
rect 9953 18751 10011 18757
rect 9953 18717 9965 18751
rect 9999 18748 10011 18751
rect 12084 18748 12112 18779
rect 12158 18776 12164 18828
rect 12216 18816 12222 18828
rect 12216 18788 12261 18816
rect 12216 18776 12222 18788
rect 12434 18776 12440 18828
rect 12492 18816 12498 18828
rect 12897 18819 12955 18825
rect 12897 18816 12909 18819
rect 12492 18788 12537 18816
rect 12728 18788 12909 18816
rect 12492 18776 12498 18788
rect 12342 18748 12348 18760
rect 9999 18720 11928 18748
rect 12084 18720 12348 18748
rect 9999 18717 10011 18720
rect 9953 18711 10011 18717
rect 11900 18689 11928 18720
rect 12342 18708 12348 18720
rect 12400 18708 12406 18760
rect 12526 18708 12532 18760
rect 12584 18748 12590 18760
rect 12728 18748 12756 18788
rect 12897 18785 12909 18788
rect 12943 18785 12955 18819
rect 13170 18816 13176 18828
rect 13131 18788 13176 18816
rect 12897 18779 12955 18785
rect 13170 18776 13176 18788
rect 13228 18776 13234 18828
rect 13648 18825 13676 18856
rect 14918 18844 14924 18856
rect 14976 18844 14982 18896
rect 15013 18887 15071 18893
rect 15013 18853 15025 18887
rect 15059 18884 15071 18887
rect 15286 18884 15292 18896
rect 15059 18856 15292 18884
rect 15059 18853 15071 18856
rect 15013 18847 15071 18853
rect 15286 18844 15292 18856
rect 15344 18844 15350 18896
rect 15470 18844 15476 18896
rect 15528 18844 15534 18896
rect 16960 18856 17908 18884
rect 13633 18819 13691 18825
rect 13633 18785 13645 18819
rect 13679 18785 13691 18819
rect 13633 18779 13691 18785
rect 16960 18760 16988 18856
rect 17126 18816 17132 18828
rect 17087 18788 17132 18816
rect 17126 18776 17132 18788
rect 17184 18816 17190 18828
rect 17880 18825 17908 18856
rect 17681 18819 17739 18825
rect 17681 18816 17693 18819
rect 17184 18788 17693 18816
rect 17184 18776 17190 18788
rect 17681 18785 17693 18788
rect 17727 18785 17739 18819
rect 17681 18779 17739 18785
rect 17865 18819 17923 18825
rect 17865 18785 17877 18819
rect 17911 18785 17923 18819
rect 17865 18779 17923 18785
rect 12584 18720 12756 18748
rect 12584 18708 12590 18720
rect 12802 18708 12808 18760
rect 12860 18748 12866 18760
rect 14642 18748 14648 18760
rect 12860 18720 14648 18748
rect 12860 18708 12866 18720
rect 14642 18708 14648 18720
rect 14700 18748 14706 18760
rect 14737 18751 14795 18757
rect 14737 18748 14749 18751
rect 14700 18720 14749 18748
rect 14700 18708 14706 18720
rect 14737 18717 14749 18720
rect 14783 18717 14795 18751
rect 16942 18748 16948 18760
rect 16903 18720 16948 18748
rect 14737 18711 14795 18717
rect 16942 18708 16948 18720
rect 17000 18708 17006 18760
rect 7616 18652 9674 18680
rect 11885 18683 11943 18689
rect 7616 18640 7622 18652
rect 11885 18649 11897 18683
rect 11931 18649 11943 18683
rect 11885 18643 11943 18649
rect 13173 18683 13231 18689
rect 13173 18649 13185 18683
rect 13219 18680 13231 18683
rect 13262 18680 13268 18692
rect 13219 18652 13268 18680
rect 13219 18649 13231 18652
rect 13173 18643 13231 18649
rect 13262 18640 13268 18652
rect 13320 18640 13326 18692
rect 4338 18612 4344 18624
rect 4299 18584 4344 18612
rect 4338 18572 4344 18584
rect 4396 18572 4402 18624
rect 7650 18612 7656 18624
rect 7611 18584 7656 18612
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 11425 18615 11483 18621
rect 11425 18581 11437 18615
rect 11471 18612 11483 18615
rect 12158 18612 12164 18624
rect 11471 18584 12164 18612
rect 11471 18581 11483 18584
rect 11425 18575 11483 18581
rect 12158 18572 12164 18584
rect 12216 18572 12222 18624
rect 16298 18572 16304 18624
rect 16356 18612 16362 18624
rect 16485 18615 16543 18621
rect 16485 18612 16497 18615
rect 16356 18584 16497 18612
rect 16356 18572 16362 18584
rect 16485 18581 16497 18584
rect 16531 18581 16543 18615
rect 16485 18575 16543 18581
rect 18141 18615 18199 18621
rect 18141 18581 18153 18615
rect 18187 18612 18199 18615
rect 18230 18612 18236 18624
rect 18187 18584 18236 18612
rect 18187 18581 18199 18584
rect 18141 18575 18199 18581
rect 18230 18572 18236 18584
rect 18288 18572 18294 18624
rect 1104 18522 19044 18544
rect 1104 18470 3972 18522
rect 4024 18470 4036 18522
rect 4088 18470 4100 18522
rect 4152 18470 4164 18522
rect 4216 18470 9952 18522
rect 10004 18470 10016 18522
rect 10068 18470 10080 18522
rect 10132 18470 10144 18522
rect 10196 18470 15932 18522
rect 15984 18470 15996 18522
rect 16048 18470 16060 18522
rect 16112 18470 16124 18522
rect 16176 18470 19044 18522
rect 1104 18448 19044 18470
rect 3694 18408 3700 18420
rect 3655 18380 3700 18408
rect 3694 18368 3700 18380
rect 3752 18368 3758 18420
rect 9030 18408 9036 18420
rect 8991 18380 9036 18408
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 12434 18408 12440 18420
rect 9646 18380 12440 18408
rect 4338 18340 4344 18352
rect 3896 18312 4344 18340
rect 3896 18213 3924 18312
rect 4338 18300 4344 18312
rect 4396 18300 4402 18352
rect 4154 18272 4160 18284
rect 4115 18244 4160 18272
rect 4154 18232 4160 18244
rect 4212 18232 4218 18284
rect 7282 18232 7288 18284
rect 7340 18272 7346 18284
rect 7340 18244 7788 18272
rect 7340 18232 7346 18244
rect 3881 18207 3939 18213
rect 3881 18173 3893 18207
rect 3927 18173 3939 18207
rect 3881 18167 3939 18173
rect 3973 18207 4031 18213
rect 3973 18173 3985 18207
rect 4019 18173 4031 18207
rect 3973 18167 4031 18173
rect 4249 18207 4307 18213
rect 4249 18173 4261 18207
rect 4295 18204 4307 18207
rect 4522 18204 4528 18216
rect 4295 18176 4528 18204
rect 4295 18173 4307 18176
rect 4249 18167 4307 18173
rect 3988 18136 4016 18167
rect 4522 18164 4528 18176
rect 4580 18164 4586 18216
rect 4614 18164 4620 18216
rect 4672 18204 4678 18216
rect 4893 18207 4951 18213
rect 4893 18204 4905 18207
rect 4672 18176 4905 18204
rect 4672 18164 4678 18176
rect 4893 18173 4905 18176
rect 4939 18173 4951 18207
rect 4893 18167 4951 18173
rect 7009 18207 7067 18213
rect 7009 18173 7021 18207
rect 7055 18204 7067 18207
rect 7466 18204 7472 18216
rect 7055 18176 7472 18204
rect 7055 18173 7067 18176
rect 7009 18167 7067 18173
rect 7466 18164 7472 18176
rect 7524 18164 7530 18216
rect 7760 18213 7788 18244
rect 7834 18232 7840 18284
rect 7892 18272 7898 18284
rect 9646 18272 9674 18380
rect 12434 18368 12440 18380
rect 12492 18408 12498 18420
rect 13170 18408 13176 18420
rect 12492 18380 13176 18408
rect 12492 18368 12498 18380
rect 13170 18368 13176 18380
rect 13228 18368 13234 18420
rect 16393 18411 16451 18417
rect 16393 18377 16405 18411
rect 16439 18408 16451 18411
rect 17126 18408 17132 18420
rect 16439 18380 17132 18408
rect 16439 18377 16451 18380
rect 16393 18371 16451 18377
rect 17126 18368 17132 18380
rect 17184 18368 17190 18420
rect 11057 18343 11115 18349
rect 11057 18309 11069 18343
rect 11103 18340 11115 18343
rect 11698 18340 11704 18352
rect 11103 18312 11704 18340
rect 11103 18309 11115 18312
rect 11057 18303 11115 18309
rect 11698 18300 11704 18312
rect 11756 18340 11762 18352
rect 18322 18340 18328 18352
rect 11756 18312 13768 18340
rect 18283 18312 18328 18340
rect 11756 18300 11762 18312
rect 7892 18244 8616 18272
rect 7892 18232 7898 18244
rect 7745 18207 7803 18213
rect 7745 18173 7757 18207
rect 7791 18173 7803 18207
rect 7926 18204 7932 18216
rect 7887 18176 7932 18204
rect 7745 18167 7803 18173
rect 7926 18164 7932 18176
rect 7984 18164 7990 18216
rect 8297 18207 8355 18213
rect 8297 18173 8309 18207
rect 8343 18173 8355 18207
rect 8478 18204 8484 18216
rect 8439 18176 8484 18204
rect 8297 18167 8355 18173
rect 4632 18136 4660 18164
rect 3988 18108 4660 18136
rect 7834 18096 7840 18148
rect 7892 18136 7898 18148
rect 8312 18136 8340 18167
rect 8478 18164 8484 18176
rect 8536 18164 8542 18216
rect 8588 18213 8616 18244
rect 8680 18244 9674 18272
rect 8573 18207 8631 18213
rect 8573 18173 8585 18207
rect 8619 18173 8631 18207
rect 8573 18167 8631 18173
rect 8680 18136 8708 18244
rect 12158 18232 12164 18284
rect 12216 18272 12222 18284
rect 12216 18244 13400 18272
rect 12216 18232 12222 18244
rect 9217 18207 9275 18213
rect 9217 18173 9229 18207
rect 9263 18173 9275 18207
rect 9217 18167 9275 18173
rect 11149 18207 11207 18213
rect 11149 18173 11161 18207
rect 11195 18204 11207 18207
rect 12176 18204 12204 18232
rect 13372 18213 13400 18244
rect 13740 18213 13768 18312
rect 18322 18300 18328 18312
rect 18380 18300 18386 18352
rect 14921 18275 14979 18281
rect 14921 18241 14933 18275
rect 14967 18272 14979 18275
rect 16942 18272 16948 18284
rect 14967 18244 16948 18272
rect 14967 18241 14979 18244
rect 14921 18235 14979 18241
rect 16942 18232 16948 18244
rect 17000 18232 17006 18284
rect 11195 18176 12204 18204
rect 12253 18207 12311 18213
rect 11195 18173 11207 18176
rect 11149 18167 11207 18173
rect 12253 18173 12265 18207
rect 12299 18173 12311 18207
rect 12253 18167 12311 18173
rect 12345 18207 12403 18213
rect 12345 18173 12357 18207
rect 12391 18204 12403 18207
rect 13357 18207 13415 18213
rect 12391 18176 12848 18204
rect 12391 18173 12403 18176
rect 12345 18167 12403 18173
rect 7892 18108 8708 18136
rect 7892 18096 7898 18108
rect 4338 18028 4344 18080
rect 4396 18068 4402 18080
rect 4801 18071 4859 18077
rect 4801 18068 4813 18071
rect 4396 18040 4813 18068
rect 4396 18028 4402 18040
rect 4801 18037 4813 18040
rect 4847 18037 4859 18071
rect 6822 18068 6828 18080
rect 6783 18040 6828 18068
rect 4801 18031 4859 18037
rect 6822 18028 6828 18040
rect 6880 18028 6886 18080
rect 7466 18028 7472 18080
rect 7524 18068 7530 18080
rect 9232 18068 9260 18167
rect 12158 18096 12164 18148
rect 12216 18136 12222 18148
rect 12268 18136 12296 18167
rect 12216 18108 12296 18136
rect 12216 18096 12222 18108
rect 12820 18080 12848 18176
rect 13357 18173 13369 18207
rect 13403 18173 13415 18207
rect 13357 18167 13415 18173
rect 13725 18207 13783 18213
rect 13725 18173 13737 18207
rect 13771 18173 13783 18207
rect 13725 18167 13783 18173
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 14642 18204 14648 18216
rect 14240 18176 14648 18204
rect 14240 18164 14246 18176
rect 14642 18164 14648 18176
rect 14700 18164 14706 18216
rect 13446 18136 13452 18148
rect 13407 18108 13452 18136
rect 13446 18096 13452 18108
rect 13504 18096 13510 18148
rect 13538 18096 13544 18148
rect 13596 18136 13602 18148
rect 17954 18136 17960 18148
rect 13596 18108 13641 18136
rect 16146 18108 17960 18136
rect 13596 18096 13602 18108
rect 17954 18096 17960 18108
rect 18012 18096 18018 18148
rect 18141 18139 18199 18145
rect 18141 18105 18153 18139
rect 18187 18136 18199 18139
rect 18414 18136 18420 18148
rect 18187 18108 18420 18136
rect 18187 18105 18199 18108
rect 18141 18099 18199 18105
rect 18414 18096 18420 18108
rect 18472 18096 18478 18148
rect 7524 18040 9260 18068
rect 7524 18028 7530 18040
rect 11790 18028 11796 18080
rect 11848 18068 11854 18080
rect 12069 18071 12127 18077
rect 12069 18068 12081 18071
rect 11848 18040 12081 18068
rect 11848 18028 11854 18040
rect 12069 18037 12081 18040
rect 12115 18037 12127 18071
rect 12069 18031 12127 18037
rect 12618 18028 12624 18080
rect 12676 18068 12682 18080
rect 12713 18071 12771 18077
rect 12713 18068 12725 18071
rect 12676 18040 12725 18068
rect 12676 18028 12682 18040
rect 12713 18037 12725 18040
rect 12759 18037 12771 18071
rect 12713 18031 12771 18037
rect 12802 18028 12808 18080
rect 12860 18068 12866 18080
rect 13173 18071 13231 18077
rect 13173 18068 13185 18071
rect 12860 18040 13185 18068
rect 12860 18028 12866 18040
rect 13173 18037 13185 18040
rect 13219 18037 13231 18071
rect 13173 18031 13231 18037
rect 1104 17978 19044 18000
rect 1104 17926 6962 17978
rect 7014 17926 7026 17978
rect 7078 17926 7090 17978
rect 7142 17926 7154 17978
rect 7206 17926 12942 17978
rect 12994 17926 13006 17978
rect 13058 17926 13070 17978
rect 13122 17926 13134 17978
rect 13186 17926 19044 17978
rect 1104 17904 19044 17926
rect 4982 17824 4988 17876
rect 5040 17864 5046 17876
rect 6546 17864 6552 17876
rect 5040 17836 6552 17864
rect 5040 17824 5046 17836
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 2774 17688 2780 17740
rect 2832 17728 2838 17740
rect 4433 17731 4491 17737
rect 2832 17700 2877 17728
rect 2832 17688 2838 17700
rect 4433 17697 4445 17731
rect 4479 17728 4491 17731
rect 4522 17728 4528 17740
rect 4479 17700 4528 17728
rect 4479 17697 4491 17700
rect 4433 17691 4491 17697
rect 4522 17688 4528 17700
rect 4580 17688 4586 17740
rect 4617 17731 4675 17737
rect 4617 17697 4629 17731
rect 4663 17728 4675 17731
rect 5442 17728 5448 17740
rect 4663 17700 5448 17728
rect 4663 17697 4675 17700
rect 4617 17691 4675 17697
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 5644 17737 5672 17836
rect 6546 17824 6552 17836
rect 6604 17824 6610 17876
rect 6822 17824 6828 17876
rect 6880 17824 6886 17876
rect 7377 17867 7435 17873
rect 7377 17833 7389 17867
rect 7423 17864 7435 17867
rect 7926 17864 7932 17876
rect 7423 17836 7932 17864
rect 7423 17833 7435 17836
rect 7377 17827 7435 17833
rect 7926 17824 7932 17836
rect 7984 17824 7990 17876
rect 12618 17864 12624 17876
rect 10704 17836 11928 17864
rect 6840 17782 6868 17824
rect 10704 17737 10732 17836
rect 10888 17768 11836 17796
rect 10888 17737 10916 17768
rect 11808 17740 11836 17768
rect 5629 17731 5687 17737
rect 5629 17697 5641 17731
rect 5675 17697 5687 17731
rect 5629 17691 5687 17697
rect 9769 17731 9827 17737
rect 9769 17697 9781 17731
rect 9815 17697 9827 17731
rect 9769 17691 9827 17697
rect 10689 17731 10747 17737
rect 10689 17697 10701 17731
rect 10735 17697 10747 17731
rect 10689 17691 10747 17697
rect 10873 17731 10931 17737
rect 10873 17697 10885 17731
rect 10919 17697 10931 17731
rect 10873 17691 10931 17697
rect 11517 17731 11575 17737
rect 11517 17697 11529 17731
rect 11563 17697 11575 17731
rect 11790 17728 11796 17740
rect 11751 17700 11796 17728
rect 11517 17691 11575 17697
rect 5905 17663 5963 17669
rect 5905 17629 5917 17663
rect 5951 17660 5963 17663
rect 7650 17660 7656 17672
rect 5951 17632 7656 17660
rect 5951 17629 5963 17632
rect 5905 17623 5963 17629
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 9674 17620 9680 17672
rect 9732 17660 9738 17672
rect 9784 17660 9812 17691
rect 11333 17663 11391 17669
rect 11333 17660 11345 17663
rect 9732 17632 11345 17660
rect 9732 17620 9738 17632
rect 11333 17629 11345 17632
rect 11379 17629 11391 17663
rect 11333 17623 11391 17629
rect 1581 17595 1639 17601
rect 1581 17561 1593 17595
rect 1627 17592 1639 17595
rect 11532 17592 11560 17691
rect 11790 17688 11796 17700
rect 11848 17688 11854 17740
rect 11900 17737 11928 17836
rect 12084 17836 12624 17864
rect 12084 17737 12112 17836
rect 12618 17824 12624 17836
rect 12676 17864 12682 17876
rect 12897 17867 12955 17873
rect 12897 17864 12909 17867
rect 12676 17836 12909 17864
rect 12676 17824 12682 17836
rect 12897 17833 12909 17836
rect 12943 17833 12955 17867
rect 12897 17827 12955 17833
rect 16942 17824 16948 17876
rect 17000 17864 17006 17876
rect 17497 17867 17555 17873
rect 17497 17864 17509 17867
rect 17000 17836 17509 17864
rect 17000 17824 17006 17836
rect 17497 17833 17509 17836
rect 17543 17833 17555 17867
rect 17954 17864 17960 17876
rect 17915 17836 17960 17864
rect 17497 17827 17555 17833
rect 17954 17824 17960 17836
rect 18012 17824 18018 17876
rect 12713 17799 12771 17805
rect 12713 17765 12725 17799
rect 12759 17796 12771 17799
rect 12802 17796 12808 17808
rect 12759 17768 12808 17796
rect 12759 17765 12771 17768
rect 12713 17759 12771 17765
rect 12802 17756 12808 17768
rect 12860 17756 12866 17808
rect 16025 17799 16083 17805
rect 16025 17765 16037 17799
rect 16071 17796 16083 17799
rect 16298 17796 16304 17808
rect 16071 17768 16304 17796
rect 16071 17765 16083 17768
rect 16025 17759 16083 17765
rect 16298 17756 16304 17768
rect 16356 17756 16362 17808
rect 17310 17796 17316 17808
rect 17250 17768 17316 17796
rect 17310 17756 17316 17768
rect 17368 17756 17374 17808
rect 11885 17731 11943 17737
rect 11885 17697 11897 17731
rect 11931 17697 11943 17731
rect 11885 17691 11943 17697
rect 12069 17731 12127 17737
rect 12069 17697 12081 17731
rect 12115 17697 12127 17731
rect 12069 17691 12127 17697
rect 11698 17660 11704 17672
rect 11659 17632 11704 17660
rect 11698 17620 11704 17632
rect 11756 17620 11762 17672
rect 11900 17660 11928 17691
rect 12158 17688 12164 17740
rect 12216 17728 12222 17740
rect 12529 17731 12587 17737
rect 12529 17728 12541 17731
rect 12216 17700 12541 17728
rect 12216 17688 12222 17700
rect 12529 17697 12541 17700
rect 12575 17697 12587 17731
rect 12529 17691 12587 17697
rect 13446 17688 13452 17740
rect 13504 17728 13510 17740
rect 13541 17731 13599 17737
rect 13541 17728 13553 17731
rect 13504 17700 13553 17728
rect 13504 17688 13510 17700
rect 13541 17697 13553 17700
rect 13587 17728 13599 17731
rect 14734 17728 14740 17740
rect 13587 17700 14740 17728
rect 13587 17697 13599 17700
rect 13541 17691 13599 17697
rect 14734 17688 14740 17700
rect 14792 17688 14798 17740
rect 14918 17728 14924 17740
rect 14879 17700 14924 17728
rect 14918 17688 14924 17700
rect 14976 17688 14982 17740
rect 18141 17731 18199 17737
rect 18141 17697 18153 17731
rect 18187 17728 18199 17731
rect 18506 17728 18512 17740
rect 18187 17700 18512 17728
rect 18187 17697 18199 17700
rect 18141 17691 18199 17697
rect 18506 17688 18512 17700
rect 18564 17688 18570 17740
rect 12710 17660 12716 17672
rect 11900 17632 12716 17660
rect 12710 17620 12716 17632
rect 12768 17620 12774 17672
rect 14182 17620 14188 17672
rect 14240 17660 14246 17672
rect 15749 17663 15807 17669
rect 15749 17660 15761 17663
rect 14240 17632 15761 17660
rect 14240 17620 14246 17632
rect 15749 17629 15761 17632
rect 15795 17629 15807 17663
rect 15749 17623 15807 17629
rect 13449 17595 13507 17601
rect 13449 17592 13461 17595
rect 1627 17564 4476 17592
rect 11532 17564 13461 17592
rect 1627 17561 1639 17564
rect 1581 17555 1639 17561
rect 2590 17524 2596 17536
rect 2551 17496 2596 17524
rect 2590 17484 2596 17496
rect 2648 17484 2654 17536
rect 3694 17484 3700 17536
rect 3752 17524 3758 17536
rect 4249 17527 4307 17533
rect 4249 17524 4261 17527
rect 3752 17496 4261 17524
rect 3752 17484 3758 17496
rect 4249 17493 4261 17496
rect 4295 17493 4307 17527
rect 4448 17524 4476 17564
rect 13449 17561 13461 17564
rect 13495 17592 13507 17595
rect 13538 17592 13544 17604
rect 13495 17564 13544 17592
rect 13495 17561 13507 17564
rect 13449 17555 13507 17561
rect 13538 17552 13544 17564
rect 13596 17552 13602 17604
rect 5994 17524 6000 17536
rect 4448 17496 6000 17524
rect 4249 17487 4307 17493
rect 5994 17484 6000 17496
rect 6052 17484 6058 17536
rect 9766 17484 9772 17536
rect 9824 17524 9830 17536
rect 9861 17527 9919 17533
rect 9861 17524 9873 17527
rect 9824 17496 9873 17524
rect 9824 17484 9830 17496
rect 9861 17493 9873 17496
rect 9907 17493 9919 17527
rect 9861 17487 9919 17493
rect 10410 17484 10416 17536
rect 10468 17524 10474 17536
rect 10781 17527 10839 17533
rect 10781 17524 10793 17527
rect 10468 17496 10793 17524
rect 10468 17484 10474 17496
rect 10781 17493 10793 17496
rect 10827 17493 10839 17527
rect 10781 17487 10839 17493
rect 14737 17527 14795 17533
rect 14737 17493 14749 17527
rect 14783 17524 14795 17527
rect 14826 17524 14832 17536
rect 14783 17496 14832 17524
rect 14783 17493 14795 17496
rect 14737 17487 14795 17493
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 1104 17434 19044 17456
rect 1104 17382 3972 17434
rect 4024 17382 4036 17434
rect 4088 17382 4100 17434
rect 4152 17382 4164 17434
rect 4216 17382 9952 17434
rect 10004 17382 10016 17434
rect 10068 17382 10080 17434
rect 10132 17382 10144 17434
rect 10196 17382 15932 17434
rect 15984 17382 15996 17434
rect 16048 17382 16060 17434
rect 16112 17382 16124 17434
rect 16176 17382 19044 17434
rect 1104 17360 19044 17382
rect 5442 17320 5448 17332
rect 5403 17292 5448 17320
rect 5442 17280 5448 17292
rect 5500 17280 5506 17332
rect 16025 17323 16083 17329
rect 16025 17320 16037 17323
rect 10060 17292 16037 17320
rect 3329 17255 3387 17261
rect 3329 17221 3341 17255
rect 3375 17252 3387 17255
rect 3375 17224 5304 17252
rect 3375 17221 3387 17224
rect 3329 17215 3387 17221
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17184 1915 17187
rect 3789 17187 3847 17193
rect 3789 17184 3801 17187
rect 1903 17156 3801 17184
rect 1903 17153 1915 17156
rect 1857 17147 1915 17153
rect 3789 17153 3801 17156
rect 3835 17153 3847 17187
rect 3789 17147 3847 17153
rect 1581 17119 1639 17125
rect 1581 17085 1593 17119
rect 1627 17085 1639 17119
rect 1581 17079 1639 17085
rect 1596 17048 1624 17079
rect 3694 17076 3700 17128
rect 3752 17116 3758 17128
rect 3973 17119 4031 17125
rect 3973 17116 3985 17119
rect 3752 17088 3985 17116
rect 3752 17076 3758 17088
rect 3973 17085 3985 17088
rect 4019 17085 4031 17119
rect 3973 17079 4031 17085
rect 1854 17048 1860 17060
rect 1596 17020 1860 17048
rect 1854 17008 1860 17020
rect 1912 17008 1918 17060
rect 2590 17008 2596 17060
rect 2648 17008 2654 17060
rect 4062 17048 4068 17060
rect 4023 17020 4068 17048
rect 4062 17008 4068 17020
rect 4120 17008 4126 17060
rect 4154 17008 4160 17060
rect 4212 17048 4218 17060
rect 4310 17057 4338 17224
rect 4982 17184 4988 17196
rect 4943 17156 4988 17184
rect 4982 17144 4988 17156
rect 5040 17144 5046 17196
rect 4433 17119 4491 17125
rect 4433 17085 4445 17119
rect 4479 17116 4491 17119
rect 4614 17116 4620 17128
rect 4479 17088 4620 17116
rect 4479 17085 4491 17088
rect 4433 17079 4491 17085
rect 4614 17076 4620 17088
rect 4672 17076 4678 17128
rect 4890 17116 4896 17128
rect 4851 17088 4896 17116
rect 4890 17076 4896 17088
rect 4948 17076 4954 17128
rect 5166 17116 5172 17128
rect 5127 17088 5172 17116
rect 5166 17076 5172 17088
rect 5224 17076 5230 17128
rect 5276 17125 5304 17224
rect 5460 17184 5488 17280
rect 10060 17252 10088 17292
rect 16025 17289 16037 17292
rect 16071 17289 16083 17323
rect 16025 17283 16083 17289
rect 16761 17323 16819 17329
rect 16761 17289 16773 17323
rect 16807 17320 16819 17323
rect 18049 17323 18107 17329
rect 18049 17320 18061 17323
rect 16807 17292 18061 17320
rect 16807 17289 16819 17292
rect 16761 17283 16819 17289
rect 18049 17289 18061 17292
rect 18095 17289 18107 17323
rect 18049 17283 18107 17289
rect 13446 17252 13452 17264
rect 9968 17224 10088 17252
rect 12544 17224 13452 17252
rect 9674 17184 9680 17196
rect 5460 17156 7052 17184
rect 9635 17156 9680 17184
rect 5261 17119 5319 17125
rect 5261 17085 5273 17119
rect 5307 17116 5319 17119
rect 5442 17116 5448 17128
rect 5307 17088 5448 17116
rect 5307 17085 5319 17088
rect 5261 17079 5319 17085
rect 5442 17076 5448 17088
rect 5500 17076 5506 17128
rect 7024 17125 7052 17156
rect 9674 17144 9680 17156
rect 9732 17144 9738 17196
rect 9858 17184 9864 17196
rect 9819 17156 9864 17184
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 9968 17193 9996 17224
rect 9953 17187 10011 17193
rect 9953 17153 9965 17187
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 10045 17187 10103 17193
rect 10045 17153 10057 17187
rect 10091 17184 10103 17187
rect 10410 17184 10416 17196
rect 10091 17156 10416 17184
rect 10091 17153 10103 17156
rect 10045 17147 10103 17153
rect 10410 17144 10416 17156
rect 10468 17144 10474 17196
rect 10505 17187 10563 17193
rect 10505 17153 10517 17187
rect 10551 17153 10563 17187
rect 10505 17147 10563 17153
rect 6273 17119 6331 17125
rect 6273 17085 6285 17119
rect 6319 17116 6331 17119
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6319 17088 6837 17116
rect 6319 17085 6331 17088
rect 6273 17079 6331 17085
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 7009 17119 7067 17125
rect 7009 17085 7021 17119
rect 7055 17085 7067 17119
rect 7466 17116 7472 17128
rect 7379 17088 7472 17116
rect 7009 17079 7067 17085
rect 7466 17076 7472 17088
rect 7524 17116 7530 17128
rect 7742 17116 7748 17128
rect 7524 17088 7748 17116
rect 7524 17076 7530 17088
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 8478 17076 8484 17128
rect 8536 17116 8542 17128
rect 9585 17119 9643 17125
rect 9585 17116 9597 17119
rect 8536 17088 9597 17116
rect 8536 17076 8542 17088
rect 9585 17085 9597 17088
rect 9631 17085 9643 17119
rect 9876 17116 9904 17144
rect 10520 17116 10548 17147
rect 9876 17088 10548 17116
rect 10689 17119 10747 17125
rect 9585 17079 9643 17085
rect 10689 17085 10701 17119
rect 10735 17085 10747 17119
rect 10689 17079 10747 17085
rect 4295 17051 4353 17057
rect 4212 17020 4257 17048
rect 4212 17008 4218 17020
rect 4295 17017 4307 17051
rect 4341 17017 4353 17051
rect 4295 17011 4353 17017
rect 8294 17008 8300 17060
rect 8352 17048 8358 17060
rect 9401 17051 9459 17057
rect 9401 17048 9413 17051
rect 8352 17020 9413 17048
rect 8352 17008 8358 17020
rect 9401 17017 9413 17020
rect 9447 17017 9459 17051
rect 10704 17048 10732 17079
rect 10778 17076 10784 17128
rect 10836 17116 10842 17128
rect 12342 17116 12348 17128
rect 10836 17088 10881 17116
rect 12303 17088 12348 17116
rect 10836 17076 10842 17088
rect 12342 17076 12348 17088
rect 12400 17076 12406 17128
rect 12544 17125 12572 17224
rect 13446 17212 13452 17224
rect 13504 17212 13510 17264
rect 16114 17212 16120 17264
rect 16172 17252 16178 17264
rect 16850 17252 16856 17264
rect 16172 17224 16856 17252
rect 16172 17212 16178 17224
rect 16850 17212 16856 17224
rect 16908 17252 16914 17264
rect 16908 17224 17724 17252
rect 16908 17212 16914 17224
rect 12630 17187 12688 17193
rect 12630 17153 12642 17187
rect 12676 17184 12688 17187
rect 12802 17184 12808 17196
rect 12676 17156 12808 17184
rect 12676 17153 12688 17156
rect 12630 17147 12688 17153
rect 12802 17144 12808 17156
rect 12860 17144 12866 17196
rect 14458 17144 14464 17196
rect 14516 17184 14522 17196
rect 15289 17187 15347 17193
rect 15289 17184 15301 17187
rect 14516 17156 15301 17184
rect 14516 17144 14522 17156
rect 15289 17153 15301 17156
rect 15335 17153 15347 17187
rect 17218 17184 17224 17196
rect 15289 17147 15347 17153
rect 16316 17156 17224 17184
rect 12529 17119 12587 17125
rect 12529 17085 12541 17119
rect 12575 17085 12587 17119
rect 12710 17116 12716 17128
rect 12671 17088 12716 17116
rect 12529 17079 12587 17085
rect 12710 17076 12716 17088
rect 12768 17076 12774 17128
rect 12897 17119 12955 17125
rect 12897 17085 12909 17119
rect 12943 17116 12955 17119
rect 13354 17116 13360 17128
rect 12943 17088 13360 17116
rect 12943 17085 12955 17088
rect 12897 17079 12955 17085
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 13538 17116 13544 17128
rect 13499 17088 13544 17116
rect 13538 17076 13544 17088
rect 13596 17076 13602 17128
rect 16316 17125 16344 17156
rect 17218 17144 17224 17156
rect 17276 17184 17282 17196
rect 17696 17193 17724 17224
rect 17589 17187 17647 17193
rect 17589 17184 17601 17187
rect 17276 17156 17601 17184
rect 17276 17144 17282 17156
rect 17589 17153 17601 17156
rect 17635 17153 17647 17187
rect 17589 17147 17647 17153
rect 17681 17187 17739 17193
rect 17681 17153 17693 17187
rect 17727 17153 17739 17187
rect 17681 17147 17739 17153
rect 15841 17119 15899 17125
rect 15841 17085 15853 17119
rect 15887 17085 15899 17119
rect 15841 17079 15899 17085
rect 16301 17119 16359 17125
rect 16301 17085 16313 17119
rect 16347 17085 16359 17119
rect 16301 17079 16359 17085
rect 13081 17051 13139 17057
rect 10704 17020 12572 17048
rect 9401 17011 9459 17017
rect 4522 16940 4528 16992
rect 4580 16980 4586 16992
rect 6273 16983 6331 16989
rect 6273 16980 6285 16983
rect 4580 16952 6285 16980
rect 4580 16940 4586 16952
rect 6273 16949 6285 16952
rect 6319 16949 6331 16983
rect 6273 16943 6331 16949
rect 6362 16940 6368 16992
rect 6420 16980 6426 16992
rect 6825 16983 6883 16989
rect 6825 16980 6837 16983
rect 6420 16952 6837 16980
rect 6420 16940 6426 16952
rect 6825 16949 6837 16952
rect 6871 16949 6883 16983
rect 6825 16943 6883 16949
rect 7558 16940 7564 16992
rect 7616 16980 7622 16992
rect 7653 16983 7711 16989
rect 7653 16980 7665 16983
rect 7616 16952 7665 16980
rect 7616 16940 7622 16952
rect 7653 16949 7665 16952
rect 7699 16949 7711 16983
rect 7653 16943 7711 16949
rect 10505 16983 10563 16989
rect 10505 16949 10517 16983
rect 10551 16980 10563 16983
rect 10778 16980 10784 16992
rect 10551 16952 10784 16980
rect 10551 16949 10563 16952
rect 10505 16943 10563 16949
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 12544 16980 12572 17020
rect 13081 17017 13093 17051
rect 13127 17048 13139 17051
rect 13817 17051 13875 17057
rect 13817 17048 13829 17051
rect 13127 17020 13829 17048
rect 13127 17017 13139 17020
rect 13081 17011 13139 17017
rect 13817 17017 13829 17020
rect 13863 17017 13875 17051
rect 13817 17011 13875 17017
rect 14826 17008 14832 17060
rect 14884 17008 14890 17060
rect 15856 17048 15884 17079
rect 16390 17076 16396 17128
rect 16448 17116 16454 17128
rect 17313 17119 17371 17125
rect 17313 17116 17325 17119
rect 16448 17088 17325 17116
rect 16448 17076 16454 17088
rect 17313 17085 17325 17088
rect 17359 17085 17371 17119
rect 17313 17079 17371 17085
rect 17497 17119 17555 17125
rect 17497 17085 17509 17119
rect 17543 17116 17555 17119
rect 17543 17088 17724 17116
rect 17543 17085 17555 17088
rect 17497 17079 17555 17085
rect 17696 17060 17724 17088
rect 17770 17076 17776 17128
rect 17828 17125 17834 17128
rect 17828 17119 17877 17125
rect 17828 17085 17831 17119
rect 17865 17085 17877 17119
rect 17828 17079 17877 17085
rect 17828 17076 17834 17079
rect 16761 17051 16819 17057
rect 16761 17048 16773 17051
rect 15856 17020 16773 17048
rect 15856 16980 15884 17020
rect 16761 17017 16773 17020
rect 16807 17017 16819 17051
rect 16761 17011 16819 17017
rect 17678 17008 17684 17060
rect 17736 17008 17742 17060
rect 12544 16952 15884 16980
rect 16209 16983 16267 16989
rect 16209 16949 16221 16983
rect 16255 16980 16267 16983
rect 17696 16980 17724 17008
rect 16255 16952 17724 16980
rect 16255 16949 16267 16952
rect 16209 16943 16267 16949
rect 1104 16890 19044 16912
rect 1104 16838 6962 16890
rect 7014 16838 7026 16890
rect 7078 16838 7090 16890
rect 7142 16838 7154 16890
rect 7206 16838 12942 16890
rect 12994 16838 13006 16890
rect 13058 16838 13070 16890
rect 13122 16838 13134 16890
rect 13186 16838 19044 16890
rect 1104 16816 19044 16838
rect 5166 16736 5172 16788
rect 5224 16776 5230 16788
rect 5810 16776 5816 16788
rect 5224 16748 5816 16776
rect 5224 16736 5230 16748
rect 5810 16736 5816 16748
rect 5868 16736 5874 16788
rect 6822 16736 6828 16788
rect 6880 16776 6886 16788
rect 6880 16748 9536 16776
rect 6880 16736 6886 16748
rect 4890 16668 4896 16720
rect 4948 16708 4954 16720
rect 5537 16711 5595 16717
rect 5537 16708 5549 16711
rect 4948 16680 5549 16708
rect 4948 16668 4954 16680
rect 5000 16649 5028 16680
rect 5537 16677 5549 16680
rect 5583 16677 5595 16711
rect 5537 16671 5595 16677
rect 7558 16668 7564 16720
rect 7616 16668 7622 16720
rect 9508 16717 9536 16748
rect 12802 16736 12808 16788
rect 12860 16776 12866 16788
rect 13357 16779 13415 16785
rect 13357 16776 13369 16779
rect 12860 16748 13369 16776
rect 12860 16736 12866 16748
rect 13357 16745 13369 16748
rect 13403 16745 13415 16779
rect 13357 16739 13415 16745
rect 13538 16736 13544 16788
rect 13596 16776 13602 16788
rect 14182 16776 14188 16788
rect 13596 16748 14188 16776
rect 13596 16736 13602 16748
rect 14182 16736 14188 16748
rect 14240 16736 14246 16788
rect 15378 16776 15384 16788
rect 15339 16748 15384 16776
rect 15378 16736 15384 16748
rect 15436 16736 15442 16788
rect 16025 16779 16083 16785
rect 16025 16745 16037 16779
rect 16071 16776 16083 16779
rect 16390 16776 16396 16788
rect 16071 16748 16396 16776
rect 16071 16745 16083 16748
rect 16025 16739 16083 16745
rect 9493 16711 9551 16717
rect 9493 16677 9505 16711
rect 9539 16677 9551 16711
rect 10410 16708 10416 16720
rect 9493 16671 9551 16677
rect 10244 16680 10416 16708
rect 4985 16643 5043 16649
rect 4985 16609 4997 16643
rect 5031 16609 5043 16643
rect 5442 16640 5448 16652
rect 5403 16612 5448 16640
rect 4985 16603 5043 16609
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 9766 16600 9772 16652
rect 9824 16640 9830 16652
rect 10244 16649 10272 16680
rect 10410 16668 10416 16680
rect 10468 16668 10474 16720
rect 12710 16668 12716 16720
rect 12768 16708 12774 16720
rect 16040 16708 16068 16739
rect 16390 16736 16396 16748
rect 16448 16736 16454 16788
rect 18138 16708 18144 16720
rect 12768 16680 13584 16708
rect 12768 16668 12774 16680
rect 9953 16643 10011 16649
rect 9953 16640 9965 16643
rect 9824 16612 9965 16640
rect 9824 16600 9830 16612
rect 9953 16609 9965 16612
rect 9999 16609 10011 16643
rect 9953 16603 10011 16609
rect 10229 16643 10287 16649
rect 10229 16609 10241 16643
rect 10275 16609 10287 16643
rect 10229 16603 10287 16609
rect 10321 16643 10379 16649
rect 10321 16609 10333 16643
rect 10367 16609 10379 16643
rect 10502 16640 10508 16652
rect 10463 16612 10508 16640
rect 10321 16603 10379 16609
rect 4062 16532 4068 16584
rect 4120 16572 4126 16584
rect 4709 16575 4767 16581
rect 4709 16572 4721 16575
rect 4120 16544 4721 16572
rect 4120 16532 4126 16544
rect 4709 16541 4721 16544
rect 4755 16572 4767 16575
rect 6362 16572 6368 16584
rect 4755 16544 6368 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 6362 16532 6368 16544
rect 6420 16532 6426 16584
rect 6546 16572 6552 16584
rect 6507 16544 6552 16572
rect 6546 16532 6552 16544
rect 6604 16532 6610 16584
rect 6825 16575 6883 16581
rect 6825 16541 6837 16575
rect 6871 16572 6883 16575
rect 6914 16572 6920 16584
rect 6871 16544 6920 16572
rect 6871 16541 6883 16544
rect 6825 16535 6883 16541
rect 6914 16532 6920 16544
rect 6972 16532 6978 16584
rect 10336 16572 10364 16603
rect 10502 16600 10508 16612
rect 10560 16600 10566 16652
rect 10778 16640 10784 16652
rect 10739 16612 10784 16640
rect 10778 16600 10784 16612
rect 10836 16600 10842 16652
rect 12069 16643 12127 16649
rect 12069 16609 12081 16643
rect 12115 16609 12127 16643
rect 12069 16603 12127 16609
rect 12253 16643 12311 16649
rect 12253 16609 12265 16643
rect 12299 16640 12311 16643
rect 12342 16640 12348 16652
rect 12299 16612 12348 16640
rect 12299 16609 12311 16612
rect 12253 16603 12311 16609
rect 10410 16572 10416 16584
rect 10336 16544 10416 16572
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 12084 16572 12112 16603
rect 12342 16600 12348 16612
rect 12400 16600 12406 16652
rect 13354 16640 13360 16652
rect 13267 16612 13360 16640
rect 13354 16600 13360 16612
rect 13412 16600 13418 16652
rect 13556 16649 13584 16680
rect 15488 16680 16068 16708
rect 18078 16680 18144 16708
rect 13541 16643 13599 16649
rect 13541 16609 13553 16643
rect 13587 16640 13599 16643
rect 14642 16640 14648 16652
rect 13587 16612 14648 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 14642 16600 14648 16612
rect 14700 16600 14706 16652
rect 15488 16649 15516 16680
rect 18138 16668 18144 16680
rect 18196 16668 18202 16720
rect 15473 16643 15531 16649
rect 15473 16609 15485 16643
rect 15519 16609 15531 16643
rect 15473 16603 15531 16609
rect 15746 16600 15752 16652
rect 15804 16640 15810 16652
rect 15933 16643 15991 16649
rect 15933 16640 15945 16643
rect 15804 16612 15945 16640
rect 15804 16600 15810 16612
rect 15933 16609 15945 16612
rect 15979 16609 15991 16643
rect 15933 16603 15991 16609
rect 16114 16600 16120 16652
rect 16172 16640 16178 16652
rect 16172 16612 16217 16640
rect 16172 16600 16178 16612
rect 12158 16572 12164 16584
rect 12071 16544 12164 16572
rect 12158 16532 12164 16544
rect 12216 16572 12222 16584
rect 13372 16572 13400 16600
rect 14458 16572 14464 16584
rect 12216 16544 14464 16572
rect 12216 16532 12222 16544
rect 14458 16532 14464 16544
rect 14516 16532 14522 16584
rect 16577 16575 16635 16581
rect 16577 16541 16589 16575
rect 16623 16541 16635 16575
rect 16577 16535 16635 16541
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16572 16911 16575
rect 16942 16572 16948 16584
rect 16899 16544 16948 16572
rect 16899 16541 16911 16544
rect 16853 16535 16911 16541
rect 4801 16507 4859 16513
rect 4801 16473 4813 16507
rect 4847 16504 4859 16507
rect 5074 16504 5080 16516
rect 4847 16476 5080 16504
rect 4847 16473 4859 16476
rect 4801 16467 4859 16473
rect 5074 16464 5080 16476
rect 5132 16464 5138 16516
rect 14182 16464 14188 16516
rect 14240 16504 14246 16516
rect 16592 16504 16620 16535
rect 16942 16532 16948 16544
rect 17000 16532 17006 16584
rect 14240 16476 16620 16504
rect 14240 16464 14246 16476
rect 4893 16439 4951 16445
rect 4893 16405 4905 16439
rect 4939 16436 4951 16439
rect 4982 16436 4988 16448
rect 4939 16408 4988 16436
rect 4939 16405 4951 16408
rect 4893 16399 4951 16405
rect 4982 16396 4988 16408
rect 5040 16436 5046 16448
rect 5718 16436 5724 16448
rect 5040 16408 5724 16436
rect 5040 16396 5046 16408
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 7834 16396 7840 16448
rect 7892 16436 7898 16448
rect 8297 16439 8355 16445
rect 8297 16436 8309 16439
rect 7892 16408 8309 16436
rect 7892 16396 7898 16408
rect 8297 16405 8309 16408
rect 8343 16405 8355 16439
rect 12250 16436 12256 16448
rect 12211 16408 12256 16436
rect 8297 16399 8355 16405
rect 12250 16396 12256 16408
rect 12308 16396 12314 16448
rect 18322 16436 18328 16448
rect 18283 16408 18328 16436
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 1104 16346 19044 16368
rect 1104 16294 3972 16346
rect 4024 16294 4036 16346
rect 4088 16294 4100 16346
rect 4152 16294 4164 16346
rect 4216 16294 9952 16346
rect 10004 16294 10016 16346
rect 10068 16294 10080 16346
rect 10132 16294 10144 16346
rect 10196 16294 15932 16346
rect 15984 16294 15996 16346
rect 16048 16294 16060 16346
rect 16112 16294 16124 16346
rect 16176 16294 19044 16346
rect 1104 16272 19044 16294
rect 5810 16232 5816 16244
rect 5771 16204 5816 16232
rect 5810 16192 5816 16204
rect 5868 16192 5874 16244
rect 6914 16232 6920 16244
rect 6875 16204 6920 16232
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 8570 16192 8576 16244
rect 8628 16232 8634 16244
rect 9582 16232 9588 16244
rect 8628 16204 9588 16232
rect 8628 16192 8634 16204
rect 9582 16192 9588 16204
rect 9640 16192 9646 16244
rect 14185 16235 14243 16241
rect 14185 16201 14197 16235
rect 14231 16232 14243 16235
rect 14231 16204 15884 16232
rect 14231 16201 14243 16204
rect 14185 16195 14243 16201
rect 10781 16167 10839 16173
rect 10781 16164 10793 16167
rect 9508 16136 10793 16164
rect 9508 16108 9536 16136
rect 10781 16133 10793 16136
rect 10827 16133 10839 16167
rect 15746 16164 15752 16176
rect 10781 16127 10839 16133
rect 14384 16136 15752 16164
rect 1854 16096 1860 16108
rect 1815 16068 1860 16096
rect 1854 16056 1860 16068
rect 1912 16056 1918 16108
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16096 3663 16099
rect 4706 16096 4712 16108
rect 3651 16068 4712 16096
rect 3651 16065 3663 16068
rect 3605 16059 3663 16065
rect 4706 16056 4712 16068
rect 4764 16056 4770 16108
rect 8202 16096 8208 16108
rect 7300 16068 8208 16096
rect 4801 16031 4859 16037
rect 4801 15997 4813 16031
rect 4847 16028 4859 16031
rect 5074 16028 5080 16040
rect 4847 16000 5080 16028
rect 4847 15997 4859 16000
rect 4801 15991 4859 15997
rect 5074 15988 5080 16000
rect 5132 15988 5138 16040
rect 5718 16028 5724 16040
rect 5631 16000 5724 16028
rect 5718 15988 5724 16000
rect 5776 16028 5782 16040
rect 6822 16028 6828 16040
rect 5776 16000 6828 16028
rect 5776 15988 5782 16000
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 7300 16037 7328 16068
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 9490 16096 9496 16108
rect 9403 16068 9496 16096
rect 9490 16056 9496 16068
rect 9548 16056 9554 16108
rect 9858 16056 9864 16108
rect 9916 16096 9922 16108
rect 10137 16099 10195 16105
rect 10137 16096 10149 16099
rect 9916 16068 10149 16096
rect 9916 16056 9922 16068
rect 10137 16065 10149 16068
rect 10183 16065 10195 16099
rect 12526 16096 12532 16108
rect 10137 16059 10195 16065
rect 12084 16068 12532 16096
rect 7101 16031 7159 16037
rect 7101 16028 7113 16031
rect 7024 16000 7113 16028
rect 2133 15963 2191 15969
rect 2133 15929 2145 15963
rect 2179 15929 2191 15963
rect 2133 15923 2191 15929
rect 2148 15892 2176 15923
rect 2866 15920 2872 15972
rect 2924 15920 2930 15972
rect 4982 15960 4988 15972
rect 4943 15932 4988 15960
rect 4982 15920 4988 15932
rect 5040 15920 5046 15972
rect 3510 15892 3516 15904
rect 2148 15864 3516 15892
rect 3510 15852 3516 15864
rect 3568 15852 3574 15904
rect 4430 15852 4436 15904
rect 4488 15892 4494 15904
rect 4617 15895 4675 15901
rect 4617 15892 4629 15895
rect 4488 15864 4629 15892
rect 4488 15852 4494 15864
rect 4617 15861 4629 15864
rect 4663 15861 4675 15895
rect 7024 15892 7052 16000
rect 7101 15997 7113 16000
rect 7147 15997 7159 16031
rect 7101 15991 7159 15997
rect 7285 16031 7343 16037
rect 7285 15997 7297 16031
rect 7331 15997 7343 16031
rect 7285 15991 7343 15997
rect 7561 16031 7619 16037
rect 7561 15997 7573 16031
rect 7607 16028 7619 16031
rect 8294 16028 8300 16040
rect 7607 16000 8300 16028
rect 7607 15997 7619 16000
rect 7561 15991 7619 15997
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 8570 16028 8576 16040
rect 8531 16000 8576 16028
rect 8570 15988 8576 16000
rect 8628 15988 8634 16040
rect 8665 16031 8723 16037
rect 8665 15997 8677 16031
rect 8711 16028 8723 16031
rect 9398 16028 9404 16040
rect 8711 16000 9404 16028
rect 8711 15997 8723 16000
rect 8665 15991 8723 15997
rect 9398 15988 9404 16000
rect 9456 15988 9462 16040
rect 9582 15988 9588 16040
rect 9640 16028 9646 16040
rect 9769 16031 9827 16037
rect 9769 16028 9781 16031
rect 9640 16000 9781 16028
rect 9640 15988 9646 16000
rect 9769 15997 9781 16000
rect 9815 15997 9827 16031
rect 9769 15991 9827 15997
rect 9953 16031 10011 16037
rect 9953 15997 9965 16031
rect 9999 15997 10011 16031
rect 10226 16028 10232 16040
rect 10187 16000 10232 16028
rect 9953 15991 10011 15997
rect 7190 15960 7196 15972
rect 7151 15932 7196 15960
rect 7190 15920 7196 15932
rect 7248 15920 7254 15972
rect 7423 15963 7481 15969
rect 7423 15929 7435 15963
rect 7469 15960 7481 15963
rect 7834 15960 7840 15972
rect 7469 15932 7840 15960
rect 7469 15929 7481 15932
rect 7423 15923 7481 15929
rect 7834 15920 7840 15932
rect 7892 15920 7898 15972
rect 9968 15960 9996 15991
rect 10226 15988 10232 16000
rect 10284 15988 10290 16040
rect 10873 16031 10931 16037
rect 10873 15997 10885 16031
rect 10919 16028 10931 16031
rect 11146 16028 11152 16040
rect 10919 16000 11152 16028
rect 10919 15997 10931 16000
rect 10873 15991 10931 15997
rect 10888 15960 10916 15991
rect 11146 15988 11152 16000
rect 11204 15988 11210 16040
rect 12084 16037 12112 16068
rect 12526 16056 12532 16068
rect 12584 16096 12590 16108
rect 12584 16068 13584 16096
rect 12584 16056 12590 16068
rect 13556 16040 13584 16068
rect 12069 16031 12127 16037
rect 12069 15997 12081 16031
rect 12115 15997 12127 16031
rect 12069 15991 12127 15997
rect 12158 15988 12164 16040
rect 12216 16028 12222 16040
rect 12253 16031 12311 16037
rect 12253 16028 12265 16031
rect 12216 16000 12265 16028
rect 12216 15988 12222 16000
rect 12253 15997 12265 16000
rect 12299 15997 12311 16031
rect 12253 15991 12311 15997
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 12492 16000 12585 16028
rect 12492 15988 12498 16000
rect 13538 15988 13544 16040
rect 13596 16028 13602 16040
rect 14384 16037 14412 16136
rect 15746 16124 15752 16136
rect 15804 16124 15810 16176
rect 15856 16164 15884 16204
rect 17218 16192 17224 16244
rect 17276 16232 17282 16244
rect 17313 16235 17371 16241
rect 17313 16232 17325 16235
rect 17276 16204 17325 16232
rect 17276 16192 17282 16204
rect 17313 16201 17325 16204
rect 17359 16201 17371 16235
rect 17313 16195 17371 16201
rect 17770 16164 17776 16176
rect 15856 16136 17776 16164
rect 17770 16124 17776 16136
rect 17828 16124 17834 16176
rect 14185 16031 14243 16037
rect 14185 16028 14197 16031
rect 13596 16000 14197 16028
rect 13596 15988 13602 16000
rect 14185 15997 14197 16000
rect 14231 16028 14243 16031
rect 14277 16031 14335 16037
rect 14277 16028 14289 16031
rect 14231 16000 14289 16028
rect 14231 15997 14243 16000
rect 14185 15991 14243 15997
rect 14277 15997 14289 16000
rect 14323 15997 14335 16031
rect 14277 15991 14335 15997
rect 14369 16031 14427 16037
rect 14369 15997 14381 16031
rect 14415 15997 14427 16031
rect 14369 15991 14427 15997
rect 14458 15988 14464 16040
rect 14516 16028 14522 16040
rect 14826 16037 14832 16040
rect 14553 16031 14611 16037
rect 14553 16028 14565 16031
rect 14516 16000 14565 16028
rect 14516 15988 14522 16000
rect 14553 15997 14565 16000
rect 14599 15997 14611 16031
rect 14553 15991 14611 15997
rect 14769 16031 14832 16037
rect 14769 15997 14781 16031
rect 14815 15997 14832 16031
rect 14769 15991 14832 15997
rect 14826 15988 14832 15991
rect 14884 15988 14890 16040
rect 14918 15988 14924 16040
rect 14976 16028 14982 16040
rect 15381 16031 15439 16037
rect 15381 16028 15393 16031
rect 14976 16000 15393 16028
rect 14976 15988 14982 16000
rect 15381 15997 15393 16000
rect 15427 15997 15439 16031
rect 16206 16028 16212 16040
rect 16167 16000 16212 16028
rect 15381 15991 15439 15997
rect 16206 15988 16212 16000
rect 16264 15988 16270 16040
rect 17494 16028 17500 16040
rect 17455 16000 17500 16028
rect 17494 15988 17500 16000
rect 17552 15988 17558 16040
rect 17586 15988 17592 16040
rect 17644 16028 17650 16040
rect 17773 16031 17831 16037
rect 17773 16028 17785 16031
rect 17644 16000 17785 16028
rect 17644 15988 17650 16000
rect 17773 15997 17785 16000
rect 17819 15997 17831 16031
rect 17773 15991 17831 15997
rect 12342 15960 12348 15972
rect 9968 15932 10916 15960
rect 12255 15932 12348 15960
rect 12342 15920 12348 15932
rect 12400 15920 12406 15972
rect 12452 15960 12480 15988
rect 13998 15960 14004 15972
rect 12452 15932 14004 15960
rect 13998 15920 14004 15932
rect 14056 15920 14062 15972
rect 14642 15920 14648 15972
rect 14700 15960 14706 15972
rect 14700 15932 14745 15960
rect 14700 15920 14706 15932
rect 7558 15892 7564 15904
rect 7024 15864 7564 15892
rect 4617 15855 4675 15861
rect 7558 15852 7564 15864
rect 7616 15852 7622 15904
rect 11974 15852 11980 15904
rect 12032 15892 12038 15904
rect 12360 15892 12388 15920
rect 12032 15864 12388 15892
rect 12621 15895 12679 15901
rect 12032 15852 12038 15864
rect 12621 15861 12633 15895
rect 12667 15892 12679 15895
rect 13446 15892 13452 15904
rect 12667 15864 13452 15892
rect 12667 15861 12679 15864
rect 12621 15855 12679 15861
rect 13446 15852 13452 15864
rect 13504 15852 13510 15904
rect 14921 15895 14979 15901
rect 14921 15861 14933 15895
rect 14967 15892 14979 15895
rect 15010 15892 15016 15904
rect 14967 15864 15016 15892
rect 14967 15861 14979 15864
rect 14921 15855 14979 15861
rect 15010 15852 15016 15864
rect 15068 15852 15074 15904
rect 15562 15892 15568 15904
rect 15523 15864 15568 15892
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 16393 15895 16451 15901
rect 16393 15861 16405 15895
rect 16439 15892 16451 15895
rect 17034 15892 17040 15904
rect 16439 15864 17040 15892
rect 16439 15861 16451 15864
rect 16393 15855 16451 15861
rect 17034 15852 17040 15864
rect 17092 15852 17098 15904
rect 17402 15852 17408 15904
rect 17460 15892 17466 15904
rect 17681 15895 17739 15901
rect 17681 15892 17693 15895
rect 17460 15864 17693 15892
rect 17460 15852 17466 15864
rect 17681 15861 17693 15864
rect 17727 15861 17739 15895
rect 17681 15855 17739 15861
rect 1104 15802 19044 15824
rect 1104 15750 6962 15802
rect 7014 15750 7026 15802
rect 7078 15750 7090 15802
rect 7142 15750 7154 15802
rect 7206 15750 12942 15802
rect 12994 15750 13006 15802
rect 13058 15750 13070 15802
rect 13122 15750 13134 15802
rect 13186 15750 19044 15802
rect 1104 15728 19044 15750
rect 2866 15648 2872 15700
rect 2924 15688 2930 15700
rect 2961 15691 3019 15697
rect 2961 15688 2973 15691
rect 2924 15660 2973 15688
rect 2924 15648 2930 15660
rect 2961 15657 2973 15660
rect 3007 15657 3019 15691
rect 2961 15651 3019 15657
rect 3510 15648 3516 15700
rect 3568 15688 3574 15700
rect 4249 15691 4307 15697
rect 4249 15688 4261 15691
rect 3568 15660 4261 15688
rect 3568 15648 3574 15660
rect 4249 15657 4261 15660
rect 4295 15657 4307 15691
rect 7558 15688 7564 15700
rect 7519 15660 7564 15688
rect 4249 15651 4307 15657
rect 7558 15648 7564 15660
rect 7616 15648 7622 15700
rect 10045 15691 10103 15697
rect 10045 15657 10057 15691
rect 10091 15688 10103 15691
rect 10502 15688 10508 15700
rect 10091 15660 10508 15688
rect 10091 15657 10103 15660
rect 10045 15651 10103 15657
rect 10502 15648 10508 15660
rect 10560 15648 10566 15700
rect 11333 15691 11391 15697
rect 11333 15657 11345 15691
rect 11379 15688 11391 15691
rect 11974 15688 11980 15700
rect 11379 15660 11980 15688
rect 11379 15657 11391 15660
rect 11333 15651 11391 15657
rect 11974 15648 11980 15660
rect 12032 15648 12038 15700
rect 14090 15688 14096 15700
rect 13004 15660 14096 15688
rect 4522 15620 4528 15632
rect 4435 15592 4528 15620
rect 4522 15580 4528 15592
rect 4580 15620 4586 15632
rect 5353 15623 5411 15629
rect 5353 15620 5365 15623
rect 4580 15592 5365 15620
rect 4580 15580 4586 15592
rect 5353 15589 5365 15592
rect 5399 15589 5411 15623
rect 5534 15620 5540 15632
rect 5447 15592 5540 15620
rect 5353 15583 5411 15589
rect 5534 15580 5540 15592
rect 5592 15620 5598 15632
rect 6273 15623 6331 15629
rect 6273 15620 6285 15623
rect 5592 15592 6285 15620
rect 5592 15580 5598 15592
rect 6273 15589 6285 15592
rect 6319 15589 6331 15623
rect 10226 15620 10232 15632
rect 6273 15583 6331 15589
rect 9692 15592 10232 15620
rect 9692 15564 9720 15592
rect 10226 15580 10232 15592
rect 10284 15580 10290 15632
rect 13004 15606 13032 15660
rect 14090 15648 14096 15660
rect 14148 15688 14154 15700
rect 14918 15688 14924 15700
rect 14148 15660 14924 15688
rect 14148 15648 14154 15660
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 16942 15688 16948 15700
rect 16903 15660 16948 15688
rect 16942 15648 16948 15660
rect 17000 15648 17006 15700
rect 18230 15688 18236 15700
rect 17144 15660 18236 15688
rect 13446 15620 13452 15632
rect 13407 15592 13452 15620
rect 13446 15580 13452 15592
rect 13504 15580 13510 15632
rect 15010 15620 15016 15632
rect 14971 15592 15016 15620
rect 15010 15580 15016 15592
rect 15068 15580 15074 15632
rect 15562 15580 15568 15632
rect 15620 15580 15626 15632
rect 17144 15564 17172 15660
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 17221 15623 17279 15629
rect 17221 15589 17233 15623
rect 17267 15620 17279 15623
rect 17267 15592 18184 15620
rect 17267 15589 17279 15592
rect 17221 15583 17279 15589
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 2774 15512 2780 15564
rect 2832 15552 2838 15564
rect 4430 15552 4436 15564
rect 2832 15524 2877 15552
rect 4391 15524 4436 15552
rect 2832 15512 2838 15524
rect 4430 15512 4436 15524
rect 4488 15512 4494 15564
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15521 4675 15555
rect 4617 15515 4675 15521
rect 4338 15444 4344 15496
rect 4396 15484 4402 15496
rect 4632 15484 4660 15515
rect 4706 15512 4712 15564
rect 4764 15561 4770 15564
rect 4764 15555 4793 15561
rect 4781 15521 4793 15555
rect 4764 15515 4793 15521
rect 4893 15555 4951 15561
rect 4893 15521 4905 15555
rect 4939 15552 4951 15555
rect 5166 15552 5172 15564
rect 4939 15524 5172 15552
rect 4939 15521 4951 15524
rect 4893 15515 4951 15521
rect 4764 15512 4770 15515
rect 4396 15456 4660 15484
rect 4396 15444 4402 15456
rect 4614 15376 4620 15428
rect 4672 15416 4678 15428
rect 4908 15416 4936 15515
rect 5166 15512 5172 15524
rect 5224 15512 5230 15564
rect 5718 15552 5724 15564
rect 5679 15524 5724 15552
rect 5718 15512 5724 15524
rect 5776 15512 5782 15564
rect 6181 15555 6239 15561
rect 6181 15521 6193 15555
rect 6227 15521 6239 15555
rect 6181 15515 6239 15521
rect 7469 15555 7527 15561
rect 7469 15521 7481 15555
rect 7515 15521 7527 15555
rect 7650 15552 7656 15564
rect 7611 15524 7656 15552
rect 7469 15515 7527 15521
rect 5074 15444 5080 15496
rect 5132 15484 5138 15496
rect 6196 15484 6224 15515
rect 5132 15456 6224 15484
rect 7484 15484 7512 15515
rect 7650 15512 7656 15524
rect 7708 15512 7714 15564
rect 9674 15552 9680 15564
rect 9587 15524 9680 15552
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 11392 15555 11450 15561
rect 11392 15521 11404 15555
rect 11438 15552 11450 15555
rect 12158 15552 12164 15564
rect 11438 15524 12164 15552
rect 11438 15521 11450 15524
rect 11392 15515 11450 15521
rect 12158 15512 12164 15524
rect 12216 15512 12222 15564
rect 17126 15552 17132 15564
rect 17039 15524 17132 15552
rect 17126 15512 17132 15524
rect 17184 15512 17190 15564
rect 17313 15555 17371 15561
rect 17313 15521 17325 15555
rect 17359 15521 17371 15555
rect 17313 15515 17371 15521
rect 17497 15555 17555 15561
rect 17497 15521 17509 15555
rect 17543 15552 17555 15555
rect 17770 15552 17776 15564
rect 17543 15524 17776 15552
rect 17543 15521 17555 15524
rect 17497 15515 17555 15521
rect 7926 15484 7932 15496
rect 7484 15456 7932 15484
rect 5132 15444 5138 15456
rect 7926 15444 7932 15456
rect 7984 15444 7990 15496
rect 9398 15444 9404 15496
rect 9456 15484 9462 15496
rect 9769 15487 9827 15493
rect 9769 15484 9781 15487
rect 9456 15456 9781 15484
rect 9456 15444 9462 15456
rect 9769 15453 9781 15456
rect 9815 15453 9827 15487
rect 9769 15447 9827 15453
rect 10873 15487 10931 15493
rect 10873 15453 10885 15487
rect 10919 15484 10931 15487
rect 12250 15484 12256 15496
rect 10919 15456 12256 15484
rect 10919 15453 10931 15456
rect 10873 15447 10931 15453
rect 12250 15444 12256 15456
rect 12308 15444 12314 15496
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 14182 15484 14188 15496
rect 13771 15456 14188 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 14182 15444 14188 15456
rect 14240 15484 14246 15496
rect 14737 15487 14795 15493
rect 14737 15484 14749 15487
rect 14240 15456 14749 15484
rect 14240 15444 14246 15456
rect 14737 15453 14749 15456
rect 14783 15453 14795 15487
rect 17328 15484 17356 15515
rect 17770 15512 17776 15524
rect 17828 15512 17834 15564
rect 18156 15561 18184 15592
rect 18141 15555 18199 15561
rect 18141 15521 18153 15555
rect 18187 15552 18199 15555
rect 18322 15552 18328 15564
rect 18187 15524 18328 15552
rect 18187 15521 18199 15524
rect 18141 15515 18199 15521
rect 18322 15512 18328 15524
rect 18380 15512 18386 15564
rect 14737 15447 14795 15453
rect 16500 15456 17356 15484
rect 4672 15388 4936 15416
rect 11517 15419 11575 15425
rect 4672 15376 4678 15388
rect 11517 15385 11529 15419
rect 11563 15416 11575 15419
rect 12066 15416 12072 15428
rect 11563 15388 12072 15416
rect 11563 15385 11575 15388
rect 11517 15379 11575 15385
rect 12066 15376 12072 15388
rect 12124 15376 12130 15428
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15348 1639 15351
rect 1762 15348 1768 15360
rect 1627 15320 1768 15348
rect 1627 15317 1639 15320
rect 1581 15311 1639 15317
rect 1762 15308 1768 15320
rect 1820 15308 1826 15360
rect 9490 15308 9496 15360
rect 9548 15348 9554 15360
rect 9677 15351 9735 15357
rect 9677 15348 9689 15351
rect 9548 15320 9689 15348
rect 9548 15308 9554 15320
rect 9677 15317 9689 15320
rect 9723 15317 9735 15351
rect 9677 15311 9735 15317
rect 10965 15351 11023 15357
rect 10965 15317 10977 15351
rect 11011 15348 11023 15351
rect 11054 15348 11060 15360
rect 11011 15320 11060 15348
rect 11011 15317 11023 15320
rect 10965 15311 11023 15317
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 11974 15348 11980 15360
rect 11935 15320 11980 15348
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 16298 15308 16304 15360
rect 16356 15348 16362 15360
rect 16500 15357 16528 15456
rect 16485 15351 16543 15357
rect 16485 15348 16497 15351
rect 16356 15320 16497 15348
rect 16356 15308 16362 15320
rect 16485 15317 16497 15320
rect 16531 15317 16543 15351
rect 16485 15311 16543 15317
rect 17586 15308 17592 15360
rect 17644 15348 17650 15360
rect 18049 15351 18107 15357
rect 18049 15348 18061 15351
rect 17644 15320 18061 15348
rect 17644 15308 17650 15320
rect 18049 15317 18061 15320
rect 18095 15317 18107 15351
rect 18049 15311 18107 15317
rect 1104 15258 19044 15280
rect 1104 15206 3972 15258
rect 4024 15206 4036 15258
rect 4088 15206 4100 15258
rect 4152 15206 4164 15258
rect 4216 15206 9952 15258
rect 10004 15206 10016 15258
rect 10068 15206 10080 15258
rect 10132 15206 10144 15258
rect 10196 15206 15932 15258
rect 15984 15206 15996 15258
rect 16048 15206 16060 15258
rect 16112 15206 16124 15258
rect 16176 15206 19044 15258
rect 1104 15184 19044 15206
rect 4709 15147 4767 15153
rect 4709 15113 4721 15147
rect 4755 15144 4767 15147
rect 4982 15144 4988 15156
rect 4755 15116 4988 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 4982 15104 4988 15116
rect 5040 15104 5046 15156
rect 5169 15147 5227 15153
rect 5169 15113 5181 15147
rect 5215 15144 5227 15147
rect 5258 15144 5264 15156
rect 5215 15116 5264 15144
rect 5215 15113 5227 15116
rect 5169 15107 5227 15113
rect 5258 15104 5264 15116
rect 5316 15104 5322 15156
rect 5718 15104 5724 15156
rect 5776 15144 5782 15156
rect 5813 15147 5871 15153
rect 5813 15144 5825 15147
rect 5776 15116 5825 15144
rect 5776 15104 5782 15116
rect 5813 15113 5825 15116
rect 5859 15113 5871 15147
rect 5813 15107 5871 15113
rect 7650 15104 7656 15156
rect 7708 15144 7714 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7708 15116 7849 15144
rect 7708 15104 7714 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 9674 15144 9680 15156
rect 9635 15116 9680 15144
rect 7837 15107 7895 15113
rect 5000 15076 5028 15104
rect 5000 15048 5764 15076
rect 4706 14900 4712 14952
rect 4764 14940 4770 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4764 14912 4905 14940
rect 4764 14900 4770 14912
rect 4893 14909 4905 14912
rect 4939 14909 4951 14943
rect 4893 14903 4951 14909
rect 4985 14943 5043 14949
rect 4985 14909 4997 14943
rect 5031 14909 5043 14943
rect 4985 14903 5043 14909
rect 5000 14872 5028 14903
rect 5074 14900 5080 14952
rect 5132 14940 5138 14952
rect 5736 14949 5764 15048
rect 5810 14968 5816 15020
rect 5868 15008 5874 15020
rect 5868 14980 7696 15008
rect 5868 14968 5874 14980
rect 5261 14943 5319 14949
rect 5261 14940 5273 14943
rect 5132 14912 5273 14940
rect 5132 14900 5138 14912
rect 5261 14909 5273 14912
rect 5307 14909 5319 14943
rect 5261 14903 5319 14909
rect 5721 14943 5779 14949
rect 5721 14909 5733 14943
rect 5767 14909 5779 14943
rect 5721 14903 5779 14909
rect 6822 14900 6828 14952
rect 6880 14940 6886 14952
rect 7668 14949 7696 14980
rect 7285 14943 7343 14949
rect 7285 14940 7297 14943
rect 6880 14912 7297 14940
rect 6880 14900 6886 14912
rect 7285 14909 7297 14912
rect 7331 14909 7343 14943
rect 7285 14903 7343 14909
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14909 7711 14943
rect 7852 14940 7880 15107
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 18138 15144 18144 15156
rect 18099 15116 18144 15144
rect 18138 15104 18144 15116
rect 18196 15104 18202 15156
rect 14458 15076 14464 15088
rect 14419 15048 14464 15076
rect 14458 15036 14464 15048
rect 14516 15036 14522 15088
rect 17494 15036 17500 15088
rect 17552 15076 17558 15088
rect 17589 15079 17647 15085
rect 17589 15076 17601 15079
rect 17552 15048 17601 15076
rect 17552 15036 17558 15048
rect 17589 15045 17601 15048
rect 17635 15045 17647 15079
rect 17589 15039 17647 15045
rect 9861 15011 9919 15017
rect 9861 14977 9873 15011
rect 9907 15008 9919 15011
rect 10321 15011 10379 15017
rect 9907 14980 10272 15008
rect 9907 14977 9919 14980
rect 9861 14971 9919 14977
rect 8110 14940 8116 14952
rect 7852 14912 8116 14940
rect 7653 14903 7711 14909
rect 8110 14900 8116 14912
rect 8168 14940 8174 14952
rect 8297 14943 8355 14949
rect 8297 14940 8309 14943
rect 8168 14912 8309 14940
rect 8168 14900 8174 14912
rect 8297 14909 8309 14912
rect 8343 14909 8355 14943
rect 8297 14903 8355 14909
rect 9953 14943 10011 14949
rect 9953 14909 9965 14943
rect 9999 14909 10011 14943
rect 10244 14940 10272 14980
rect 10321 14977 10333 15011
rect 10367 15008 10379 15011
rect 10410 15008 10416 15020
rect 10367 14980 10416 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 10410 14968 10416 14980
rect 10468 15008 10474 15020
rect 10781 15011 10839 15017
rect 10781 15008 10793 15011
rect 10468 14980 10793 15008
rect 10468 14968 10474 14980
rect 10781 14977 10793 14980
rect 10827 14977 10839 15011
rect 10781 14971 10839 14977
rect 11974 14968 11980 15020
rect 12032 15008 12038 15020
rect 14826 15008 14832 15020
rect 12032 14980 12572 15008
rect 12032 14968 12038 14980
rect 10870 14940 10876 14952
rect 10244 14912 10876 14940
rect 9953 14903 10011 14909
rect 5810 14872 5816 14884
rect 5000 14844 5816 14872
rect 5810 14832 5816 14844
rect 5868 14832 5874 14884
rect 7466 14872 7472 14884
rect 7427 14844 7472 14872
rect 7466 14832 7472 14844
rect 7524 14832 7530 14884
rect 7561 14875 7619 14881
rect 7561 14841 7573 14875
rect 7607 14872 7619 14875
rect 7834 14872 7840 14884
rect 7607 14844 7840 14872
rect 7607 14841 7619 14844
rect 7561 14835 7619 14841
rect 7834 14832 7840 14844
rect 7892 14832 7898 14884
rect 7926 14832 7932 14884
rect 7984 14872 7990 14884
rect 8481 14875 8539 14881
rect 8481 14872 8493 14875
rect 7984 14844 8493 14872
rect 7984 14832 7990 14844
rect 8481 14841 8493 14844
rect 8527 14841 8539 14875
rect 9968 14872 9996 14903
rect 10870 14900 10876 14912
rect 10928 14940 10934 14952
rect 11149 14943 11207 14949
rect 11149 14940 11161 14943
rect 10928 14912 11161 14940
rect 10928 14900 10934 14912
rect 11149 14909 11161 14912
rect 11195 14909 11207 14943
rect 12250 14940 12256 14952
rect 12211 14912 12256 14940
rect 11149 14903 11207 14909
rect 12250 14900 12256 14912
rect 12308 14900 12314 14952
rect 12544 14949 12572 14980
rect 14752 14980 14832 15008
rect 12529 14943 12587 14949
rect 12529 14909 12541 14943
rect 12575 14909 12587 14943
rect 14642 14940 14648 14952
rect 14603 14912 14648 14940
rect 12529 14903 12587 14909
rect 14642 14900 14648 14912
rect 14700 14900 14706 14952
rect 14752 14949 14780 14980
rect 14826 14968 14832 14980
rect 14884 14968 14890 15020
rect 14737 14943 14795 14949
rect 14737 14909 14749 14943
rect 14783 14909 14795 14943
rect 14737 14903 14795 14909
rect 16206 14900 16212 14952
rect 16264 14940 16270 14952
rect 17402 14940 17408 14952
rect 16264 14912 17408 14940
rect 16264 14900 16270 14912
rect 17402 14900 17408 14912
rect 17460 14900 17466 14952
rect 17586 14940 17592 14952
rect 17547 14912 17592 14940
rect 17586 14900 17592 14912
rect 17644 14900 17650 14952
rect 18325 14943 18383 14949
rect 18325 14909 18337 14943
rect 18371 14940 18383 14943
rect 18506 14940 18512 14952
rect 18371 14912 18512 14940
rect 18371 14909 18383 14912
rect 18325 14903 18383 14909
rect 18506 14900 18512 14912
rect 18564 14900 18570 14952
rect 10962 14872 10968 14884
rect 9968 14844 10968 14872
rect 8481 14835 8539 14841
rect 10962 14832 10968 14844
rect 11020 14832 11026 14884
rect 12437 14875 12495 14881
rect 12437 14841 12449 14875
rect 12483 14872 12495 14875
rect 14458 14872 14464 14884
rect 12483 14844 14464 14872
rect 12483 14841 12495 14844
rect 12437 14835 12495 14841
rect 14458 14832 14464 14844
rect 14516 14832 14522 14884
rect 14829 14875 14887 14881
rect 14829 14841 14841 14875
rect 14875 14872 14887 14875
rect 15102 14872 15108 14884
rect 14875 14844 15108 14872
rect 14875 14841 14887 14844
rect 14829 14835 14887 14841
rect 15102 14832 15108 14844
rect 15160 14832 15166 14884
rect 7282 14764 7288 14816
rect 7340 14804 7346 14816
rect 8665 14807 8723 14813
rect 8665 14804 8677 14807
rect 7340 14776 8677 14804
rect 7340 14764 7346 14776
rect 8665 14773 8677 14776
rect 8711 14773 8723 14807
rect 8665 14767 8723 14773
rect 11514 14764 11520 14816
rect 11572 14804 11578 14816
rect 12069 14807 12127 14813
rect 12069 14804 12081 14807
rect 11572 14776 12081 14804
rect 11572 14764 11578 14776
rect 12069 14773 12081 14776
rect 12115 14773 12127 14807
rect 12069 14767 12127 14773
rect 15013 14807 15071 14813
rect 15013 14773 15025 14807
rect 15059 14804 15071 14807
rect 15194 14804 15200 14816
rect 15059 14776 15200 14804
rect 15059 14773 15071 14776
rect 15013 14767 15071 14773
rect 15194 14764 15200 14776
rect 15252 14764 15258 14816
rect 1104 14714 19044 14736
rect 1104 14662 6962 14714
rect 7014 14662 7026 14714
rect 7078 14662 7090 14714
rect 7142 14662 7154 14714
rect 7206 14662 12942 14714
rect 12994 14662 13006 14714
rect 13058 14662 13070 14714
rect 13122 14662 13134 14714
rect 13186 14662 19044 14714
rect 1104 14640 19044 14662
rect 5813 14603 5871 14609
rect 5813 14569 5825 14603
rect 5859 14569 5871 14603
rect 5813 14563 5871 14569
rect 5828 14532 5856 14563
rect 10870 14560 10876 14612
rect 10928 14600 10934 14612
rect 10965 14603 11023 14609
rect 10965 14600 10977 14603
rect 10928 14572 10977 14600
rect 10928 14560 10934 14572
rect 10965 14569 10977 14572
rect 11011 14569 11023 14603
rect 10965 14563 11023 14569
rect 11149 14603 11207 14609
rect 11149 14569 11161 14603
rect 11195 14600 11207 14603
rect 11514 14600 11520 14612
rect 11195 14572 11520 14600
rect 11195 14569 11207 14572
rect 11149 14563 11207 14569
rect 11514 14560 11520 14572
rect 11572 14560 11578 14612
rect 14642 14560 14648 14612
rect 14700 14600 14706 14612
rect 14921 14603 14979 14609
rect 14921 14600 14933 14603
rect 14700 14572 14933 14600
rect 14700 14560 14706 14572
rect 14921 14569 14933 14572
rect 14967 14569 14979 14603
rect 14921 14563 14979 14569
rect 15746 14560 15752 14612
rect 15804 14600 15810 14612
rect 16206 14600 16212 14612
rect 15804 14572 16212 14600
rect 15804 14560 15810 14572
rect 16206 14560 16212 14572
rect 16264 14560 16270 14612
rect 16850 14560 16856 14612
rect 16908 14600 16914 14612
rect 17037 14603 17095 14609
rect 17037 14600 17049 14603
rect 16908 14572 17049 14600
rect 16908 14560 16914 14572
rect 17037 14569 17049 14572
rect 17083 14569 17095 14603
rect 17037 14563 17095 14569
rect 17221 14603 17279 14609
rect 17221 14569 17233 14603
rect 17267 14600 17279 14603
rect 17310 14600 17316 14612
rect 17267 14572 17316 14600
rect 17267 14569 17279 14572
rect 17221 14563 17279 14569
rect 5828 14504 7788 14532
rect 1486 14464 1492 14476
rect 1447 14436 1492 14464
rect 1486 14424 1492 14436
rect 1544 14424 1550 14476
rect 2041 14467 2099 14473
rect 2041 14433 2053 14467
rect 2087 14464 2099 14467
rect 2682 14464 2688 14476
rect 2087 14436 2688 14464
rect 2087 14433 2099 14436
rect 2041 14427 2099 14433
rect 2682 14424 2688 14436
rect 2740 14424 2746 14476
rect 3050 14464 3056 14476
rect 3011 14436 3056 14464
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 4709 14467 4767 14473
rect 4709 14433 4721 14467
rect 4755 14464 4767 14467
rect 5074 14464 5080 14476
rect 4755 14436 5080 14464
rect 4755 14433 4767 14436
rect 4709 14427 4767 14433
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 5169 14467 5227 14473
rect 5169 14433 5181 14467
rect 5215 14464 5227 14467
rect 5258 14464 5264 14476
rect 5215 14436 5264 14464
rect 5215 14433 5227 14436
rect 5169 14427 5227 14433
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 5445 14467 5503 14473
rect 5445 14433 5457 14467
rect 5491 14464 5503 14467
rect 5534 14464 5540 14476
rect 5491 14436 5540 14464
rect 5491 14433 5503 14436
rect 5445 14427 5503 14433
rect 5534 14424 5540 14436
rect 5592 14424 5598 14476
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14464 5687 14467
rect 5718 14464 5724 14476
rect 5675 14436 5724 14464
rect 5675 14433 5687 14436
rect 5629 14427 5687 14433
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 6917 14467 6975 14473
rect 6917 14433 6929 14467
rect 6963 14464 6975 14467
rect 7466 14464 7472 14476
rect 6963 14436 7472 14464
rect 6963 14433 6975 14436
rect 6917 14427 6975 14433
rect 7466 14424 7472 14436
rect 7524 14424 7530 14476
rect 7653 14467 7711 14473
rect 7653 14433 7665 14467
rect 7699 14433 7711 14467
rect 7760 14464 7788 14504
rect 7926 14464 7932 14476
rect 7760 14436 7932 14464
rect 7653 14427 7711 14433
rect 4433 14399 4491 14405
rect 4433 14365 4445 14399
rect 4479 14396 4491 14399
rect 4522 14396 4528 14408
rect 4479 14368 4528 14396
rect 4479 14365 4491 14368
rect 4433 14359 4491 14365
rect 4522 14356 4528 14368
rect 4580 14356 4586 14408
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14396 4675 14399
rect 5276 14396 5304 14424
rect 4663 14368 5304 14396
rect 4663 14365 4675 14368
rect 4617 14359 4675 14365
rect 2041 14331 2099 14337
rect 2041 14297 2053 14331
rect 2087 14328 2099 14331
rect 2866 14328 2872 14340
rect 2087 14300 2872 14328
rect 2087 14297 2099 14300
rect 2041 14291 2099 14297
rect 2866 14288 2872 14300
rect 2924 14288 2930 14340
rect 2590 14220 2596 14272
rect 2648 14260 2654 14272
rect 2961 14263 3019 14269
rect 2961 14260 2973 14263
rect 2648 14232 2973 14260
rect 2648 14220 2654 14232
rect 2961 14229 2973 14232
rect 3007 14229 3019 14263
rect 4522 14260 4528 14272
rect 4483 14232 4528 14260
rect 2961 14223 3019 14229
rect 4522 14220 4528 14232
rect 4580 14220 4586 14272
rect 5276 14260 5304 14368
rect 5353 14399 5411 14405
rect 5353 14365 5365 14399
rect 5399 14396 5411 14399
rect 5810 14396 5816 14408
rect 5399 14368 5816 14396
rect 5399 14365 5411 14368
rect 5353 14359 5411 14365
rect 5810 14356 5816 14368
rect 5868 14356 5874 14408
rect 6822 14356 6828 14408
rect 6880 14396 6886 14408
rect 7009 14399 7067 14405
rect 7009 14396 7021 14399
rect 6880 14368 7021 14396
rect 6880 14356 6886 14368
rect 7009 14365 7021 14368
rect 7055 14365 7067 14399
rect 7009 14359 7067 14365
rect 7193 14399 7251 14405
rect 7193 14365 7205 14399
rect 7239 14396 7251 14399
rect 7282 14396 7288 14408
rect 7239 14368 7288 14396
rect 7239 14365 7251 14368
rect 7193 14359 7251 14365
rect 5534 14328 5540 14340
rect 5495 14300 5540 14328
rect 5534 14288 5540 14300
rect 5592 14288 5598 14340
rect 7024 14328 7052 14359
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 7668 14340 7696 14427
rect 7926 14424 7932 14436
rect 7984 14424 7990 14476
rect 8110 14464 8116 14476
rect 8071 14436 8116 14464
rect 8110 14424 8116 14436
rect 8168 14424 8174 14476
rect 9214 14464 9220 14476
rect 8312 14436 9220 14464
rect 8312 14405 8340 14436
rect 9214 14424 9220 14436
rect 9272 14464 9278 14476
rect 9493 14467 9551 14473
rect 9493 14464 9505 14467
rect 9272 14436 9505 14464
rect 9272 14424 9278 14436
rect 9493 14433 9505 14436
rect 9539 14433 9551 14467
rect 9493 14427 9551 14433
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 11146 14467 11204 14473
rect 11146 14464 11158 14467
rect 11112 14436 11158 14464
rect 11112 14424 11118 14436
rect 11146 14433 11158 14436
rect 11192 14464 11204 14467
rect 11514 14464 11520 14476
rect 11192 14436 11376 14464
rect 11475 14436 11520 14464
rect 11192 14433 11204 14436
rect 11146 14427 11204 14433
rect 7837 14399 7895 14405
rect 7837 14365 7849 14399
rect 7883 14365 7895 14399
rect 7837 14359 7895 14365
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14365 8355 14399
rect 11348 14396 11376 14436
rect 11514 14424 11520 14436
rect 11572 14424 11578 14476
rect 13354 14464 13360 14476
rect 13315 14436 13360 14464
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 15010 14464 15016 14476
rect 14971 14436 15016 14464
rect 15010 14424 15016 14436
rect 15068 14424 15074 14476
rect 16117 14467 16175 14473
rect 16117 14433 16129 14467
rect 16163 14464 16175 14467
rect 16298 14464 16304 14476
rect 16163 14436 16304 14464
rect 16163 14433 16175 14436
rect 16117 14427 16175 14433
rect 16298 14424 16304 14436
rect 16356 14424 16362 14476
rect 16761 14467 16819 14473
rect 16761 14433 16773 14467
rect 16807 14433 16819 14467
rect 16761 14427 16819 14433
rect 16945 14467 17003 14473
rect 16945 14433 16957 14467
rect 16991 14464 17003 14467
rect 17236 14464 17264 14563
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 17678 14560 17684 14612
rect 17736 14600 17742 14612
rect 18141 14603 18199 14609
rect 18141 14600 18153 14603
rect 17736 14572 18153 14600
rect 17736 14560 17742 14572
rect 18141 14569 18153 14572
rect 18187 14569 18199 14603
rect 18141 14563 18199 14569
rect 16991 14436 17264 14464
rect 17313 14467 17371 14473
rect 16991 14433 17003 14436
rect 16945 14427 17003 14433
rect 17313 14433 17325 14467
rect 17359 14464 17371 14467
rect 17494 14464 17500 14476
rect 17359 14436 17500 14464
rect 17359 14433 17371 14436
rect 17313 14427 17371 14433
rect 11609 14399 11667 14405
rect 11609 14396 11621 14399
rect 11348 14368 11621 14396
rect 8297 14359 8355 14365
rect 11609 14365 11621 14368
rect 11655 14396 11667 14399
rect 11698 14396 11704 14408
rect 11655 14368 11704 14396
rect 11655 14365 11667 14368
rect 11609 14359 11667 14365
rect 7650 14328 7656 14340
rect 7024 14300 7656 14328
rect 5442 14260 5448 14272
rect 5276 14232 5448 14260
rect 5442 14220 5448 14232
rect 5500 14260 5506 14272
rect 7024 14260 7052 14300
rect 7650 14288 7656 14300
rect 7708 14288 7714 14340
rect 5500 14232 7052 14260
rect 5500 14220 5506 14232
rect 7098 14220 7104 14272
rect 7156 14260 7162 14272
rect 7852 14260 7880 14359
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 16776 14396 16804 14427
rect 17328 14396 17356 14427
rect 17494 14424 17500 14436
rect 17552 14424 17558 14476
rect 17862 14424 17868 14476
rect 17920 14464 17926 14476
rect 18325 14467 18383 14473
rect 18325 14464 18337 14467
rect 17920 14436 18337 14464
rect 17920 14424 17926 14436
rect 18325 14433 18337 14436
rect 18371 14433 18383 14467
rect 18325 14427 18383 14433
rect 16776 14368 17356 14396
rect 8018 14328 8024 14340
rect 7979 14300 8024 14328
rect 8018 14288 8024 14300
rect 8076 14288 8082 14340
rect 8386 14260 8392 14272
rect 7156 14232 7201 14260
rect 7852 14232 8392 14260
rect 7156 14220 7162 14232
rect 8386 14220 8392 14232
rect 8444 14220 8450 14272
rect 9306 14220 9312 14272
rect 9364 14260 9370 14272
rect 9585 14263 9643 14269
rect 9585 14260 9597 14263
rect 9364 14232 9597 14260
rect 9364 14220 9370 14232
rect 9585 14229 9597 14232
rect 9631 14229 9643 14263
rect 13262 14260 13268 14272
rect 13223 14232 13268 14260
rect 9585 14223 9643 14229
rect 13262 14220 13268 14232
rect 13320 14220 13326 14272
rect 1104 14170 19044 14192
rect 1104 14118 3972 14170
rect 4024 14118 4036 14170
rect 4088 14118 4100 14170
rect 4152 14118 4164 14170
rect 4216 14118 9952 14170
rect 10004 14118 10016 14170
rect 10068 14118 10080 14170
rect 10132 14118 10144 14170
rect 10196 14118 15932 14170
rect 15984 14118 15996 14170
rect 16048 14118 16060 14170
rect 16112 14118 16124 14170
rect 16176 14118 19044 14170
rect 1104 14096 19044 14118
rect 3050 14056 3056 14068
rect 3011 14028 3056 14056
rect 3050 14016 3056 14028
rect 3108 14016 3114 14068
rect 7466 14016 7472 14068
rect 7524 14056 7530 14068
rect 8110 14056 8116 14068
rect 7524 14028 8116 14056
rect 7524 14016 7530 14028
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 10229 14059 10287 14065
rect 10229 14056 10241 14059
rect 8260 14028 10241 14056
rect 8260 14016 8266 14028
rect 10229 14025 10241 14028
rect 10275 14025 10287 14059
rect 10229 14019 10287 14025
rect 11146 14016 11152 14068
rect 11204 14056 11210 14068
rect 12621 14059 12679 14065
rect 12621 14056 12633 14059
rect 11204 14028 12633 14056
rect 11204 14016 11210 14028
rect 12621 14025 12633 14028
rect 12667 14025 12679 14059
rect 12621 14019 12679 14025
rect 1581 13991 1639 13997
rect 1581 13957 1593 13991
rect 1627 13988 1639 13991
rect 1670 13988 1676 14000
rect 1627 13960 1676 13988
rect 1627 13957 1639 13960
rect 1581 13951 1639 13957
rect 1670 13948 1676 13960
rect 1728 13948 1734 14000
rect 5166 13948 5172 14000
rect 5224 13988 5230 14000
rect 9585 13991 9643 13997
rect 5224 13960 7880 13988
rect 5224 13948 5230 13960
rect 2590 13920 2596 13932
rect 2551 13892 2596 13920
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13920 4215 13923
rect 4203 13892 5028 13920
rect 4203 13889 4215 13892
rect 4157 13883 4215 13889
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 1486 13812 1492 13864
rect 1544 13852 1550 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1544 13824 2053 13852
rect 1544 13812 1550 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 2501 13855 2559 13861
rect 2501 13821 2513 13855
rect 2547 13852 2559 13855
rect 2866 13852 2872 13864
rect 2547 13824 2872 13852
rect 2547 13821 2559 13824
rect 2501 13815 2559 13821
rect 2866 13812 2872 13824
rect 2924 13812 2930 13864
rect 3050 13852 3056 13864
rect 3011 13824 3056 13852
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 3234 13812 3240 13864
rect 3292 13852 3298 13864
rect 3421 13855 3479 13861
rect 3421 13852 3433 13855
rect 3292 13824 3433 13852
rect 3292 13812 3298 13824
rect 3421 13821 3433 13824
rect 3467 13821 3479 13855
rect 3421 13815 3479 13821
rect 4249 13855 4307 13861
rect 4249 13821 4261 13855
rect 4295 13852 4307 13855
rect 4522 13852 4528 13864
rect 4295 13824 4528 13852
rect 4295 13821 4307 13824
rect 4249 13815 4307 13821
rect 4522 13812 4528 13824
rect 4580 13852 4586 13864
rect 4847 13855 4905 13861
rect 4847 13852 4859 13855
rect 4580 13824 4859 13852
rect 4580 13812 4586 13824
rect 4847 13821 4859 13824
rect 4893 13821 4905 13855
rect 5000 13852 5028 13892
rect 5368 13861 5396 13960
rect 7742 13920 7748 13932
rect 7392 13892 7748 13920
rect 5205 13855 5263 13861
rect 5205 13852 5217 13855
rect 5000 13824 5217 13852
rect 4847 13815 4905 13821
rect 5205 13821 5217 13824
rect 5251 13821 5263 13855
rect 5205 13815 5263 13821
rect 5353 13855 5411 13861
rect 5353 13821 5365 13855
rect 5399 13821 5411 13855
rect 5353 13815 5411 13821
rect 7098 13812 7104 13864
rect 7156 13861 7162 13864
rect 7156 13855 7205 13861
rect 7156 13821 7159 13855
rect 7193 13852 7205 13855
rect 7392 13852 7420 13892
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 7852 13920 7880 13960
rect 9585 13957 9597 13991
rect 9631 13988 9643 13991
rect 13725 13991 13783 13997
rect 13725 13988 13737 13991
rect 9631 13960 10088 13988
rect 9631 13957 9643 13960
rect 9585 13951 9643 13957
rect 8294 13920 8300 13932
rect 7852 13892 8300 13920
rect 7558 13852 7564 13864
rect 7193 13824 7420 13852
rect 7519 13824 7564 13852
rect 7193 13821 7205 13824
rect 7156 13815 7205 13821
rect 7156 13812 7162 13815
rect 7558 13812 7564 13824
rect 7616 13812 7622 13864
rect 7653 13855 7711 13861
rect 7653 13821 7665 13855
rect 7699 13852 7711 13855
rect 7852 13852 7880 13892
rect 8294 13880 8300 13892
rect 8352 13920 8358 13932
rect 10060 13929 10088 13960
rect 13188 13960 13737 13988
rect 13188 13929 13216 13960
rect 13725 13957 13737 13960
rect 13771 13957 13783 13991
rect 17865 13991 17923 13997
rect 17865 13988 17877 13991
rect 13725 13951 13783 13957
rect 14292 13960 17877 13988
rect 10045 13923 10103 13929
rect 8352 13892 8984 13920
rect 8352 13880 8358 13892
rect 7699 13824 7880 13852
rect 7699 13821 7711 13824
rect 7653 13815 7711 13821
rect 8018 13812 8024 13864
rect 8076 13852 8082 13864
rect 8956 13861 8984 13892
rect 10045 13889 10057 13923
rect 10091 13889 10103 13923
rect 13173 13923 13231 13929
rect 13173 13920 13185 13923
rect 10045 13883 10103 13889
rect 12912 13892 13185 13920
rect 9122 13861 9128 13864
rect 8113 13855 8171 13861
rect 8113 13852 8125 13855
rect 8076 13824 8125 13852
rect 8076 13812 8082 13824
rect 8113 13821 8125 13824
rect 8159 13821 8171 13855
rect 8113 13815 8171 13821
rect 8941 13855 8999 13861
rect 8941 13821 8953 13855
rect 8987 13821 8999 13855
rect 8941 13815 8999 13821
rect 9089 13855 9128 13861
rect 9089 13821 9101 13855
rect 9089 13815 9128 13821
rect 9122 13812 9128 13815
rect 9180 13812 9186 13864
rect 9306 13852 9312 13864
rect 9267 13824 9312 13852
rect 9306 13812 9312 13824
rect 9364 13812 9370 13864
rect 9490 13861 9496 13864
rect 9447 13855 9496 13861
rect 9447 13821 9459 13855
rect 9493 13821 9496 13855
rect 9447 13815 9496 13821
rect 9490 13812 9496 13815
rect 9548 13812 9554 13864
rect 10321 13855 10379 13861
rect 10321 13821 10333 13855
rect 10367 13852 10379 13855
rect 10778 13852 10784 13864
rect 10367 13824 10784 13852
rect 10367 13821 10379 13824
rect 10321 13815 10379 13821
rect 10778 13812 10784 13824
rect 10836 13812 10842 13864
rect 12912 13861 12940 13892
rect 13173 13889 13185 13892
rect 13219 13889 13231 13923
rect 13173 13883 13231 13889
rect 13265 13923 13323 13929
rect 13265 13889 13277 13923
rect 13311 13920 13323 13923
rect 13354 13920 13360 13932
rect 13311 13892 13360 13920
rect 13311 13889 13323 13892
rect 13265 13883 13323 13889
rect 12805 13855 12863 13861
rect 12805 13821 12817 13855
rect 12851 13821 12863 13855
rect 12805 13815 12863 13821
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13821 12955 13855
rect 13280 13852 13308 13883
rect 13354 13880 13360 13892
rect 13412 13920 13418 13932
rect 14292 13920 14320 13960
rect 17865 13957 17877 13960
rect 17911 13957 17923 13991
rect 17865 13951 17923 13957
rect 13412 13892 14320 13920
rect 13412 13880 13418 13892
rect 14458 13880 14464 13932
rect 14516 13920 14522 13932
rect 14737 13923 14795 13929
rect 14737 13920 14749 13923
rect 14516 13892 14749 13920
rect 14516 13880 14522 13892
rect 14737 13889 14749 13892
rect 14783 13889 14795 13923
rect 15102 13920 15108 13932
rect 15063 13892 15108 13920
rect 14737 13883 14795 13889
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 12897 13815 12955 13821
rect 13004 13824 13308 13852
rect 4982 13784 4988 13796
rect 4943 13756 4988 13784
rect 4982 13744 4988 13756
rect 5040 13744 5046 13796
rect 5077 13787 5135 13793
rect 5077 13753 5089 13787
rect 5123 13784 5135 13787
rect 5534 13784 5540 13796
rect 5123 13756 5540 13784
rect 5123 13753 5135 13756
rect 5077 13747 5135 13753
rect 5534 13744 5540 13756
rect 5592 13744 5598 13796
rect 7285 13787 7343 13793
rect 7285 13753 7297 13787
rect 7331 13753 7343 13787
rect 7285 13747 7343 13753
rect 7377 13787 7435 13793
rect 7377 13753 7389 13787
rect 7423 13784 7435 13787
rect 8036 13784 8064 13812
rect 9214 13784 9220 13796
rect 7423 13756 8064 13784
rect 9175 13756 9220 13784
rect 7423 13753 7435 13756
rect 7377 13747 7435 13753
rect 4709 13719 4767 13725
rect 4709 13685 4721 13719
rect 4755 13716 4767 13719
rect 4798 13716 4804 13728
rect 4755 13688 4804 13716
rect 4755 13685 4767 13688
rect 4709 13679 4767 13685
rect 4798 13676 4804 13688
rect 4856 13676 4862 13728
rect 6822 13676 6828 13728
rect 6880 13716 6886 13728
rect 7009 13719 7067 13725
rect 7009 13716 7021 13719
rect 6880 13688 7021 13716
rect 6880 13676 6886 13688
rect 7009 13685 7021 13688
rect 7055 13685 7067 13719
rect 7300 13716 7328 13747
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 12820 13784 12848 13815
rect 13004 13784 13032 13824
rect 13906 13812 13912 13864
rect 13964 13852 13970 13864
rect 14001 13855 14059 13861
rect 14001 13852 14013 13855
rect 13964 13824 14013 13852
rect 13964 13812 13970 13824
rect 14001 13821 14013 13824
rect 14047 13821 14059 13855
rect 14918 13852 14924 13864
rect 14879 13824 14924 13852
rect 14001 13815 14059 13821
rect 14918 13812 14924 13824
rect 14976 13812 14982 13864
rect 15010 13812 15016 13864
rect 15068 13852 15074 13864
rect 15194 13852 15200 13864
rect 15068 13824 15113 13852
rect 15155 13824 15200 13852
rect 15068 13812 15074 13824
rect 15194 13812 15200 13824
rect 15252 13852 15258 13864
rect 16117 13855 16175 13861
rect 16117 13852 16129 13855
rect 15252 13824 16129 13852
rect 15252 13812 15258 13824
rect 16117 13821 16129 13824
rect 16163 13821 16175 13855
rect 16117 13815 16175 13821
rect 16301 13855 16359 13861
rect 16301 13821 16313 13855
rect 16347 13852 16359 13855
rect 16390 13852 16396 13864
rect 16347 13824 16396 13852
rect 16347 13821 16359 13824
rect 16301 13815 16359 13821
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 17310 13852 17316 13864
rect 17271 13824 17316 13852
rect 17310 13812 17316 13824
rect 17368 13812 17374 13864
rect 17494 13852 17500 13864
rect 17455 13824 17500 13852
rect 17494 13812 17500 13824
rect 17552 13812 17558 13864
rect 17678 13852 17684 13864
rect 17639 13824 17684 13852
rect 17678 13812 17684 13824
rect 17736 13812 17742 13864
rect 13722 13784 13728 13796
rect 12820 13756 13032 13784
rect 13683 13756 13728 13784
rect 13722 13744 13728 13756
rect 13780 13744 13786 13796
rect 15930 13784 15936 13796
rect 15891 13756 15936 13784
rect 15930 13744 15936 13756
rect 15988 13744 15994 13796
rect 17586 13784 17592 13796
rect 17547 13756 17592 13784
rect 17586 13744 17592 13756
rect 17644 13744 17650 13796
rect 8205 13719 8263 13725
rect 8205 13716 8217 13719
rect 7300 13688 8217 13716
rect 7009 13679 7067 13685
rect 8205 13685 8217 13688
rect 8251 13685 8263 13719
rect 10042 13716 10048 13728
rect 10003 13688 10048 13716
rect 8205 13679 8263 13685
rect 10042 13676 10048 13688
rect 10100 13676 10106 13728
rect 13814 13676 13820 13728
rect 13872 13716 13878 13728
rect 13909 13719 13967 13725
rect 13909 13716 13921 13719
rect 13872 13688 13921 13716
rect 13872 13676 13878 13688
rect 13909 13685 13921 13688
rect 13955 13685 13967 13719
rect 13909 13679 13967 13685
rect 13998 13676 14004 13728
rect 14056 13716 14062 13728
rect 15102 13716 15108 13728
rect 14056 13688 15108 13716
rect 14056 13676 14062 13688
rect 15102 13676 15108 13688
rect 15160 13716 15166 13728
rect 17126 13716 17132 13728
rect 15160 13688 17132 13716
rect 15160 13676 15166 13688
rect 17126 13676 17132 13688
rect 17184 13676 17190 13728
rect 1104 13626 19044 13648
rect 1104 13574 6962 13626
rect 7014 13574 7026 13626
rect 7078 13574 7090 13626
rect 7142 13574 7154 13626
rect 7206 13574 12942 13626
rect 12994 13574 13006 13626
rect 13058 13574 13070 13626
rect 13122 13574 13134 13626
rect 13186 13574 19044 13626
rect 1104 13552 19044 13574
rect 1486 13512 1492 13524
rect 1447 13484 1492 13512
rect 1486 13472 1492 13484
rect 1544 13472 1550 13524
rect 1949 13515 2007 13521
rect 1949 13481 1961 13515
rect 1995 13512 2007 13515
rect 3142 13512 3148 13524
rect 1995 13484 3148 13512
rect 1995 13481 2007 13484
rect 1949 13475 2007 13481
rect 3142 13472 3148 13484
rect 3200 13472 3206 13524
rect 4982 13472 4988 13524
rect 5040 13512 5046 13524
rect 5629 13515 5687 13521
rect 5629 13512 5641 13515
rect 5040 13484 5641 13512
rect 5040 13472 5046 13484
rect 5629 13481 5641 13484
rect 5675 13481 5687 13515
rect 5629 13475 5687 13481
rect 7558 13472 7564 13524
rect 7616 13512 7622 13524
rect 7837 13515 7895 13521
rect 7837 13512 7849 13515
rect 7616 13484 7849 13512
rect 7616 13472 7622 13484
rect 7837 13481 7849 13484
rect 7883 13481 7895 13515
rect 7837 13475 7895 13481
rect 9122 13472 9128 13524
rect 9180 13512 9186 13524
rect 9585 13515 9643 13521
rect 9585 13512 9597 13515
rect 9180 13484 9597 13512
rect 9180 13472 9186 13484
rect 9585 13481 9597 13484
rect 9631 13481 9643 13515
rect 9585 13475 9643 13481
rect 11698 13472 11704 13524
rect 11756 13512 11762 13524
rect 12529 13515 12587 13521
rect 12529 13512 12541 13515
rect 11756 13484 12541 13512
rect 11756 13472 11762 13484
rect 12529 13481 12541 13484
rect 12575 13481 12587 13515
rect 12529 13475 12587 13481
rect 12713 13515 12771 13521
rect 12713 13481 12725 13515
rect 12759 13481 12771 13515
rect 13722 13512 13728 13524
rect 13683 13484 13728 13512
rect 12713 13475 12771 13481
rect 2777 13447 2835 13453
rect 2777 13413 2789 13447
rect 2823 13444 2835 13447
rect 2958 13444 2964 13456
rect 2823 13416 2964 13444
rect 2823 13413 2835 13416
rect 2777 13407 2835 13413
rect 2958 13404 2964 13416
rect 3016 13404 3022 13456
rect 10042 13404 10048 13456
rect 10100 13444 10106 13456
rect 10413 13447 10471 13453
rect 10413 13444 10425 13447
rect 10100 13416 10425 13444
rect 10100 13404 10106 13416
rect 10413 13413 10425 13416
rect 10459 13413 10471 13447
rect 10413 13407 10471 13413
rect 11422 13404 11428 13456
rect 11480 13404 11486 13456
rect 12728 13444 12756 13475
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 14737 13515 14795 13521
rect 14737 13481 14749 13515
rect 14783 13512 14795 13515
rect 15010 13512 15016 13524
rect 14783 13484 15016 13512
rect 14783 13481 14795 13484
rect 14737 13475 14795 13481
rect 15010 13472 15016 13484
rect 15068 13472 15074 13524
rect 15565 13515 15623 13521
rect 15565 13481 15577 13515
rect 15611 13512 15623 13515
rect 15930 13512 15936 13524
rect 15611 13484 15936 13512
rect 15611 13481 15623 13484
rect 15565 13475 15623 13481
rect 15930 13472 15936 13484
rect 15988 13472 15994 13524
rect 17310 13472 17316 13524
rect 17368 13512 17374 13524
rect 17497 13515 17555 13521
rect 17497 13512 17509 13515
rect 17368 13484 17509 13512
rect 17368 13472 17374 13484
rect 17497 13481 17509 13484
rect 17543 13481 17555 13515
rect 17678 13512 17684 13524
rect 17591 13484 17684 13512
rect 17497 13475 17555 13481
rect 17678 13472 17684 13484
rect 17736 13512 17742 13524
rect 18322 13512 18328 13524
rect 17736 13484 18328 13512
rect 17736 13472 17742 13484
rect 18322 13472 18328 13484
rect 18380 13472 18386 13524
rect 13906 13444 13912 13456
rect 12728 13416 13912 13444
rect 1857 13379 1915 13385
rect 1857 13345 1869 13379
rect 1903 13376 1915 13379
rect 2682 13376 2688 13388
rect 1903 13348 2544 13376
rect 2643 13348 2688 13376
rect 1903 13345 1915 13348
rect 1857 13339 1915 13345
rect 1578 13268 1584 13320
rect 1636 13308 1642 13320
rect 2041 13311 2099 13317
rect 2041 13308 2053 13311
rect 1636 13280 2053 13308
rect 1636 13268 1642 13280
rect 2041 13277 2053 13280
rect 2087 13277 2099 13311
rect 2516 13308 2544 13348
rect 2682 13336 2688 13348
rect 2740 13336 2746 13388
rect 3234 13376 3240 13388
rect 3195 13348 3240 13376
rect 3234 13336 3240 13348
rect 3292 13336 3298 13388
rect 5077 13379 5135 13385
rect 5077 13345 5089 13379
rect 5123 13345 5135 13379
rect 5534 13376 5540 13388
rect 5495 13348 5540 13376
rect 5077 13339 5135 13345
rect 4430 13308 4436 13320
rect 2516 13280 4436 13308
rect 2041 13271 2099 13277
rect 4430 13268 4436 13280
rect 4488 13268 4494 13320
rect 4798 13308 4804 13320
rect 4759 13280 4804 13308
rect 4798 13268 4804 13280
rect 4856 13268 4862 13320
rect 5092 13308 5120 13339
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 7285 13379 7343 13385
rect 7285 13345 7297 13379
rect 7331 13376 7343 13379
rect 7466 13376 7472 13388
rect 7331 13348 7472 13376
rect 7331 13345 7343 13348
rect 7285 13339 7343 13345
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 7742 13376 7748 13388
rect 7703 13348 7748 13376
rect 7742 13336 7748 13348
rect 7800 13336 7806 13388
rect 9490 13376 9496 13388
rect 9451 13348 9496 13376
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 12710 13379 12768 13385
rect 12710 13345 12722 13379
rect 12756 13376 12768 13379
rect 13081 13379 13139 13385
rect 12756 13348 13032 13376
rect 12756 13345 12768 13348
rect 12710 13339 12768 13345
rect 5718 13308 5724 13320
rect 5092 13280 5724 13308
rect 5718 13268 5724 13280
rect 5776 13268 5782 13320
rect 6822 13268 6828 13320
rect 6880 13308 6886 13320
rect 7009 13311 7067 13317
rect 7009 13308 7021 13311
rect 6880 13280 7021 13308
rect 6880 13268 6886 13280
rect 7009 13277 7021 13280
rect 7055 13277 7067 13311
rect 7009 13271 7067 13277
rect 7193 13311 7251 13317
rect 7193 13277 7205 13311
rect 7239 13308 7251 13311
rect 8202 13308 8208 13320
rect 7239 13280 8208 13308
rect 7239 13277 7251 13280
rect 7193 13271 7251 13277
rect 4338 13200 4344 13252
rect 4396 13240 4402 13252
rect 7101 13243 7159 13249
rect 4396 13212 5028 13240
rect 4396 13200 4402 13212
rect 4522 13132 4528 13184
rect 4580 13172 4586 13184
rect 5000 13181 5028 13212
rect 7101 13209 7113 13243
rect 7147 13240 7159 13243
rect 7282 13240 7288 13252
rect 7147 13212 7288 13240
rect 7147 13209 7159 13212
rect 7101 13203 7159 13209
rect 7282 13200 7288 13212
rect 7340 13200 7346 13252
rect 4893 13175 4951 13181
rect 4893 13172 4905 13175
rect 4580 13144 4905 13172
rect 4580 13132 4586 13144
rect 4893 13141 4905 13144
rect 4939 13141 4951 13175
rect 4893 13135 4951 13141
rect 4985 13175 5043 13181
rect 4985 13141 4997 13175
rect 5031 13172 5043 13175
rect 7392 13172 7420 13280
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 10137 13311 10195 13317
rect 10137 13277 10149 13311
rect 10183 13308 10195 13311
rect 10410 13308 10416 13320
rect 10183 13280 10416 13308
rect 10183 13277 10195 13280
rect 10137 13271 10195 13277
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 13004 13240 13032 13348
rect 13081 13345 13093 13379
rect 13127 13376 13139 13379
rect 13262 13376 13268 13388
rect 13127 13348 13268 13376
rect 13127 13345 13139 13348
rect 13081 13339 13139 13345
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 13648 13385 13676 13416
rect 13906 13404 13912 13416
rect 13964 13404 13970 13456
rect 16853 13447 16911 13453
rect 16853 13444 16865 13447
rect 15764 13416 16865 13444
rect 13633 13379 13691 13385
rect 13633 13345 13645 13379
rect 13679 13345 13691 13379
rect 13814 13376 13820 13388
rect 13727 13348 13820 13376
rect 13633 13339 13691 13345
rect 13814 13336 13820 13348
rect 13872 13336 13878 13388
rect 15102 13376 15108 13388
rect 15063 13348 15108 13376
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 15764 13385 15792 13416
rect 16853 13413 16865 13416
rect 16899 13413 16911 13447
rect 16853 13407 16911 13413
rect 15749 13379 15807 13385
rect 15749 13345 15761 13379
rect 15795 13345 15807 13379
rect 15749 13339 15807 13345
rect 13173 13311 13231 13317
rect 13173 13277 13185 13311
rect 13219 13308 13231 13311
rect 13722 13308 13728 13320
rect 13219 13280 13728 13308
rect 13219 13277 13231 13280
rect 13173 13271 13231 13277
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 13832 13240 13860 13336
rect 15010 13308 15016 13320
rect 14923 13280 15016 13308
rect 15010 13268 15016 13280
rect 15068 13308 15074 13320
rect 15764 13308 15792 13339
rect 15838 13336 15844 13388
rect 15896 13376 15902 13388
rect 15933 13379 15991 13385
rect 15933 13376 15945 13379
rect 15896 13348 15945 13376
rect 15896 13336 15902 13348
rect 15933 13345 15945 13348
rect 15979 13345 15991 13379
rect 15933 13339 15991 13345
rect 16117 13379 16175 13385
rect 16117 13345 16129 13379
rect 16163 13345 16175 13379
rect 16117 13339 16175 13345
rect 16301 13379 16359 13385
rect 16301 13345 16313 13379
rect 16347 13376 16359 13379
rect 16945 13379 17003 13385
rect 16347 13348 16528 13376
rect 16347 13345 16359 13348
rect 16301 13339 16359 13345
rect 15068 13280 15792 13308
rect 15068 13268 15074 13280
rect 15746 13240 15752 13252
rect 13004 13212 15752 13240
rect 15746 13200 15752 13212
rect 15804 13200 15810 13252
rect 5031 13144 7420 13172
rect 5031 13141 5043 13144
rect 4985 13135 5043 13141
rect 7834 13132 7840 13184
rect 7892 13172 7898 13184
rect 8202 13172 8208 13184
rect 7892 13144 8208 13172
rect 7892 13132 7898 13144
rect 8202 13132 8208 13144
rect 8260 13132 8266 13184
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 11885 13175 11943 13181
rect 11885 13172 11897 13175
rect 11112 13144 11897 13172
rect 11112 13132 11118 13144
rect 11885 13141 11897 13144
rect 11931 13141 11943 13175
rect 11885 13135 11943 13141
rect 15105 13175 15163 13181
rect 15105 13141 15117 13175
rect 15151 13172 15163 13175
rect 15286 13172 15292 13184
rect 15151 13144 15292 13172
rect 15151 13141 15163 13144
rect 15105 13135 15163 13141
rect 15286 13132 15292 13144
rect 15344 13172 15350 13184
rect 15856 13172 15884 13336
rect 16025 13311 16083 13317
rect 16025 13277 16037 13311
rect 16071 13277 16083 13311
rect 16132 13308 16160 13339
rect 16500 13308 16528 13348
rect 16945 13345 16957 13379
rect 16991 13376 17003 13379
rect 17678 13376 17684 13388
rect 16991 13348 17684 13376
rect 16991 13345 17003 13348
rect 16945 13339 17003 13345
rect 17126 13308 17132 13320
rect 16132 13280 16436 13308
rect 16500 13280 17132 13308
rect 16025 13271 16083 13277
rect 16040 13240 16068 13271
rect 16298 13240 16304 13252
rect 16040 13212 16304 13240
rect 16298 13200 16304 13212
rect 16356 13200 16362 13252
rect 16408 13240 16436 13280
rect 17126 13268 17132 13280
rect 17184 13268 17190 13320
rect 17236 13240 17264 13348
rect 17678 13336 17684 13348
rect 17736 13376 17742 13388
rect 18141 13379 18199 13385
rect 18141 13376 18153 13379
rect 17736 13348 18153 13376
rect 17736 13336 17742 13348
rect 18141 13345 18153 13348
rect 18187 13345 18199 13379
rect 18141 13339 18199 13345
rect 16408 13212 17264 13240
rect 15344 13144 15884 13172
rect 18049 13175 18107 13181
rect 15344 13132 15350 13144
rect 18049 13141 18061 13175
rect 18095 13172 18107 13175
rect 18322 13172 18328 13184
rect 18095 13144 18328 13172
rect 18095 13141 18107 13144
rect 18049 13135 18107 13141
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 1104 13082 19044 13104
rect 1104 13030 3972 13082
rect 4024 13030 4036 13082
rect 4088 13030 4100 13082
rect 4152 13030 4164 13082
rect 4216 13030 9952 13082
rect 10004 13030 10016 13082
rect 10068 13030 10080 13082
rect 10132 13030 10144 13082
rect 10196 13030 15932 13082
rect 15984 13030 15996 13082
rect 16048 13030 16060 13082
rect 16112 13030 16124 13082
rect 16176 13030 19044 13082
rect 1104 13008 19044 13030
rect 3050 12928 3056 12980
rect 3108 12968 3114 12980
rect 3145 12971 3203 12977
rect 3145 12968 3157 12971
rect 3108 12940 3157 12968
rect 3108 12928 3114 12940
rect 3145 12937 3157 12940
rect 3191 12937 3203 12971
rect 3145 12931 3203 12937
rect 5169 12971 5227 12977
rect 5169 12937 5181 12971
rect 5215 12968 5227 12971
rect 5534 12968 5540 12980
rect 5215 12940 5540 12968
rect 5215 12937 5227 12940
rect 5169 12931 5227 12937
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 5629 12971 5687 12977
rect 5629 12937 5641 12971
rect 5675 12968 5687 12971
rect 5902 12968 5908 12980
rect 5675 12940 5908 12968
rect 5675 12937 5687 12940
rect 5629 12931 5687 12937
rect 5902 12928 5908 12940
rect 5960 12968 5966 12980
rect 7558 12968 7564 12980
rect 5960 12940 7564 12968
rect 5960 12928 5966 12940
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 8018 12968 8024 12980
rect 7979 12940 8024 12968
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 14918 12968 14924 12980
rect 14879 12940 14924 12968
rect 14918 12928 14924 12940
rect 14976 12928 14982 12980
rect 15013 12971 15071 12977
rect 15013 12937 15025 12971
rect 15059 12968 15071 12971
rect 15286 12968 15292 12980
rect 15059 12940 15292 12968
rect 15059 12937 15071 12940
rect 15013 12931 15071 12937
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 3234 12860 3240 12912
rect 3292 12900 3298 12912
rect 8941 12903 8999 12909
rect 8941 12900 8953 12903
rect 3292 12872 8953 12900
rect 3292 12860 3298 12872
rect 8941 12869 8953 12872
rect 8987 12869 8999 12903
rect 8941 12863 8999 12869
rect 11057 12903 11115 12909
rect 11057 12869 11069 12903
rect 11103 12900 11115 12903
rect 13538 12900 13544 12912
rect 11103 12872 13544 12900
rect 11103 12869 11115 12872
rect 11057 12863 11115 12869
rect 13538 12860 13544 12872
rect 13596 12860 13602 12912
rect 15102 12860 15108 12912
rect 15160 12860 15166 12912
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12832 9459 12835
rect 9766 12832 9772 12844
rect 9447 12804 9772 12832
rect 9447 12801 9459 12804
rect 9401 12795 9459 12801
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 13906 12832 13912 12844
rect 12820 12804 13912 12832
rect 2682 12724 2688 12776
rect 2740 12764 2746 12776
rect 3142 12764 3148 12776
rect 2740 12736 3148 12764
rect 2740 12724 2746 12736
rect 3142 12724 3148 12736
rect 3200 12764 3206 12776
rect 3329 12767 3387 12773
rect 3329 12764 3341 12767
rect 3200 12736 3341 12764
rect 3200 12724 3206 12736
rect 3329 12733 3341 12736
rect 3375 12733 3387 12767
rect 5350 12764 5356 12776
rect 5311 12736 5356 12764
rect 3329 12727 3387 12733
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 5442 12724 5448 12776
rect 5500 12764 5506 12776
rect 5718 12764 5724 12776
rect 5500 12736 5545 12764
rect 5679 12736 5724 12764
rect 5500 12724 5506 12736
rect 5718 12724 5724 12736
rect 5776 12724 5782 12776
rect 7466 12764 7472 12776
rect 7427 12736 7472 12764
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 7650 12724 7656 12776
rect 7708 12764 7714 12776
rect 7745 12767 7803 12773
rect 7745 12764 7757 12767
rect 7708 12736 7757 12764
rect 7708 12724 7714 12736
rect 7745 12733 7757 12736
rect 7791 12733 7803 12767
rect 7745 12727 7803 12733
rect 7834 12724 7840 12776
rect 7892 12764 7898 12776
rect 12820 12773 12848 12804
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 14829 12835 14887 12841
rect 14829 12801 14841 12835
rect 14875 12832 14887 12835
rect 15120 12832 15148 12860
rect 15657 12835 15715 12841
rect 15657 12832 15669 12835
rect 14875 12804 15669 12832
rect 14875 12801 14887 12804
rect 14829 12795 14887 12801
rect 15657 12801 15669 12804
rect 15703 12801 15715 12835
rect 15657 12795 15715 12801
rect 10965 12767 11023 12773
rect 7892 12736 7937 12764
rect 7892 12724 7898 12736
rect 10965 12733 10977 12767
rect 11011 12764 11023 12767
rect 12713 12767 12771 12773
rect 12713 12764 12725 12767
rect 11011 12736 12725 12764
rect 11011 12733 11023 12736
rect 10965 12727 11023 12733
rect 12713 12733 12725 12736
rect 12759 12733 12771 12767
rect 12713 12727 12771 12733
rect 12805 12767 12863 12773
rect 12805 12733 12817 12767
rect 12851 12733 12863 12767
rect 12805 12727 12863 12733
rect 13081 12767 13139 12773
rect 13081 12733 13093 12767
rect 13127 12764 13139 12767
rect 13538 12764 13544 12776
rect 13127 12736 13544 12764
rect 13127 12733 13139 12736
rect 13081 12727 13139 12733
rect 9493 12699 9551 12705
rect 9493 12665 9505 12699
rect 9539 12696 9551 12699
rect 11514 12696 11520 12708
rect 9539 12668 11520 12696
rect 9539 12665 9551 12668
rect 9493 12659 9551 12665
rect 11514 12656 11520 12668
rect 11572 12656 11578 12708
rect 9401 12631 9459 12637
rect 9401 12597 9413 12631
rect 9447 12628 9459 12631
rect 10686 12628 10692 12640
rect 9447 12600 10692 12628
rect 9447 12597 9459 12600
rect 9401 12591 9459 12597
rect 10686 12588 10692 12600
rect 10744 12588 10750 12640
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12529 12631 12587 12637
rect 12529 12628 12541 12631
rect 12492 12600 12541 12628
rect 12492 12588 12498 12600
rect 12529 12597 12541 12600
rect 12575 12597 12587 12631
rect 12728 12628 12756 12727
rect 13538 12724 13544 12736
rect 13596 12724 13602 12776
rect 15010 12724 15016 12776
rect 15068 12764 15074 12776
rect 15105 12767 15163 12773
rect 15105 12764 15117 12767
rect 15068 12736 15117 12764
rect 15068 12724 15074 12736
rect 15105 12733 15117 12736
rect 15151 12733 15163 12767
rect 15746 12764 15752 12776
rect 15707 12736 15752 12764
rect 15105 12727 15163 12733
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 17126 12724 17132 12776
rect 17184 12764 17190 12776
rect 17497 12767 17555 12773
rect 17497 12764 17509 12767
rect 17184 12736 17509 12764
rect 17184 12724 17190 12736
rect 17497 12733 17509 12736
rect 17543 12733 17555 12767
rect 17497 12727 17555 12733
rect 17770 12724 17776 12776
rect 17828 12764 17834 12776
rect 17865 12767 17923 12773
rect 17865 12764 17877 12767
rect 17828 12736 17877 12764
rect 17828 12724 17834 12736
rect 17865 12733 17877 12736
rect 17911 12733 17923 12767
rect 17865 12727 17923 12733
rect 12897 12699 12955 12705
rect 12897 12665 12909 12699
rect 12943 12696 12955 12699
rect 13814 12696 13820 12708
rect 12943 12668 13820 12696
rect 12943 12665 12955 12668
rect 12897 12659 12955 12665
rect 13814 12656 13820 12668
rect 13872 12656 13878 12708
rect 17589 12699 17647 12705
rect 17589 12665 17601 12699
rect 17635 12665 17647 12699
rect 17589 12659 17647 12665
rect 13998 12628 14004 12640
rect 12728 12600 14004 12628
rect 12529 12591 12587 12597
rect 13998 12588 14004 12600
rect 14056 12588 14062 12640
rect 16850 12588 16856 12640
rect 16908 12628 16914 12640
rect 17313 12631 17371 12637
rect 17313 12628 17325 12631
rect 16908 12600 17325 12628
rect 16908 12588 16914 12600
rect 17313 12597 17325 12600
rect 17359 12597 17371 12631
rect 17604 12628 17632 12659
rect 17678 12656 17684 12708
rect 17736 12696 17742 12708
rect 17736 12668 17781 12696
rect 17736 12656 17742 12668
rect 18322 12628 18328 12640
rect 17604 12600 18328 12628
rect 17313 12591 17371 12597
rect 18322 12588 18328 12600
rect 18380 12588 18386 12640
rect 1104 12538 19044 12560
rect 1104 12486 6962 12538
rect 7014 12486 7026 12538
rect 7078 12486 7090 12538
rect 7142 12486 7154 12538
rect 7206 12486 12942 12538
rect 12994 12486 13006 12538
rect 13058 12486 13070 12538
rect 13122 12486 13134 12538
rect 13186 12486 19044 12538
rect 1104 12464 19044 12486
rect 8202 12384 8208 12436
rect 8260 12424 8266 12436
rect 11333 12427 11391 12433
rect 8260 12396 10640 12424
rect 8260 12384 8266 12396
rect 2225 12359 2283 12365
rect 2225 12325 2237 12359
rect 2271 12356 2283 12359
rect 3142 12356 3148 12368
rect 2271 12328 3004 12356
rect 3103 12328 3148 12356
rect 2271 12325 2283 12328
rect 2225 12319 2283 12325
rect 2976 12300 3004 12328
rect 3142 12316 3148 12328
rect 3200 12316 3206 12368
rect 4522 12356 4528 12368
rect 4483 12328 4528 12356
rect 4522 12316 4528 12328
rect 4580 12316 4586 12368
rect 7650 12316 7656 12368
rect 7708 12356 7714 12368
rect 7708 12328 9812 12356
rect 7708 12316 7714 12328
rect 1765 12291 1823 12297
rect 1765 12257 1777 12291
rect 1811 12288 1823 12291
rect 2130 12288 2136 12300
rect 1811 12260 2136 12288
rect 1811 12257 1823 12260
rect 1765 12251 1823 12257
rect 2130 12248 2136 12260
rect 2188 12248 2194 12300
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12288 2375 12291
rect 2958 12288 2964 12300
rect 2363 12260 2774 12288
rect 2919 12260 2964 12288
rect 2363 12257 2375 12260
rect 2317 12251 2375 12257
rect 2746 12220 2774 12260
rect 2958 12248 2964 12260
rect 3016 12248 3022 12300
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 6549 12291 6607 12297
rect 5592 12260 5658 12288
rect 5592 12248 5598 12260
rect 6549 12257 6561 12291
rect 6595 12288 6607 12291
rect 6595 12260 6776 12288
rect 6595 12257 6607 12260
rect 6549 12251 6607 12257
rect 3142 12220 3148 12232
rect 2746 12192 3148 12220
rect 3142 12180 3148 12192
rect 3200 12180 3206 12232
rect 4249 12223 4307 12229
rect 4249 12189 4261 12223
rect 4295 12220 4307 12223
rect 4295 12192 5580 12220
rect 4295 12189 4307 12192
rect 4249 12183 4307 12189
rect 5552 12152 5580 12192
rect 5718 12180 5724 12232
rect 5776 12220 5782 12232
rect 6270 12220 6276 12232
rect 5776 12192 6276 12220
rect 5776 12180 5782 12192
rect 6270 12180 6276 12192
rect 6328 12220 6334 12232
rect 6641 12223 6699 12229
rect 6641 12220 6653 12223
rect 6328 12192 6653 12220
rect 6328 12180 6334 12192
rect 6641 12189 6653 12192
rect 6687 12189 6699 12223
rect 6641 12183 6699 12189
rect 5902 12152 5908 12164
rect 5552 12124 5908 12152
rect 5902 12112 5908 12124
rect 5960 12112 5966 12164
rect 6748 12152 6776 12260
rect 6914 12248 6920 12300
rect 6972 12288 6978 12300
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 6972 12260 7481 12288
rect 6972 12248 6978 12260
rect 7469 12257 7481 12260
rect 7515 12288 7527 12291
rect 8018 12288 8024 12300
rect 7515 12260 8024 12288
rect 7515 12257 7527 12260
rect 7469 12251 7527 12257
rect 8018 12248 8024 12260
rect 8076 12288 8082 12300
rect 8202 12288 8208 12300
rect 8076 12260 8208 12288
rect 8076 12248 8082 12260
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 8481 12291 8539 12297
rect 8481 12257 8493 12291
rect 8527 12288 8539 12291
rect 8754 12288 8760 12300
rect 8527 12260 8760 12288
rect 8527 12257 8539 12260
rect 8481 12251 8539 12257
rect 8754 12248 8760 12260
rect 8812 12248 8818 12300
rect 9398 12248 9404 12300
rect 9456 12288 9462 12300
rect 9784 12297 9812 12328
rect 9677 12291 9735 12297
rect 9677 12288 9689 12291
rect 9456 12260 9689 12288
rect 9456 12248 9462 12260
rect 9677 12257 9689 12260
rect 9723 12257 9735 12291
rect 9677 12251 9735 12257
rect 9769 12291 9827 12297
rect 9769 12257 9781 12291
rect 9815 12257 9827 12291
rect 9769 12251 9827 12257
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12288 10103 12291
rect 10505 12291 10563 12297
rect 10505 12288 10517 12291
rect 10091 12260 10517 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 10505 12257 10517 12260
rect 10551 12257 10563 12291
rect 10612 12288 10640 12396
rect 11333 12393 11345 12427
rect 11379 12424 11391 12427
rect 11422 12424 11428 12436
rect 11379 12396 11428 12424
rect 11379 12393 11391 12396
rect 11333 12387 11391 12393
rect 11422 12384 11428 12396
rect 11480 12384 11486 12436
rect 13817 12427 13875 12433
rect 13817 12393 13829 12427
rect 13863 12424 13875 12427
rect 13906 12424 13912 12436
rect 13863 12396 13912 12424
rect 13863 12393 13875 12396
rect 13817 12387 13875 12393
rect 13906 12384 13912 12396
rect 13964 12384 13970 12436
rect 18322 12424 18328 12436
rect 18283 12396 18328 12424
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 12345 12359 12403 12365
rect 12345 12325 12357 12359
rect 12391 12356 12403 12359
rect 12434 12356 12440 12368
rect 12391 12328 12440 12356
rect 12391 12325 12403 12328
rect 12345 12319 12403 12325
rect 12434 12316 12440 12328
rect 12492 12316 12498 12368
rect 13354 12316 13360 12368
rect 13412 12316 13418 12368
rect 14918 12316 14924 12368
rect 14976 12356 14982 12368
rect 16850 12356 16856 12368
rect 14976 12328 16620 12356
rect 16811 12328 16856 12356
rect 14976 12316 14982 12328
rect 11146 12288 11152 12300
rect 10612 12260 11152 12288
rect 10505 12251 10563 12257
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 9953 12223 10011 12229
rect 9953 12220 9965 12223
rect 7616 12192 9965 12220
rect 7616 12180 7622 12192
rect 9953 12189 9965 12192
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 8478 12152 8484 12164
rect 6748 12124 8484 12152
rect 5258 12044 5264 12096
rect 5316 12084 5322 12096
rect 5997 12087 6055 12093
rect 5997 12084 6009 12087
rect 5316 12056 6009 12084
rect 5316 12044 5322 12056
rect 5997 12053 6009 12056
rect 6043 12084 6055 12087
rect 6748 12084 6776 12124
rect 8478 12112 8484 12124
rect 8536 12112 8542 12164
rect 9493 12155 9551 12161
rect 9493 12121 9505 12155
rect 9539 12152 9551 12155
rect 9582 12152 9588 12164
rect 9539 12124 9588 12152
rect 9539 12121 9551 12124
rect 9493 12115 9551 12121
rect 9582 12112 9588 12124
rect 9640 12112 9646 12164
rect 9674 12112 9680 12164
rect 9732 12152 9738 12164
rect 10060 12152 10088 12251
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 13998 12248 14004 12300
rect 14056 12288 14062 12300
rect 16592 12297 16620 12328
rect 16850 12316 16856 12328
rect 16908 12316 16914 12368
rect 15105 12291 15163 12297
rect 15105 12288 15117 12291
rect 14056 12260 15117 12288
rect 14056 12248 14062 12260
rect 15105 12257 15117 12260
rect 15151 12257 15163 12291
rect 15105 12251 15163 12257
rect 16577 12291 16635 12297
rect 16577 12257 16589 12291
rect 16623 12257 16635 12291
rect 16577 12251 16635 12257
rect 17954 12248 17960 12300
rect 18012 12248 18018 12300
rect 10410 12180 10416 12232
rect 10468 12220 10474 12232
rect 12069 12223 12127 12229
rect 12069 12220 12081 12223
rect 10468 12192 12081 12220
rect 10468 12180 10474 12192
rect 12069 12189 12081 12192
rect 12115 12220 12127 12223
rect 14182 12220 14188 12232
rect 12115 12192 14188 12220
rect 12115 12189 12127 12192
rect 12069 12183 12127 12189
rect 14182 12180 14188 12192
rect 14240 12180 14246 12232
rect 11054 12152 11060 12164
rect 9732 12124 11060 12152
rect 9732 12112 9738 12124
rect 11054 12112 11060 12124
rect 11112 12112 11118 12164
rect 7650 12084 7656 12096
rect 6043 12056 6776 12084
rect 7611 12056 7656 12084
rect 6043 12053 6055 12056
rect 5997 12047 6055 12053
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 8294 12044 8300 12096
rect 8352 12084 8358 12096
rect 8389 12087 8447 12093
rect 8389 12084 8401 12087
rect 8352 12056 8401 12084
rect 8352 12044 8358 12056
rect 8389 12053 8401 12056
rect 8435 12053 8447 12087
rect 8389 12047 8447 12053
rect 9398 12044 9404 12096
rect 9456 12084 9462 12096
rect 10597 12087 10655 12093
rect 10597 12084 10609 12087
rect 9456 12056 10609 12084
rect 9456 12044 9462 12056
rect 10597 12053 10609 12056
rect 10643 12084 10655 12087
rect 10778 12084 10784 12096
rect 10643 12056 10784 12084
rect 10643 12053 10655 12056
rect 10597 12047 10655 12053
rect 10778 12044 10784 12056
rect 10836 12044 10842 12096
rect 15194 12044 15200 12096
rect 15252 12084 15258 12096
rect 15289 12087 15347 12093
rect 15289 12084 15301 12087
rect 15252 12056 15301 12084
rect 15252 12044 15258 12056
rect 15289 12053 15301 12056
rect 15335 12053 15347 12087
rect 15289 12047 15347 12053
rect 1104 11994 19044 12016
rect 1104 11942 3972 11994
rect 4024 11942 4036 11994
rect 4088 11942 4100 11994
rect 4152 11942 4164 11994
rect 4216 11942 9952 11994
rect 10004 11942 10016 11994
rect 10068 11942 10080 11994
rect 10132 11942 10144 11994
rect 10196 11942 15932 11994
rect 15984 11942 15996 11994
rect 16048 11942 16060 11994
rect 16112 11942 16124 11994
rect 16176 11942 19044 11994
rect 1104 11920 19044 11942
rect 2130 11840 2136 11892
rect 2188 11880 2194 11892
rect 2225 11883 2283 11889
rect 2225 11880 2237 11883
rect 2188 11852 2237 11880
rect 2188 11840 2194 11852
rect 2225 11849 2237 11852
rect 2271 11849 2283 11883
rect 2225 11843 2283 11849
rect 1578 11744 1584 11756
rect 1539 11716 1584 11744
rect 1578 11704 1584 11716
rect 1636 11704 1642 11756
rect 1762 11744 1768 11756
rect 1723 11716 1768 11744
rect 1762 11704 1768 11716
rect 1820 11704 1826 11756
rect 2240 11744 2268 11843
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3053 11883 3111 11889
rect 3053 11880 3065 11883
rect 3016 11852 3065 11880
rect 3016 11840 3022 11852
rect 3053 11849 3065 11852
rect 3099 11849 3111 11883
rect 3053 11843 3111 11849
rect 4430 11840 4436 11892
rect 4488 11880 4494 11892
rect 4525 11883 4583 11889
rect 4525 11880 4537 11883
rect 4488 11852 4537 11880
rect 4488 11840 4494 11852
rect 4525 11849 4537 11852
rect 4571 11849 4583 11883
rect 5350 11880 5356 11892
rect 4525 11843 4583 11849
rect 4816 11852 5356 11880
rect 4816 11753 4844 11852
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 5534 11880 5540 11892
rect 5495 11852 5540 11880
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 6914 11840 6920 11892
rect 6972 11840 6978 11892
rect 7088 11883 7146 11889
rect 7088 11849 7100 11883
rect 7134 11880 7146 11883
rect 7190 11880 7196 11892
rect 7134 11852 7196 11880
rect 7134 11849 7146 11852
rect 7088 11843 7146 11849
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 7282 11840 7288 11892
rect 7340 11880 7346 11892
rect 7834 11880 7840 11892
rect 7340 11852 7840 11880
rect 7340 11840 7346 11852
rect 7834 11840 7840 11852
rect 7892 11880 7898 11892
rect 8573 11883 8631 11889
rect 8573 11880 8585 11883
rect 7892 11852 8585 11880
rect 7892 11840 7898 11852
rect 8573 11849 8585 11852
rect 8619 11849 8631 11883
rect 8573 11843 8631 11849
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 9861 11883 9919 11889
rect 9861 11880 9873 11883
rect 9824 11852 9873 11880
rect 9824 11840 9830 11852
rect 9861 11849 9873 11852
rect 9907 11849 9919 11883
rect 13354 11880 13360 11892
rect 13315 11852 13360 11880
rect 9861 11843 9919 11849
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 17954 11880 17960 11892
rect 17915 11852 17960 11880
rect 17954 11840 17960 11852
rect 18012 11840 18018 11892
rect 4982 11772 4988 11824
rect 5040 11812 5046 11824
rect 6932 11812 6960 11840
rect 5040 11784 5120 11812
rect 5040 11772 5046 11784
rect 2685 11747 2743 11753
rect 2685 11744 2697 11747
rect 2240 11716 2697 11744
rect 2685 11713 2697 11716
rect 2731 11713 2743 11747
rect 2685 11707 2743 11713
rect 4801 11747 4859 11753
rect 4801 11713 4813 11747
rect 4847 11713 4859 11747
rect 4801 11707 4859 11713
rect 3050 11676 3056 11688
rect 3011 11648 3056 11676
rect 3050 11636 3056 11648
rect 3108 11636 3114 11688
rect 4614 11636 4620 11688
rect 4672 11676 4678 11688
rect 4709 11679 4767 11685
rect 4709 11676 4721 11679
rect 4672 11648 4721 11676
rect 4672 11636 4678 11648
rect 4709 11645 4721 11648
rect 4755 11645 4767 11679
rect 4709 11639 4767 11645
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11645 4951 11679
rect 4893 11639 4951 11645
rect 4985 11679 5043 11685
rect 4985 11645 4997 11679
rect 5031 11676 5043 11679
rect 5092 11676 5120 11784
rect 5736 11784 6960 11812
rect 5736 11685 5764 11784
rect 8478 11772 8484 11824
rect 8536 11812 8542 11824
rect 9490 11812 9496 11824
rect 8536 11784 9496 11812
rect 8536 11772 8542 11784
rect 9490 11772 9496 11784
rect 9548 11772 9554 11824
rect 5902 11704 5908 11756
rect 5960 11744 5966 11756
rect 6546 11744 6552 11756
rect 5960 11716 6552 11744
rect 5960 11704 5966 11716
rect 6546 11704 6552 11716
rect 6604 11744 6610 11756
rect 6825 11747 6883 11753
rect 6825 11744 6837 11747
rect 6604 11716 6837 11744
rect 6604 11704 6610 11716
rect 6825 11713 6837 11716
rect 6871 11744 6883 11747
rect 7742 11744 7748 11756
rect 6871 11716 7748 11744
rect 6871 11713 6883 11716
rect 6825 11707 6883 11713
rect 7742 11704 7748 11716
rect 7800 11704 7806 11756
rect 7834 11704 7840 11756
rect 7892 11744 7898 11756
rect 9398 11744 9404 11756
rect 7892 11716 9260 11744
rect 9359 11716 9404 11744
rect 7892 11704 7898 11716
rect 5031 11648 5120 11676
rect 5721 11679 5779 11685
rect 5031 11645 5043 11648
rect 4985 11639 5043 11645
rect 5721 11645 5733 11679
rect 5767 11645 5779 11679
rect 9122 11676 9128 11688
rect 9083 11648 9128 11676
rect 5721 11639 5779 11645
rect 1857 11611 1915 11617
rect 1857 11577 1869 11611
rect 1903 11608 1915 11611
rect 4246 11608 4252 11620
rect 1903 11580 4252 11608
rect 1903 11577 1915 11580
rect 1857 11571 1915 11577
rect 4246 11568 4252 11580
rect 4304 11568 4310 11620
rect 4908 11608 4936 11639
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 9232 11676 9260 11716
rect 9398 11704 9404 11716
rect 9456 11704 9462 11756
rect 14458 11744 14464 11756
rect 14419 11716 14464 11744
rect 14458 11704 14464 11716
rect 14516 11704 14522 11756
rect 15746 11704 15752 11756
rect 15804 11744 15810 11756
rect 16209 11747 16267 11753
rect 16209 11744 16221 11747
rect 15804 11716 16221 11744
rect 15804 11704 15810 11716
rect 16209 11713 16221 11716
rect 16255 11713 16267 11747
rect 16209 11707 16267 11713
rect 9309 11679 9367 11685
rect 9309 11676 9321 11679
rect 9232 11648 9321 11676
rect 9309 11645 9321 11648
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11676 9643 11679
rect 10318 11676 10324 11688
rect 9631 11648 10324 11676
rect 9631 11645 9643 11648
rect 9585 11639 9643 11645
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 10594 11676 10600 11688
rect 10555 11648 10600 11676
rect 10594 11636 10600 11648
rect 10652 11636 10658 11688
rect 10778 11676 10784 11688
rect 10739 11648 10784 11676
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 11146 11636 11152 11688
rect 11204 11676 11210 11688
rect 13541 11679 13599 11685
rect 13541 11676 13553 11679
rect 11204 11648 13553 11676
rect 11204 11636 11210 11648
rect 13541 11645 13553 11648
rect 13587 11676 13599 11679
rect 13998 11676 14004 11688
rect 13587 11648 14004 11676
rect 13587 11645 13599 11648
rect 13541 11639 13599 11645
rect 13998 11636 14004 11648
rect 14056 11636 14062 11688
rect 14182 11676 14188 11688
rect 14143 11648 14188 11676
rect 14182 11636 14188 11648
rect 14240 11636 14246 11688
rect 17497 11679 17555 11685
rect 17497 11676 17509 11679
rect 16546 11648 17509 11676
rect 7374 11608 7380 11620
rect 4908 11580 7380 11608
rect 7374 11568 7380 11580
rect 7432 11568 7438 11620
rect 7650 11568 7656 11620
rect 7708 11568 7714 11620
rect 11330 11608 11336 11620
rect 8496 11580 11336 11608
rect 4890 11500 4896 11552
rect 4948 11540 4954 11552
rect 8496 11540 8524 11580
rect 11330 11568 11336 11580
rect 11388 11568 11394 11620
rect 4948 11512 8524 11540
rect 10781 11543 10839 11549
rect 4948 11500 4954 11512
rect 10781 11509 10793 11543
rect 10827 11540 10839 11543
rect 11146 11540 11152 11552
rect 10827 11512 11152 11540
rect 10827 11509 10839 11512
rect 10781 11503 10839 11509
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 14016 11540 14044 11636
rect 15194 11568 15200 11620
rect 15252 11568 15258 11620
rect 16546 11540 16574 11648
rect 17497 11645 17509 11648
rect 17543 11676 17555 11679
rect 18141 11679 18199 11685
rect 18141 11676 18153 11679
rect 17543 11648 18153 11676
rect 17543 11645 17555 11648
rect 17497 11639 17555 11645
rect 18141 11645 18153 11648
rect 18187 11676 18199 11679
rect 18506 11676 18512 11688
rect 18187 11648 18512 11676
rect 18187 11645 18199 11648
rect 18141 11639 18199 11645
rect 18506 11636 18512 11648
rect 18564 11636 18570 11688
rect 14016 11512 16574 11540
rect 17313 11543 17371 11549
rect 17313 11509 17325 11543
rect 17359 11540 17371 11543
rect 17402 11540 17408 11552
rect 17359 11512 17408 11540
rect 17359 11509 17371 11512
rect 17313 11503 17371 11509
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 1104 11450 19044 11472
rect 1104 11398 6962 11450
rect 7014 11398 7026 11450
rect 7078 11398 7090 11450
rect 7142 11398 7154 11450
rect 7206 11398 12942 11450
rect 12994 11398 13006 11450
rect 13058 11398 13070 11450
rect 13122 11398 13134 11450
rect 13186 11398 19044 11450
rect 1104 11376 19044 11398
rect 1486 11336 1492 11348
rect 1447 11308 1492 11336
rect 1486 11296 1492 11308
rect 1544 11296 1550 11348
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 3050 11336 3056 11348
rect 2915 11308 3056 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 3050 11296 3056 11308
rect 3108 11296 3114 11348
rect 4246 11336 4252 11348
rect 4207 11308 4252 11336
rect 4246 11296 4252 11308
rect 4304 11296 4310 11348
rect 5074 11296 5080 11348
rect 5132 11336 5138 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 5132 11308 5181 11336
rect 5132 11296 5138 11308
rect 5169 11305 5181 11308
rect 5215 11336 5227 11339
rect 5215 11308 6132 11336
rect 5215 11305 5227 11308
rect 5169 11299 5227 11305
rect 4522 11228 4528 11280
rect 4580 11228 4586 11280
rect 6104 11277 6132 11308
rect 7466 11296 7472 11348
rect 7524 11336 7530 11348
rect 7653 11339 7711 11345
rect 7653 11336 7665 11339
rect 7524 11308 7665 11336
rect 7524 11296 7530 11308
rect 7653 11305 7665 11308
rect 7699 11305 7711 11339
rect 7653 11299 7711 11305
rect 8573 11339 8631 11345
rect 8573 11305 8585 11339
rect 8619 11336 8631 11339
rect 10229 11339 10287 11345
rect 10229 11336 10241 11339
rect 8619 11308 10241 11336
rect 8619 11305 8631 11308
rect 8573 11299 8631 11305
rect 10229 11305 10241 11308
rect 10275 11336 10287 11339
rect 10594 11336 10600 11348
rect 10275 11308 10600 11336
rect 10275 11305 10287 11308
rect 10229 11299 10287 11305
rect 6089 11271 6147 11277
rect 6089 11237 6101 11271
rect 6135 11237 6147 11271
rect 6270 11268 6276 11280
rect 6231 11240 6276 11268
rect 6089 11231 6147 11237
rect 6270 11228 6276 11240
rect 6328 11228 6334 11280
rect 7668 11268 7696 11299
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 11330 11336 11336 11348
rect 11291 11308 11336 11336
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 11793 11339 11851 11345
rect 11793 11305 11805 11339
rect 11839 11336 11851 11339
rect 12618 11336 12624 11348
rect 11839 11308 12624 11336
rect 11839 11305 11851 11308
rect 11793 11299 11851 11305
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 17678 11296 17684 11348
rect 17736 11336 17742 11348
rect 17865 11339 17923 11345
rect 17865 11336 17877 11339
rect 17736 11308 17877 11336
rect 17736 11296 17742 11308
rect 17865 11305 17877 11308
rect 17911 11305 17923 11339
rect 17865 11299 17923 11305
rect 9122 11268 9128 11280
rect 7668 11240 9128 11268
rect 1581 11203 1639 11209
rect 1581 11169 1593 11203
rect 1627 11169 1639 11203
rect 1581 11163 1639 11169
rect 1596 11064 1624 11163
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 4540 11200 4568 11228
rect 4617 11203 4675 11209
rect 4617 11200 4629 11203
rect 2832 11172 2877 11200
rect 4540 11172 4629 11200
rect 2832 11160 2838 11172
rect 4617 11169 4629 11172
rect 4663 11169 4675 11203
rect 4617 11163 4675 11169
rect 4706 11160 4712 11212
rect 4764 11200 4770 11212
rect 5074 11200 5080 11212
rect 4764 11172 5080 11200
rect 4764 11160 4770 11172
rect 5074 11160 5080 11172
rect 5132 11200 5138 11212
rect 5261 11203 5319 11209
rect 5261 11200 5273 11203
rect 5132 11172 5273 11200
rect 5132 11160 5138 11172
rect 5261 11169 5273 11172
rect 5307 11169 5319 11203
rect 5261 11163 5319 11169
rect 5350 11160 5356 11212
rect 5408 11200 5414 11212
rect 6917 11203 6975 11209
rect 6917 11200 6929 11203
rect 5408 11172 6929 11200
rect 5408 11160 5414 11172
rect 6917 11169 6929 11172
rect 6963 11200 6975 11203
rect 7190 11200 7196 11212
rect 6963 11172 7196 11200
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7374 11160 7380 11212
rect 7432 11200 7438 11212
rect 7561 11203 7619 11209
rect 7561 11200 7573 11203
rect 7432 11172 7573 11200
rect 7432 11160 7438 11172
rect 7561 11169 7573 11172
rect 7607 11169 7619 11203
rect 8202 11200 8208 11212
rect 8163 11172 8208 11200
rect 7561 11163 7619 11169
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 8312 11209 8340 11240
rect 9122 11228 9128 11240
rect 9180 11228 9186 11280
rect 10137 11271 10195 11277
rect 10137 11237 10149 11271
rect 10183 11268 10195 11271
rect 11054 11268 11060 11280
rect 10183 11240 11060 11268
rect 10183 11237 10195 11240
rect 10137 11231 10195 11237
rect 11054 11228 11060 11240
rect 11112 11268 11118 11280
rect 12437 11271 12495 11277
rect 12437 11268 12449 11271
rect 11112 11240 12449 11268
rect 11112 11228 11118 11240
rect 12437 11237 12449 11240
rect 12483 11237 12495 11271
rect 16390 11268 16396 11280
rect 16351 11240 16396 11268
rect 12437 11231 12495 11237
rect 16390 11228 16396 11240
rect 16448 11228 16454 11280
rect 17402 11228 17408 11280
rect 17460 11228 17466 11280
rect 8297 11203 8355 11209
rect 8297 11169 8309 11203
rect 8343 11169 8355 11203
rect 11422 11200 11428 11212
rect 11383 11172 11428 11200
rect 8297 11163 8355 11169
rect 11422 11160 11428 11172
rect 11480 11160 11486 11212
rect 11514 11160 11520 11212
rect 11572 11160 11578 11212
rect 12250 11160 12256 11212
rect 12308 11200 12314 11212
rect 12621 11203 12679 11209
rect 12621 11200 12633 11203
rect 12308 11172 12633 11200
rect 12308 11160 12314 11172
rect 12621 11169 12633 11172
rect 12667 11169 12679 11203
rect 12621 11163 12679 11169
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11132 4583 11135
rect 4890 11132 4896 11144
rect 4571 11104 4896 11132
rect 4571 11101 4583 11104
rect 4525 11095 4583 11101
rect 4890 11092 4896 11104
rect 4948 11092 4954 11144
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11132 6515 11135
rect 8220 11132 8248 11160
rect 6503 11104 8248 11132
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 9306 11092 9312 11144
rect 9364 11132 9370 11144
rect 9674 11132 9680 11144
rect 9364 11104 9680 11132
rect 9364 11092 9370 11104
rect 9674 11092 9680 11104
rect 9732 11132 9738 11144
rect 9953 11135 10011 11141
rect 9953 11132 9965 11135
rect 9732 11104 9965 11132
rect 9732 11092 9738 11104
rect 9953 11101 9965 11104
rect 9999 11101 10011 11135
rect 9953 11095 10011 11101
rect 11241 11135 11299 11141
rect 11241 11101 11253 11135
rect 11287 11132 11299 11135
rect 11532 11132 11560 11160
rect 11698 11132 11704 11144
rect 11287 11104 11704 11132
rect 11287 11101 11299 11104
rect 11241 11095 11299 11101
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 14182 11092 14188 11144
rect 14240 11132 14246 11144
rect 14918 11132 14924 11144
rect 14240 11104 14924 11132
rect 14240 11092 14246 11104
rect 14918 11092 14924 11104
rect 14976 11132 14982 11144
rect 16117 11135 16175 11141
rect 16117 11132 16129 11135
rect 14976 11104 16129 11132
rect 14976 11092 14982 11104
rect 16117 11101 16129 11104
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 5718 11064 5724 11076
rect 1596 11036 5724 11064
rect 5718 11024 5724 11036
rect 5776 11024 5782 11076
rect 7009 11067 7067 11073
rect 7009 11033 7021 11067
rect 7055 11033 7067 11067
rect 7009 11027 7067 11033
rect 4617 10999 4675 11005
rect 4617 10965 4629 10999
rect 4663 10996 4675 10999
rect 5258 10996 5264 11008
rect 4663 10968 5264 10996
rect 4663 10965 4675 10968
rect 4617 10959 4675 10965
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 7024 10996 7052 11027
rect 7190 11024 7196 11076
rect 7248 11064 7254 11076
rect 7926 11064 7932 11076
rect 7248 11036 7932 11064
rect 7248 11024 7254 11036
rect 7926 11024 7932 11036
rect 7984 11024 7990 11076
rect 10597 11067 10655 11073
rect 10597 11033 10609 11067
rect 10643 11064 10655 11067
rect 10643 11036 11192 11064
rect 10643 11033 10655 11036
rect 10597 11027 10655 11033
rect 7282 10996 7288 11008
rect 7024 10968 7288 10996
rect 7282 10956 7288 10968
rect 7340 10996 7346 11008
rect 8110 10996 8116 11008
rect 7340 10968 8116 10996
rect 7340 10956 7346 10968
rect 8110 10956 8116 10968
rect 8168 10996 8174 11008
rect 8297 10999 8355 11005
rect 8297 10996 8309 10999
rect 8168 10968 8309 10996
rect 8168 10956 8174 10968
rect 8297 10965 8309 10968
rect 8343 10965 8355 10999
rect 11164 10996 11192 11036
rect 11514 10996 11520 11008
rect 11164 10968 11520 10996
rect 8297 10959 8355 10965
rect 11514 10956 11520 10968
rect 11572 10956 11578 11008
rect 12802 10996 12808 11008
rect 12763 10968 12808 10996
rect 12802 10956 12808 10968
rect 12860 10956 12866 11008
rect 1104 10906 19044 10928
rect 1104 10854 3972 10906
rect 4024 10854 4036 10906
rect 4088 10854 4100 10906
rect 4152 10854 4164 10906
rect 4216 10854 9952 10906
rect 10004 10854 10016 10906
rect 10068 10854 10080 10906
rect 10132 10854 10144 10906
rect 10196 10854 15932 10906
rect 15984 10854 15996 10906
rect 16048 10854 16060 10906
rect 16112 10854 16124 10906
rect 16176 10854 19044 10906
rect 1104 10832 19044 10854
rect 4614 10752 4620 10804
rect 4672 10792 4678 10804
rect 4893 10795 4951 10801
rect 4893 10792 4905 10795
rect 4672 10764 4905 10792
rect 4672 10752 4678 10764
rect 4893 10761 4905 10764
rect 4939 10792 4951 10795
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 4939 10764 5641 10792
rect 4939 10761 4951 10764
rect 4893 10755 4951 10761
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 5810 10792 5816 10804
rect 5771 10764 5816 10792
rect 5629 10755 5687 10761
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 9677 10795 9735 10801
rect 9677 10792 9689 10795
rect 7984 10764 9689 10792
rect 7984 10752 7990 10764
rect 9677 10761 9689 10764
rect 9723 10761 9735 10795
rect 11054 10792 11060 10804
rect 11015 10764 11060 10792
rect 9677 10755 9735 10761
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 11422 10752 11428 10804
rect 11480 10792 11486 10804
rect 12069 10795 12127 10801
rect 12069 10792 12081 10795
rect 11480 10764 12081 10792
rect 11480 10752 11486 10764
rect 12069 10761 12081 10764
rect 12115 10761 12127 10795
rect 12069 10755 12127 10761
rect 2777 10727 2835 10733
rect 2777 10693 2789 10727
rect 2823 10724 2835 10727
rect 3237 10727 3295 10733
rect 3237 10724 3249 10727
rect 2823 10696 3249 10724
rect 2823 10693 2835 10696
rect 2777 10687 2835 10693
rect 3237 10693 3249 10696
rect 3283 10693 3295 10727
rect 3237 10687 3295 10693
rect 4798 10684 4804 10736
rect 4856 10724 4862 10736
rect 18141 10727 18199 10733
rect 18141 10724 18153 10727
rect 4856 10696 18153 10724
rect 4856 10684 4862 10696
rect 18141 10693 18153 10696
rect 18187 10693 18199 10727
rect 18141 10687 18199 10693
rect 8389 10659 8447 10665
rect 8389 10656 8401 10659
rect 7392 10628 8401 10656
rect 7392 10600 7420 10628
rect 8389 10625 8401 10628
rect 8435 10625 8447 10659
rect 9398 10656 9404 10668
rect 8389 10619 8447 10625
rect 8588 10628 9404 10656
rect 2406 10588 2412 10600
rect 2367 10560 2412 10588
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 3050 10548 3056 10600
rect 3108 10588 3114 10600
rect 3421 10591 3479 10597
rect 3421 10588 3433 10591
rect 3108 10560 3433 10588
rect 3108 10548 3114 10560
rect 3421 10557 3433 10560
rect 3467 10557 3479 10591
rect 3421 10551 3479 10557
rect 4617 10591 4675 10597
rect 4617 10557 4629 10591
rect 4663 10588 4675 10591
rect 5074 10588 5080 10600
rect 4663 10560 5080 10588
rect 4663 10557 4675 10560
rect 4617 10551 4675 10557
rect 5074 10548 5080 10560
rect 5132 10548 5138 10600
rect 5629 10591 5687 10597
rect 5629 10557 5641 10591
rect 5675 10588 5687 10591
rect 5721 10591 5779 10597
rect 5721 10588 5733 10591
rect 5675 10560 5733 10588
rect 5675 10557 5687 10560
rect 5629 10551 5687 10557
rect 5721 10557 5733 10560
rect 5767 10588 5779 10591
rect 7009 10591 7067 10597
rect 5767 10560 6960 10588
rect 5767 10557 5779 10560
rect 5721 10551 5779 10557
rect 4801 10523 4859 10529
rect 4801 10489 4813 10523
rect 4847 10520 4859 10523
rect 5258 10520 5264 10532
rect 4847 10492 5264 10520
rect 4847 10489 4859 10492
rect 4801 10483 4859 10489
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 5350 10480 5356 10532
rect 5408 10520 5414 10532
rect 6825 10523 6883 10529
rect 6825 10520 6837 10523
rect 5408 10492 6837 10520
rect 5408 10480 5414 10492
rect 6825 10489 6837 10492
rect 6871 10489 6883 10523
rect 6932 10520 6960 10560
rect 7009 10557 7021 10591
rect 7055 10588 7067 10591
rect 7374 10588 7380 10600
rect 7055 10560 7380 10588
rect 7055 10557 7067 10560
rect 7009 10551 7067 10557
rect 7374 10548 7380 10560
rect 7432 10548 7438 10600
rect 8110 10548 8116 10600
rect 8168 10588 8174 10600
rect 8297 10591 8355 10597
rect 8297 10588 8309 10591
rect 8168 10560 8309 10588
rect 8168 10548 8174 10560
rect 8297 10557 8309 10560
rect 8343 10557 8355 10591
rect 8297 10551 8355 10557
rect 8478 10548 8484 10600
rect 8536 10588 8542 10600
rect 8588 10597 8616 10628
rect 9398 10616 9404 10628
rect 9456 10656 9462 10668
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 9456 10628 9781 10656
rect 9456 10616 9462 10628
rect 9769 10625 9781 10628
rect 9815 10625 9827 10659
rect 9769 10619 9827 10625
rect 11146 10616 11152 10668
rect 11204 10656 11210 10668
rect 11204 10628 11468 10656
rect 11204 10616 11210 10628
rect 8573 10591 8631 10597
rect 8573 10588 8585 10591
rect 8536 10560 8585 10588
rect 8536 10548 8542 10560
rect 8573 10557 8585 10560
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 9122 10548 9128 10600
rect 9180 10588 9186 10600
rect 9493 10591 9551 10597
rect 9493 10588 9505 10591
rect 9180 10560 9505 10588
rect 9180 10548 9186 10560
rect 9493 10557 9505 10560
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 9953 10591 10011 10597
rect 9953 10557 9965 10591
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 10229 10591 10287 10597
rect 10229 10557 10241 10591
rect 10275 10588 10287 10591
rect 11440 10588 11468 10628
rect 11514 10616 11520 10668
rect 11572 10656 11578 10668
rect 12437 10659 12495 10665
rect 12437 10656 12449 10659
rect 11572 10628 12449 10656
rect 11572 10616 11578 10628
rect 12437 10625 12449 10628
rect 12483 10625 12495 10659
rect 13538 10656 13544 10668
rect 13499 10628 13544 10656
rect 12437 10619 12495 10625
rect 13538 10616 13544 10628
rect 13596 10616 13602 10668
rect 12253 10591 12311 10597
rect 12253 10588 12265 10591
rect 10275 10560 11376 10588
rect 11440 10560 12265 10588
rect 10275 10557 10287 10560
rect 10229 10551 10287 10557
rect 9030 10520 9036 10532
rect 6932 10492 8892 10520
rect 8991 10492 9036 10520
rect 6825 10483 6883 10489
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 2832 10424 2877 10452
rect 2832 10412 2838 10424
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 7101 10455 7159 10461
rect 7101 10452 7113 10455
rect 4580 10424 7113 10452
rect 4580 10412 4586 10424
rect 7101 10421 7113 10424
rect 7147 10452 7159 10455
rect 8754 10452 8760 10464
rect 7147 10424 8760 10452
rect 7147 10421 7159 10424
rect 7101 10415 7159 10421
rect 8754 10412 8760 10424
rect 8812 10412 8818 10464
rect 8864 10452 8892 10492
rect 9030 10480 9036 10492
rect 9088 10480 9094 10532
rect 9490 10452 9496 10464
rect 8864 10424 9496 10452
rect 9490 10412 9496 10424
rect 9548 10452 9554 10464
rect 9876 10452 9904 10551
rect 9968 10520 9996 10551
rect 10318 10520 10324 10532
rect 9968 10492 10324 10520
rect 10318 10480 10324 10492
rect 10376 10480 10382 10532
rect 10686 10520 10692 10532
rect 10647 10492 10692 10520
rect 10686 10480 10692 10492
rect 10744 10480 10750 10532
rect 10873 10523 10931 10529
rect 10873 10489 10885 10523
rect 10919 10489 10931 10523
rect 11348 10520 11376 10560
rect 12253 10557 12265 10560
rect 12299 10557 12311 10591
rect 12253 10551 12311 10557
rect 12802 10548 12808 10600
rect 12860 10588 12866 10600
rect 13357 10591 13415 10597
rect 13357 10588 13369 10591
rect 12860 10560 13369 10588
rect 12860 10548 12866 10560
rect 13357 10557 13369 10560
rect 13403 10557 13415 10591
rect 13357 10551 13415 10557
rect 13449 10591 13507 10597
rect 13449 10557 13461 10591
rect 13495 10588 13507 10591
rect 14366 10588 14372 10600
rect 13495 10560 14372 10588
rect 13495 10557 13507 10560
rect 13449 10551 13507 10557
rect 14366 10548 14372 10560
rect 14424 10548 14430 10600
rect 14829 10591 14887 10597
rect 14829 10557 14841 10591
rect 14875 10588 14887 10591
rect 15102 10588 15108 10600
rect 14875 10560 15108 10588
rect 14875 10557 14887 10560
rect 14829 10551 14887 10557
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 15378 10588 15384 10600
rect 15339 10560 15384 10588
rect 15378 10548 15384 10560
rect 15436 10548 15442 10600
rect 18322 10588 18328 10600
rect 18283 10560 18328 10588
rect 18322 10548 18328 10560
rect 18380 10548 18386 10600
rect 15010 10520 15016 10532
rect 11348 10492 15016 10520
rect 10873 10483 10931 10489
rect 10888 10452 10916 10483
rect 15010 10480 15016 10492
rect 15068 10480 15074 10532
rect 15286 10520 15292 10532
rect 15247 10492 15292 10520
rect 15286 10480 15292 10492
rect 15344 10480 15350 10532
rect 9548 10424 10916 10452
rect 12989 10455 13047 10461
rect 9548 10412 9554 10424
rect 12989 10421 13001 10455
rect 13035 10452 13047 10455
rect 13262 10452 13268 10464
rect 13035 10424 13268 10452
rect 13035 10421 13047 10424
rect 12989 10415 13047 10421
rect 13262 10412 13268 10424
rect 13320 10412 13326 10464
rect 13446 10412 13452 10464
rect 13504 10452 13510 10464
rect 16482 10452 16488 10464
rect 13504 10424 16488 10452
rect 13504 10412 13510 10424
rect 16482 10412 16488 10424
rect 16540 10412 16546 10464
rect 1104 10362 19044 10384
rect 1104 10310 6962 10362
rect 7014 10310 7026 10362
rect 7078 10310 7090 10362
rect 7142 10310 7154 10362
rect 7206 10310 12942 10362
rect 12994 10310 13006 10362
rect 13058 10310 13070 10362
rect 13122 10310 13134 10362
rect 13186 10310 19044 10362
rect 1104 10288 19044 10310
rect 2406 10248 2412 10260
rect 2240 10220 2412 10248
rect 2240 10121 2268 10220
rect 2406 10208 2412 10220
rect 2464 10248 2470 10260
rect 10855 10251 10913 10257
rect 10855 10248 10867 10251
rect 2464 10220 10867 10248
rect 2464 10208 2470 10220
rect 10855 10217 10867 10220
rect 10901 10217 10913 10251
rect 10855 10211 10913 10217
rect 11333 10251 11391 10257
rect 11333 10217 11345 10251
rect 11379 10248 11391 10251
rect 17034 10248 17040 10260
rect 11379 10220 16574 10248
rect 16995 10220 17040 10248
rect 11379 10217 11391 10220
rect 11333 10211 11391 10217
rect 4798 10180 4804 10192
rect 4759 10152 4804 10180
rect 4798 10140 4804 10152
rect 4856 10140 4862 10192
rect 5258 10140 5264 10192
rect 5316 10180 5322 10192
rect 11146 10180 11152 10192
rect 5316 10152 6040 10180
rect 5316 10140 5322 10152
rect 2225 10115 2283 10121
rect 2225 10081 2237 10115
rect 2271 10081 2283 10115
rect 2225 10075 2283 10081
rect 2777 10115 2835 10121
rect 2777 10081 2789 10115
rect 2823 10112 2835 10115
rect 3050 10112 3056 10124
rect 2823 10084 3056 10112
rect 2823 10081 2835 10084
rect 2777 10075 2835 10081
rect 3050 10072 3056 10084
rect 3108 10072 3114 10124
rect 4706 10072 4712 10124
rect 4764 10112 4770 10124
rect 4893 10115 4951 10121
rect 4893 10112 4905 10115
rect 4764 10084 4905 10112
rect 4764 10072 4770 10084
rect 4893 10081 4905 10084
rect 4939 10081 4951 10115
rect 4893 10075 4951 10081
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 5905 10115 5963 10121
rect 5905 10112 5917 10115
rect 5592 10084 5917 10112
rect 5592 10072 5598 10084
rect 5905 10081 5917 10084
rect 5951 10081 5963 10115
rect 5905 10075 5963 10081
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 2774 9936 2780 9988
rect 2832 9976 2838 9988
rect 4816 9976 4844 10007
rect 5350 10004 5356 10056
rect 5408 10044 5414 10056
rect 5629 10047 5687 10053
rect 5629 10044 5641 10047
rect 5408 10016 5641 10044
rect 5408 10004 5414 10016
rect 5629 10013 5641 10016
rect 5675 10013 5687 10047
rect 5629 10007 5687 10013
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10044 5871 10047
rect 6012 10044 6040 10152
rect 6748 10152 7328 10180
rect 6270 10072 6276 10124
rect 6328 10112 6334 10124
rect 6748 10121 6776 10152
rect 6733 10115 6791 10121
rect 6733 10112 6745 10115
rect 6328 10084 6745 10112
rect 6328 10072 6334 10084
rect 6733 10081 6745 10084
rect 6779 10081 6791 10115
rect 6733 10075 6791 10081
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10112 6883 10115
rect 7190 10112 7196 10124
rect 6871 10084 7196 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 7190 10072 7196 10084
rect 7248 10072 7254 10124
rect 7300 10121 7328 10152
rect 8128 10152 9812 10180
rect 11107 10152 11152 10180
rect 7285 10115 7343 10121
rect 7285 10081 7297 10115
rect 7331 10081 7343 10115
rect 7285 10075 7343 10081
rect 8128 10056 8156 10152
rect 8294 10112 8300 10124
rect 8255 10084 8300 10112
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 8444 10084 8489 10112
rect 8444 10072 8450 10084
rect 9030 10072 9036 10124
rect 9088 10112 9094 10124
rect 9582 10112 9588 10124
rect 9088 10084 9588 10112
rect 9088 10072 9094 10084
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 9784 10121 9812 10152
rect 11146 10140 11152 10152
rect 11204 10140 11210 10192
rect 11716 10152 13400 10180
rect 9769 10115 9827 10121
rect 9769 10081 9781 10115
rect 9815 10081 9827 10115
rect 9769 10075 9827 10081
rect 11716 10056 11744 10152
rect 12250 10112 12256 10124
rect 12211 10084 12256 10112
rect 12250 10072 12256 10084
rect 12308 10072 12314 10124
rect 13265 10115 13323 10121
rect 13265 10112 13277 10115
rect 12452 10084 13277 10112
rect 5859 10016 6040 10044
rect 6549 10047 6607 10053
rect 5859 10013 5871 10016
rect 5813 10007 5871 10013
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 6638 10044 6644 10056
rect 6595 10016 6644 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 5445 9979 5503 9985
rect 5445 9976 5457 9979
rect 2832 9948 2877 9976
rect 4816 9948 5457 9976
rect 2832 9936 2838 9948
rect 5445 9945 5457 9948
rect 5491 9945 5503 9979
rect 5445 9939 5503 9945
rect 4341 9911 4399 9917
rect 4341 9877 4353 9911
rect 4387 9908 4399 9911
rect 4430 9908 4436 9920
rect 4387 9880 4436 9908
rect 4387 9877 4399 9880
rect 4341 9871 4399 9877
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 5074 9868 5080 9920
rect 5132 9908 5138 9920
rect 5736 9908 5764 10007
rect 6638 10004 6644 10016
rect 6696 10044 6702 10056
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 6696 10016 7389 10044
rect 6696 10004 6702 10016
rect 7377 10013 7389 10016
rect 7423 10013 7435 10047
rect 7558 10044 7564 10056
rect 7519 10016 7564 10044
rect 7377 10007 7435 10013
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 8110 10044 8116 10056
rect 8071 10016 8116 10044
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 9490 10044 9496 10056
rect 9451 10016 9496 10044
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10044 11483 10047
rect 11698 10044 11704 10056
rect 11471 10016 11704 10044
rect 11471 10013 11483 10016
rect 11425 10007 11483 10013
rect 11698 10004 11704 10016
rect 11756 10004 11762 10056
rect 12452 9985 12480 10084
rect 13265 10081 13277 10084
rect 13311 10081 13323 10115
rect 13372 10112 13400 10152
rect 13446 10140 13452 10192
rect 13504 10180 13510 10192
rect 13504 10152 13549 10180
rect 13504 10140 13510 10152
rect 15010 10140 15016 10192
rect 15068 10180 15074 10192
rect 15473 10183 15531 10189
rect 15473 10180 15485 10183
rect 15068 10152 15485 10180
rect 15068 10140 15074 10152
rect 15473 10149 15485 10152
rect 15519 10149 15531 10183
rect 16546 10180 16574 10220
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 18138 10180 18144 10192
rect 16546 10152 18144 10180
rect 15473 10143 15531 10149
rect 18138 10140 18144 10152
rect 18196 10140 18202 10192
rect 13538 10112 13544 10124
rect 13372 10084 13544 10112
rect 13265 10075 13323 10081
rect 13538 10072 13544 10084
rect 13596 10112 13602 10124
rect 15565 10115 15623 10121
rect 13596 10084 15332 10112
rect 13596 10072 13602 10084
rect 12526 10004 12532 10056
rect 12584 10044 12590 10056
rect 12971 10047 13029 10053
rect 12971 10044 12983 10047
rect 12584 10016 12983 10044
rect 12584 10004 12590 10016
rect 12971 10013 12983 10016
rect 13017 10013 13029 10047
rect 15304 10044 15332 10084
rect 15565 10081 15577 10115
rect 15611 10112 15623 10115
rect 16942 10112 16948 10124
rect 15611 10084 16948 10112
rect 15611 10081 15623 10084
rect 15565 10075 15623 10081
rect 16942 10072 16948 10084
rect 17000 10072 17006 10124
rect 17129 10115 17187 10121
rect 17129 10081 17141 10115
rect 17175 10081 17187 10115
rect 17129 10075 17187 10081
rect 15657 10047 15715 10053
rect 15657 10044 15669 10047
rect 15304 10016 15669 10044
rect 12971 10007 13029 10013
rect 15657 10013 15669 10016
rect 15703 10044 15715 10047
rect 16853 10047 16911 10053
rect 16853 10044 16865 10047
rect 15703 10016 16865 10044
rect 15703 10013 15715 10016
rect 15657 10007 15715 10013
rect 16853 10013 16865 10016
rect 16899 10013 16911 10047
rect 16853 10007 16911 10013
rect 9953 9979 10011 9985
rect 9953 9945 9965 9979
rect 9999 9976 10011 9979
rect 12437 9979 12495 9985
rect 9999 9948 11192 9976
rect 9999 9945 10011 9948
rect 9953 9939 10011 9945
rect 5132 9880 5764 9908
rect 6641 9911 6699 9917
rect 5132 9868 5138 9880
rect 6641 9877 6653 9911
rect 6687 9908 6699 9911
rect 6822 9908 6828 9920
rect 6687 9880 6828 9908
rect 6687 9877 6699 9880
rect 6641 9871 6699 9877
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 7466 9868 7472 9920
rect 7524 9908 7530 9920
rect 11164 9908 11192 9948
rect 12437 9945 12449 9979
rect 12483 9945 12495 9979
rect 15102 9976 15108 9988
rect 12437 9939 12495 9945
rect 12544 9948 14964 9976
rect 15063 9948 15108 9976
rect 12544 9908 12572 9948
rect 7524 9880 7569 9908
rect 11164 9880 12572 9908
rect 14936 9908 14964 9948
rect 15102 9936 15108 9948
rect 15160 9936 15166 9988
rect 17144 9976 17172 10075
rect 16546 9948 17172 9976
rect 16546 9908 16574 9948
rect 17494 9908 17500 9920
rect 14936 9880 16574 9908
rect 17455 9880 17500 9908
rect 7524 9868 7530 9880
rect 17494 9868 17500 9880
rect 17552 9868 17558 9920
rect 1104 9818 19044 9840
rect 1104 9766 3972 9818
rect 4024 9766 4036 9818
rect 4088 9766 4100 9818
rect 4152 9766 4164 9818
rect 4216 9766 9952 9818
rect 10004 9766 10016 9818
rect 10068 9766 10080 9818
rect 10132 9766 10144 9818
rect 10196 9766 15932 9818
rect 15984 9766 15996 9818
rect 16048 9766 16060 9818
rect 16112 9766 16124 9818
rect 16176 9766 19044 9818
rect 1104 9744 19044 9766
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 7653 9707 7711 9713
rect 7653 9704 7665 9707
rect 7616 9676 7665 9704
rect 7616 9664 7622 9676
rect 7653 9673 7665 9676
rect 7699 9673 7711 9707
rect 7653 9667 7711 9673
rect 4982 9596 4988 9648
rect 5040 9636 5046 9648
rect 5445 9639 5503 9645
rect 5445 9636 5457 9639
rect 5040 9608 5457 9636
rect 5040 9596 5046 9608
rect 5445 9605 5457 9608
rect 5491 9636 5503 9639
rect 5534 9636 5540 9648
rect 5491 9608 5540 9636
rect 5491 9605 5503 9608
rect 5445 9599 5503 9605
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 7282 9596 7288 9648
rect 7340 9636 7346 9648
rect 15381 9639 15439 9645
rect 7340 9608 7420 9636
rect 7340 9596 7346 9608
rect 1578 9528 1584 9580
rect 1636 9568 1642 9580
rect 7392 9577 7420 9608
rect 15381 9605 15393 9639
rect 15427 9636 15439 9639
rect 15841 9639 15899 9645
rect 15841 9636 15853 9639
rect 15427 9608 15853 9636
rect 15427 9605 15439 9608
rect 15381 9599 15439 9605
rect 15841 9605 15853 9608
rect 15887 9605 15899 9639
rect 18138 9636 18144 9648
rect 18099 9608 18144 9636
rect 15841 9599 15899 9605
rect 18138 9596 18144 9608
rect 18196 9596 18202 9648
rect 1673 9571 1731 9577
rect 1673 9568 1685 9571
rect 1636 9540 1685 9568
rect 1636 9528 1642 9540
rect 1673 9537 1685 9540
rect 1719 9537 1731 9571
rect 1673 9531 1731 9537
rect 4617 9571 4675 9577
rect 4617 9537 4629 9571
rect 4663 9568 4675 9571
rect 7377 9571 7435 9577
rect 4663 9540 7328 9568
rect 4663 9537 4675 9540
rect 4617 9531 4675 9537
rect 2866 9500 2872 9512
rect 2827 9472 2872 9500
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 3326 9460 3332 9512
rect 3384 9500 3390 9512
rect 4709 9503 4767 9509
rect 4709 9500 4721 9503
rect 3384 9472 4721 9500
rect 3384 9460 3390 9472
rect 4709 9469 4721 9472
rect 4755 9469 4767 9503
rect 4709 9463 4767 9469
rect 4801 9503 4859 9509
rect 4801 9469 4813 9503
rect 4847 9469 4859 9503
rect 4801 9463 4859 9469
rect 1670 9392 1676 9444
rect 1728 9432 1734 9444
rect 1765 9435 1823 9441
rect 1765 9432 1777 9435
rect 1728 9404 1777 9432
rect 1728 9392 1734 9404
rect 1765 9401 1777 9404
rect 1811 9401 1823 9435
rect 1765 9395 1823 9401
rect 2314 9392 2320 9444
rect 2372 9432 2378 9444
rect 2685 9435 2743 9441
rect 2685 9432 2697 9435
rect 2372 9404 2697 9432
rect 2372 9392 2378 9404
rect 2685 9401 2697 9404
rect 2731 9401 2743 9435
rect 2685 9395 2743 9401
rect 1854 9364 1860 9376
rect 1815 9336 1860 9364
rect 1854 9324 1860 9336
rect 1912 9324 1918 9376
rect 1946 9324 1952 9376
rect 2004 9364 2010 9376
rect 2225 9367 2283 9373
rect 2225 9364 2237 9367
rect 2004 9336 2237 9364
rect 2004 9324 2010 9336
rect 2225 9333 2237 9336
rect 2271 9333 2283 9367
rect 2225 9327 2283 9333
rect 4338 9324 4344 9376
rect 4396 9364 4402 9376
rect 4433 9367 4491 9373
rect 4433 9364 4445 9367
rect 4396 9336 4445 9364
rect 4396 9324 4402 9336
rect 4433 9333 4445 9336
rect 4479 9333 4491 9367
rect 4724 9364 4752 9463
rect 4816 9432 4844 9463
rect 4890 9460 4896 9512
rect 4948 9500 4954 9512
rect 5828 9509 5856 9540
rect 7300 9512 7328 9540
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 13262 9568 13268 9580
rect 8260 9540 9444 9568
rect 13223 9540 13268 9568
rect 8260 9528 8266 9540
rect 5629 9503 5687 9509
rect 5629 9500 5641 9503
rect 4948 9472 5641 9500
rect 4948 9460 4954 9472
rect 5629 9469 5641 9472
rect 5675 9469 5687 9503
rect 5629 9463 5687 9469
rect 5813 9503 5871 9509
rect 5813 9469 5825 9503
rect 5859 9469 5871 9503
rect 5813 9463 5871 9469
rect 5350 9432 5356 9444
rect 4816 9404 5356 9432
rect 5350 9392 5356 9404
rect 5408 9392 5414 9444
rect 5644 9432 5672 9463
rect 6638 9460 6644 9512
rect 6696 9500 6702 9512
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 6696 9472 7205 9500
rect 6696 9460 6702 9472
rect 7193 9469 7205 9472
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 7282 9460 7288 9512
rect 7340 9500 7346 9512
rect 7469 9503 7527 9509
rect 7340 9472 7433 9500
rect 7340 9460 7346 9472
rect 7469 9469 7481 9503
rect 7515 9500 7527 9503
rect 8386 9500 8392 9512
rect 7515 9472 8392 9500
rect 7515 9469 7527 9472
rect 7469 9463 7527 9469
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 8662 9500 8668 9512
rect 8575 9472 8668 9500
rect 8588 9432 8616 9472
rect 8662 9460 8668 9472
rect 8720 9460 8726 9512
rect 8849 9503 8907 9509
rect 8849 9469 8861 9503
rect 8895 9469 8907 9503
rect 8849 9463 8907 9469
rect 5644 9404 8616 9432
rect 5258 9364 5264 9376
rect 4724 9336 5264 9364
rect 4433 9327 4491 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 8478 9364 8484 9376
rect 8439 9336 8484 9364
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 8864 9364 8892 9463
rect 8938 9460 8944 9512
rect 8996 9500 9002 9512
rect 9416 9509 9444 9540
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 15013 9571 15071 9577
rect 15013 9537 15025 9571
rect 15059 9568 15071 9571
rect 15102 9568 15108 9580
rect 15059 9540 15108 9568
rect 15059 9537 15071 9540
rect 15013 9531 15071 9537
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 9401 9503 9459 9509
rect 8996 9472 9041 9500
rect 8996 9460 9002 9472
rect 9401 9469 9413 9503
rect 9447 9469 9459 9503
rect 9401 9463 9459 9469
rect 12802 9460 12808 9512
rect 12860 9500 12866 9512
rect 12897 9503 12955 9509
rect 12897 9500 12909 9503
rect 12860 9472 12909 9500
rect 12860 9460 12866 9472
rect 12897 9469 12909 9472
rect 12943 9469 12955 9503
rect 12897 9463 12955 9469
rect 15378 9460 15384 9512
rect 15436 9500 15442 9512
rect 16025 9503 16083 9509
rect 16025 9500 16037 9503
rect 15436 9472 16037 9500
rect 15436 9460 15442 9472
rect 16025 9469 16037 9472
rect 16071 9469 16083 9503
rect 18322 9500 18328 9512
rect 18283 9472 18328 9500
rect 16025 9463 16083 9469
rect 18322 9460 18328 9472
rect 18380 9460 18386 9512
rect 8956 9432 8984 9460
rect 9674 9432 9680 9444
rect 8956 9404 9680 9432
rect 9674 9392 9680 9404
rect 9732 9432 9738 9444
rect 10686 9432 10692 9444
rect 9732 9404 10692 9432
rect 9732 9392 9738 9404
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 9490 9364 9496 9376
rect 8864 9336 9496 9364
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 12710 9324 12716 9376
rect 12768 9364 12774 9376
rect 12897 9367 12955 9373
rect 12897 9364 12909 9367
rect 12768 9336 12909 9364
rect 12768 9324 12774 9336
rect 12897 9333 12909 9336
rect 12943 9333 12955 9367
rect 12897 9327 12955 9333
rect 15286 9324 15292 9376
rect 15344 9364 15350 9376
rect 15381 9367 15439 9373
rect 15381 9364 15393 9367
rect 15344 9336 15393 9364
rect 15344 9324 15350 9336
rect 15381 9333 15393 9336
rect 15427 9333 15439 9367
rect 15381 9327 15439 9333
rect 1104 9274 19044 9296
rect 1104 9222 6962 9274
rect 7014 9222 7026 9274
rect 7078 9222 7090 9274
rect 7142 9222 7154 9274
rect 7206 9222 12942 9274
rect 12994 9222 13006 9274
rect 13058 9222 13070 9274
rect 13122 9222 13134 9274
rect 13186 9222 19044 9274
rect 1104 9200 19044 9222
rect 1854 9120 1860 9172
rect 1912 9160 1918 9172
rect 2869 9163 2927 9169
rect 2869 9160 2881 9163
rect 1912 9132 2881 9160
rect 1912 9120 1918 9132
rect 2869 9129 2881 9132
rect 2915 9129 2927 9163
rect 2869 9123 2927 9129
rect 9582 9120 9588 9172
rect 9640 9160 9646 9172
rect 9698 9163 9756 9169
rect 9698 9160 9710 9163
rect 9640 9132 9710 9160
rect 9640 9120 9646 9132
rect 9698 9129 9710 9132
rect 9744 9129 9756 9163
rect 11238 9160 11244 9172
rect 11199 9132 11244 9160
rect 9698 9123 9756 9129
rect 11238 9120 11244 9132
rect 11296 9120 11302 9172
rect 15286 9120 15292 9172
rect 15344 9160 15350 9172
rect 15565 9163 15623 9169
rect 15565 9160 15577 9163
rect 15344 9132 15577 9160
rect 15344 9120 15350 9132
rect 15565 9129 15577 9132
rect 15611 9129 15623 9163
rect 15565 9123 15623 9129
rect 17589 9163 17647 9169
rect 17589 9129 17601 9163
rect 17635 9160 17647 9163
rect 17678 9160 17684 9172
rect 17635 9132 17684 9160
rect 17635 9129 17647 9132
rect 17589 9123 17647 9129
rect 17678 9120 17684 9132
rect 17736 9120 17742 9172
rect 5810 9052 5816 9104
rect 5868 9092 5874 9104
rect 5868 9064 6592 9092
rect 5868 9052 5874 9064
rect 1581 9027 1639 9033
rect 1581 8993 1593 9027
rect 1627 9024 1639 9027
rect 2498 9024 2504 9036
rect 1627 8996 2504 9024
rect 1627 8993 1639 8996
rect 1581 8987 1639 8993
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 3053 9027 3111 9033
rect 3053 8993 3065 9027
rect 3099 9024 3111 9027
rect 4890 9024 4896 9036
rect 3099 8996 4896 9024
rect 3099 8993 3111 8996
rect 3053 8987 3111 8993
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 5166 9033 5172 9036
rect 5158 9027 5172 9033
rect 5158 8993 5170 9027
rect 5224 9024 5230 9036
rect 5224 8996 5258 9024
rect 5158 8987 5172 8993
rect 5166 8984 5172 8987
rect 5224 8984 5230 8996
rect 5534 8984 5540 9036
rect 5592 9024 5598 9036
rect 6564 9033 6592 9064
rect 8662 9052 8668 9104
rect 8720 9092 8726 9104
rect 9306 9092 9312 9104
rect 8720 9064 9312 9092
rect 8720 9052 8726 9064
rect 9306 9052 9312 9064
rect 9364 9092 9370 9104
rect 9493 9095 9551 9101
rect 9493 9092 9505 9095
rect 9364 9064 9505 9092
rect 9364 9052 9370 9064
rect 9493 9061 9505 9064
rect 9539 9061 9551 9095
rect 9493 9055 9551 9061
rect 12621 9095 12679 9101
rect 12621 9061 12633 9095
rect 12667 9092 12679 9095
rect 12710 9092 12716 9104
rect 12667 9064 12716 9092
rect 12667 9061 12679 9064
rect 12621 9055 12679 9061
rect 12710 9052 12716 9064
rect 12768 9092 12774 9104
rect 14829 9095 14887 9101
rect 14829 9092 14841 9095
rect 12768 9064 14841 9092
rect 12768 9052 12774 9064
rect 14829 9061 14841 9064
rect 14875 9061 14887 9095
rect 14829 9055 14887 9061
rect 15013 9095 15071 9101
rect 15013 9061 15025 9095
rect 15059 9092 15071 9095
rect 15378 9092 15384 9104
rect 15059 9064 15384 9092
rect 15059 9061 15071 9064
rect 15013 9055 15071 9061
rect 15378 9052 15384 9064
rect 15436 9052 15442 9104
rect 5905 9027 5963 9033
rect 5905 9024 5917 9027
rect 5592 8996 5917 9024
rect 5592 8984 5598 8996
rect 5905 8993 5917 8996
rect 5951 8993 5963 9027
rect 5905 8987 5963 8993
rect 6549 9027 6607 9033
rect 6549 8993 6561 9027
rect 6595 8993 6607 9027
rect 6549 8987 6607 8993
rect 7285 9027 7343 9033
rect 7285 8993 7297 9027
rect 7331 9024 7343 9027
rect 7558 9024 7564 9036
rect 7331 8996 7564 9024
rect 7331 8993 7343 8996
rect 7285 8987 7343 8993
rect 3326 8956 3332 8968
rect 3287 8928 3332 8956
rect 3326 8916 3332 8928
rect 3384 8916 3390 8968
rect 4982 8916 4988 8968
rect 5040 8956 5046 8968
rect 5077 8959 5135 8965
rect 5077 8956 5089 8959
rect 5040 8928 5089 8956
rect 5040 8916 5046 8928
rect 5077 8925 5089 8928
rect 5123 8925 5135 8959
rect 5258 8956 5264 8968
rect 5219 8928 5264 8956
rect 5077 8919 5135 8925
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 5353 8959 5411 8965
rect 5353 8925 5365 8959
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8956 6055 8959
rect 6638 8956 6644 8968
rect 6043 8928 6644 8956
rect 6043 8925 6055 8928
rect 5997 8919 6055 8925
rect 1394 8888 1400 8900
rect 1355 8860 1400 8888
rect 1394 8848 1400 8860
rect 1452 8848 1458 8900
rect 3237 8823 3295 8829
rect 3237 8789 3249 8823
rect 3283 8820 3295 8823
rect 4522 8820 4528 8832
rect 3283 8792 4528 8820
rect 3283 8789 3295 8792
rect 3237 8783 3295 8789
rect 4522 8780 4528 8792
rect 4580 8780 4586 8832
rect 4614 8780 4620 8832
rect 4672 8820 4678 8832
rect 4893 8823 4951 8829
rect 4893 8820 4905 8823
rect 4672 8792 4905 8820
rect 4672 8780 4678 8792
rect 4893 8789 4905 8792
rect 4939 8789 4951 8823
rect 5368 8820 5396 8919
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 6825 8959 6883 8965
rect 6825 8925 6837 8959
rect 6871 8956 6883 8959
rect 7300 8956 7328 8987
rect 7558 8984 7564 8996
rect 7616 8984 7622 9036
rect 8202 8984 8208 9036
rect 8260 9024 8266 9036
rect 8297 9027 8355 9033
rect 8297 9024 8309 9027
rect 8260 8996 8309 9024
rect 8260 8984 8266 8996
rect 8297 8993 8309 8996
rect 8343 8993 8355 9027
rect 11333 9027 11391 9033
rect 11333 9024 11345 9027
rect 8297 8987 8355 8993
rect 8404 8996 11345 9024
rect 6871 8928 7328 8956
rect 7377 8959 7435 8965
rect 6871 8925 6883 8928
rect 6825 8919 6883 8925
rect 7377 8925 7389 8959
rect 7423 8956 7435 8959
rect 8404 8956 8432 8996
rect 11333 8993 11345 8996
rect 11379 8993 11391 9027
rect 11333 8987 11391 8993
rect 11790 8984 11796 9036
rect 11848 9024 11854 9036
rect 12529 9027 12587 9033
rect 12529 9024 12541 9027
rect 11848 8996 12541 9024
rect 11848 8984 11854 8996
rect 12529 8993 12541 8996
rect 12575 8993 12587 9027
rect 12529 8987 12587 8993
rect 13081 9027 13139 9033
rect 13081 8993 13093 9027
rect 13127 9024 13139 9027
rect 13262 9024 13268 9036
rect 13127 8996 13268 9024
rect 13127 8993 13139 8996
rect 13081 8987 13139 8993
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 16482 9024 16488 9036
rect 16443 8996 16488 9024
rect 16482 8984 16488 8996
rect 16540 8984 16546 9036
rect 17221 9027 17279 9033
rect 17221 8993 17233 9027
rect 17267 9024 17279 9027
rect 17494 9024 17500 9036
rect 17267 8996 17500 9024
rect 17267 8993 17279 8996
rect 17221 8987 17279 8993
rect 17494 8984 17500 8996
rect 17552 8984 17558 9036
rect 17862 8984 17868 9036
rect 17920 9024 17926 9036
rect 18233 9027 18291 9033
rect 18233 9024 18245 9027
rect 17920 8996 18245 9024
rect 17920 8984 17926 8996
rect 18233 8993 18245 8996
rect 18279 8993 18291 9027
rect 18233 8987 18291 8993
rect 7423 8928 8432 8956
rect 8573 8959 8631 8965
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 9490 8956 9496 8968
rect 8619 8928 9496 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 6546 8848 6552 8900
rect 6604 8888 6610 8900
rect 6733 8891 6791 8897
rect 6733 8888 6745 8891
rect 6604 8860 6745 8888
rect 6604 8848 6610 8860
rect 6733 8857 6745 8860
rect 6779 8857 6791 8891
rect 6733 8851 6791 8857
rect 7392 8820 7420 8919
rect 9490 8916 9496 8928
rect 9548 8916 9554 8968
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8956 11207 8959
rect 11698 8956 11704 8968
rect 11195 8928 11704 8956
rect 11195 8925 11207 8928
rect 11149 8919 11207 8925
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 8481 8891 8539 8897
rect 8481 8857 8493 8891
rect 8527 8888 8539 8891
rect 9582 8888 9588 8900
rect 8527 8860 9588 8888
rect 8527 8857 8539 8860
rect 8481 8851 8539 8857
rect 9582 8848 9588 8860
rect 9640 8848 9646 8900
rect 17589 8891 17647 8897
rect 17589 8857 17601 8891
rect 17635 8888 17647 8891
rect 18049 8891 18107 8897
rect 18049 8888 18061 8891
rect 17635 8860 18061 8888
rect 17635 8857 17647 8860
rect 17589 8851 17647 8857
rect 18049 8857 18061 8860
rect 18095 8857 18107 8891
rect 18049 8851 18107 8857
rect 5368 8792 7420 8820
rect 4893 8783 4951 8789
rect 8018 8780 8024 8832
rect 8076 8820 8082 8832
rect 8113 8823 8171 8829
rect 8113 8820 8125 8823
rect 8076 8792 8125 8820
rect 8076 8780 8082 8792
rect 8113 8789 8125 8792
rect 8159 8789 8171 8823
rect 9674 8820 9680 8832
rect 9635 8792 9680 8820
rect 8113 8783 8171 8789
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 9861 8823 9919 8829
rect 9861 8789 9873 8823
rect 9907 8820 9919 8823
rect 10318 8820 10324 8832
rect 9907 8792 10324 8820
rect 9907 8789 9919 8792
rect 9861 8783 9919 8789
rect 10318 8780 10324 8792
rect 10376 8820 10382 8832
rect 10686 8820 10692 8832
rect 10376 8792 10692 8820
rect 10376 8780 10382 8792
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 11701 8823 11759 8829
rect 11701 8789 11713 8823
rect 11747 8820 11759 8823
rect 14458 8820 14464 8832
rect 11747 8792 14464 8820
rect 11747 8789 11759 8792
rect 11701 8783 11759 8789
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 15654 8820 15660 8832
rect 15615 8792 15660 8820
rect 15654 8780 15660 8792
rect 15712 8780 15718 8832
rect 16574 8780 16580 8832
rect 16632 8820 16638 8832
rect 16632 8792 16677 8820
rect 16632 8780 16638 8792
rect 1104 8730 19044 8752
rect 1104 8678 3972 8730
rect 4024 8678 4036 8730
rect 4088 8678 4100 8730
rect 4152 8678 4164 8730
rect 4216 8678 9952 8730
rect 10004 8678 10016 8730
rect 10068 8678 10080 8730
rect 10132 8678 10144 8730
rect 10196 8678 15932 8730
rect 15984 8678 15996 8730
rect 16048 8678 16060 8730
rect 16112 8678 16124 8730
rect 16176 8678 19044 8730
rect 1104 8656 19044 8678
rect 2225 8619 2283 8625
rect 2225 8585 2237 8619
rect 2271 8616 2283 8619
rect 2590 8616 2596 8628
rect 2271 8588 2596 8616
rect 2271 8585 2283 8588
rect 2225 8579 2283 8585
rect 2590 8576 2596 8588
rect 2648 8616 2654 8628
rect 2685 8619 2743 8625
rect 2685 8616 2697 8619
rect 2648 8588 2697 8616
rect 2648 8576 2654 8588
rect 2685 8585 2697 8588
rect 2731 8585 2743 8619
rect 2685 8579 2743 8585
rect 5169 8619 5227 8625
rect 5169 8585 5181 8619
rect 5215 8616 5227 8619
rect 5442 8616 5448 8628
rect 5215 8588 5448 8616
rect 5215 8585 5227 8588
rect 5169 8579 5227 8585
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 9401 8619 9459 8625
rect 9401 8585 9413 8619
rect 9447 8616 9459 8619
rect 9582 8616 9588 8628
rect 9447 8588 9588 8616
rect 9447 8585 9459 8588
rect 9401 8579 9459 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8616 11207 8619
rect 12069 8619 12127 8625
rect 12069 8616 12081 8619
rect 11195 8588 12081 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 12069 8585 12081 8588
rect 12115 8616 12127 8619
rect 12115 8588 12572 8616
rect 12115 8585 12127 8588
rect 12069 8579 12127 8585
rect 4433 8551 4491 8557
rect 4433 8517 4445 8551
rect 4479 8548 4491 8551
rect 9769 8551 9827 8557
rect 4479 8520 9720 8548
rect 4479 8517 4491 8520
rect 4433 8511 4491 8517
rect 3053 8483 3111 8489
rect 3053 8480 3065 8483
rect 1964 8452 3065 8480
rect 1964 8424 1992 8452
rect 3053 8449 3065 8452
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8480 4123 8483
rect 4338 8480 4344 8492
rect 4111 8452 4344 8480
rect 4111 8449 4123 8452
rect 4065 8443 4123 8449
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 5626 8480 5632 8492
rect 5587 8452 5632 8480
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 7558 8480 7564 8492
rect 5859 8452 7564 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 8754 8440 8760 8492
rect 8812 8480 8818 8492
rect 8812 8452 8857 8480
rect 9232 8452 9628 8480
rect 8812 8440 8818 8452
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 1946 8412 1952 8424
rect 1719 8384 1952 8412
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 2225 8415 2283 8421
rect 2225 8381 2237 8415
rect 2271 8412 2283 8415
rect 2314 8412 2320 8424
rect 2271 8384 2320 8412
rect 2271 8381 2283 8384
rect 2225 8375 2283 8381
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 2682 8412 2688 8424
rect 2643 8384 2688 8412
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 3510 8372 3516 8424
rect 3568 8412 3574 8424
rect 7101 8415 7159 8421
rect 3568 8384 4016 8412
rect 3568 8372 3574 8384
rect 3988 8353 4016 8384
rect 7101 8381 7113 8415
rect 7147 8412 7159 8415
rect 8294 8412 8300 8424
rect 7147 8384 8300 8412
rect 7147 8381 7159 8384
rect 7101 8375 7159 8381
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 9232 8412 9260 8452
rect 8496 8384 9260 8412
rect 9309 8415 9367 8421
rect 3881 8347 3939 8353
rect 3881 8313 3893 8347
rect 3927 8313 3939 8347
rect 3881 8307 3939 8313
rect 3973 8347 4031 8353
rect 3973 8313 3985 8347
rect 4019 8313 4031 8347
rect 3973 8307 4031 8313
rect 5537 8347 5595 8353
rect 5537 8313 5549 8347
rect 5583 8344 5595 8347
rect 8202 8344 8208 8356
rect 5583 8316 8208 8344
rect 5583 8313 5595 8316
rect 5537 8307 5595 8313
rect 3896 8276 3924 8307
rect 8202 8304 8208 8316
rect 8260 8344 8266 8356
rect 8496 8344 8524 8384
rect 9309 8381 9321 8415
rect 9355 8412 9367 8415
rect 9398 8412 9404 8424
rect 9355 8384 9404 8412
rect 9355 8381 9367 8384
rect 9309 8375 9367 8381
rect 9398 8372 9404 8384
rect 9456 8372 9462 8424
rect 9600 8421 9628 8452
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8381 9643 8415
rect 9692 8412 9720 8520
rect 9769 8517 9781 8551
rect 9815 8548 9827 8551
rect 12434 8548 12440 8560
rect 9815 8520 12440 8548
rect 9815 8517 9827 8520
rect 9769 8511 9827 8517
rect 12434 8508 12440 8520
rect 12492 8508 12498 8560
rect 10612 8452 12480 8480
rect 10612 8421 10640 8452
rect 10597 8415 10655 8421
rect 10597 8412 10609 8415
rect 9692 8384 10609 8412
rect 9585 8375 9643 8381
rect 10597 8381 10609 8384
rect 10643 8381 10655 8415
rect 10597 8375 10655 8381
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8412 11207 8415
rect 11790 8412 11796 8424
rect 11195 8384 11796 8412
rect 11195 8381 11207 8384
rect 11149 8375 11207 8381
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 12066 8412 12072 8424
rect 12027 8384 12072 8412
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 12452 8421 12480 8452
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8381 12495 8415
rect 12544 8412 12572 8588
rect 12802 8576 12808 8628
rect 12860 8616 12866 8628
rect 12989 8619 13047 8625
rect 12989 8616 13001 8619
rect 12860 8588 13001 8616
rect 12860 8576 12866 8588
rect 12989 8585 13001 8588
rect 13035 8585 13047 8619
rect 12989 8579 13047 8585
rect 15654 8508 15660 8560
rect 15712 8548 15718 8560
rect 15841 8551 15899 8557
rect 15841 8548 15853 8551
rect 15712 8520 15853 8548
rect 15712 8508 15718 8520
rect 15841 8517 15853 8520
rect 15887 8517 15899 8551
rect 15841 8511 15899 8517
rect 15473 8483 15531 8489
rect 15473 8480 15485 8483
rect 14476 8452 15485 8480
rect 14476 8424 14504 8452
rect 15473 8449 15485 8452
rect 15519 8449 15531 8483
rect 17678 8480 17684 8492
rect 17639 8452 17684 8480
rect 15473 8443 15531 8449
rect 17678 8440 17684 8452
rect 17736 8440 17742 8492
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 12544 8384 12909 8412
rect 12437 8375 12495 8381
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 14458 8412 14464 8424
rect 14419 8384 14464 8412
rect 12897 8375 12955 8381
rect 14458 8372 14464 8384
rect 14516 8372 14522 8424
rect 15013 8415 15071 8421
rect 15013 8381 15025 8415
rect 15059 8412 15071 8415
rect 15378 8412 15384 8424
rect 15059 8384 15384 8412
rect 15059 8381 15071 8384
rect 15013 8375 15071 8381
rect 15378 8372 15384 8384
rect 15436 8372 15442 8424
rect 17313 8415 17371 8421
rect 17313 8381 17325 8415
rect 17359 8412 17371 8415
rect 17494 8412 17500 8424
rect 17359 8384 17500 8412
rect 17359 8381 17371 8384
rect 17313 8375 17371 8381
rect 17494 8372 17500 8384
rect 17552 8372 17558 8424
rect 17862 8412 17868 8424
rect 17775 8384 17868 8412
rect 17862 8372 17868 8384
rect 17920 8372 17926 8424
rect 8260 8316 8524 8344
rect 8573 8347 8631 8353
rect 8260 8304 8266 8316
rect 8573 8313 8585 8347
rect 8619 8344 8631 8347
rect 10410 8344 10416 8356
rect 8619 8316 10416 8344
rect 8619 8313 8631 8316
rect 8573 8307 8631 8313
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 14921 8347 14979 8353
rect 14921 8313 14933 8347
rect 14967 8344 14979 8347
rect 16482 8344 16488 8356
rect 14967 8316 16488 8344
rect 14967 8313 14979 8316
rect 14921 8307 14979 8313
rect 4338 8276 4344 8288
rect 3896 8248 4344 8276
rect 4338 8236 4344 8248
rect 4396 8276 4402 8288
rect 4706 8276 4712 8288
rect 4396 8248 4712 8276
rect 4396 8236 4402 8248
rect 4706 8236 4712 8248
rect 4764 8236 4770 8288
rect 6917 8279 6975 8285
rect 6917 8245 6929 8279
rect 6963 8276 6975 8279
rect 7282 8276 7288 8288
rect 6963 8248 7288 8276
rect 6963 8245 6975 8248
rect 6917 8239 6975 8245
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 8110 8276 8116 8288
rect 8071 8248 8116 8276
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 8478 8276 8484 8288
rect 8439 8248 8484 8276
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 15856 8285 15884 8316
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 17880 8344 17908 8372
rect 16632 8316 17908 8344
rect 16632 8304 16638 8316
rect 15841 8279 15899 8285
rect 15841 8245 15853 8279
rect 15887 8245 15899 8279
rect 15841 8239 15899 8245
rect 1104 8186 19044 8208
rect 1104 8134 6962 8186
rect 7014 8134 7026 8186
rect 7078 8134 7090 8186
rect 7142 8134 7154 8186
rect 7206 8134 12942 8186
rect 12994 8134 13006 8186
rect 13058 8134 13070 8186
rect 13122 8134 13134 8186
rect 13186 8134 19044 8186
rect 1104 8112 19044 8134
rect 2682 8072 2688 8084
rect 2643 8044 2688 8072
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 11977 8075 12035 8081
rect 11977 8041 11989 8075
rect 12023 8072 12035 8075
rect 12066 8072 12072 8084
rect 12023 8044 12072 8072
rect 12023 8041 12035 8044
rect 11977 8035 12035 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 13265 8075 13323 8081
rect 13265 8041 13277 8075
rect 13311 8072 13323 8075
rect 13354 8072 13360 8084
rect 13311 8044 13360 8072
rect 13311 8041 13323 8044
rect 13265 8035 13323 8041
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 17589 8075 17647 8081
rect 17589 8041 17601 8075
rect 17635 8072 17647 8075
rect 17678 8072 17684 8084
rect 17635 8044 17684 8072
rect 17635 8041 17647 8044
rect 17589 8035 17647 8041
rect 17678 8032 17684 8044
rect 17736 8032 17742 8084
rect 2590 7964 2596 8016
rect 2648 8004 2654 8016
rect 3145 8007 3203 8013
rect 3145 8004 3157 8007
rect 2648 7976 3157 8004
rect 2648 7964 2654 7976
rect 3145 7973 3157 7976
rect 3191 7973 3203 8007
rect 3145 7967 3203 7973
rect 4433 8007 4491 8013
rect 4433 7973 4445 8007
rect 4479 7973 4491 8007
rect 4614 8004 4620 8016
rect 4575 7976 4620 8004
rect 4433 7967 4491 7973
rect 2314 7896 2320 7948
rect 2372 7936 2378 7948
rect 2501 7939 2559 7945
rect 2501 7936 2513 7939
rect 2372 7908 2513 7936
rect 2372 7896 2378 7908
rect 2501 7905 2513 7908
rect 2547 7905 2559 7939
rect 4448 7936 4476 7967
rect 4614 7964 4620 7976
rect 4672 7964 4678 8016
rect 7469 8007 7527 8013
rect 7469 7973 7481 8007
rect 7515 8004 7527 8007
rect 7742 8004 7748 8016
rect 7515 7976 7748 8004
rect 7515 7973 7527 7976
rect 7469 7967 7527 7973
rect 7742 7964 7748 7976
rect 7800 7964 7806 8016
rect 11149 8007 11207 8013
rect 11149 8004 11161 8007
rect 9508 7976 11161 8004
rect 7282 7936 7288 7948
rect 2501 7899 2559 7905
rect 2608 7908 4476 7936
rect 7243 7908 7288 7936
rect 2406 7828 2412 7880
rect 2464 7868 2470 7880
rect 2608 7868 2636 7908
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 9306 7896 9312 7948
rect 9364 7936 9370 7948
rect 9508 7945 9536 7976
rect 11149 7973 11161 7976
rect 11195 8004 11207 8007
rect 12250 8004 12256 8016
rect 11195 7976 12256 8004
rect 11195 7973 11207 7976
rect 11149 7967 11207 7973
rect 12250 7964 12256 7976
rect 12308 7964 12314 8016
rect 9493 7939 9551 7945
rect 9493 7936 9505 7939
rect 9364 7908 9505 7936
rect 9364 7896 9370 7908
rect 9493 7905 9505 7908
rect 9539 7905 9551 7939
rect 9674 7936 9680 7948
rect 9635 7908 9680 7936
rect 9493 7899 9551 7905
rect 9674 7896 9680 7908
rect 9732 7936 9738 7948
rect 10965 7939 11023 7945
rect 10965 7936 10977 7939
rect 9732 7908 10977 7936
rect 9732 7896 9738 7908
rect 10965 7905 10977 7908
rect 11011 7905 11023 7939
rect 11790 7936 11796 7948
rect 11751 7908 11796 7936
rect 10965 7899 11023 7905
rect 11790 7896 11796 7908
rect 11848 7896 11854 7948
rect 12618 7896 12624 7948
rect 12676 7936 12682 7948
rect 12897 7939 12955 7945
rect 12897 7936 12909 7939
rect 12676 7908 12909 7936
rect 12676 7896 12682 7908
rect 12897 7905 12909 7908
rect 12943 7905 12955 7939
rect 12897 7899 12955 7905
rect 16761 7939 16819 7945
rect 16761 7905 16773 7939
rect 16807 7936 16819 7939
rect 17405 7939 17463 7945
rect 17405 7936 17417 7939
rect 16807 7908 17417 7936
rect 16807 7905 16819 7908
rect 16761 7899 16819 7905
rect 17405 7905 17417 7908
rect 17451 7905 17463 7939
rect 17405 7899 17463 7905
rect 4338 7868 4344 7880
rect 2464 7840 2636 7868
rect 4299 7840 4344 7868
rect 2464 7828 2470 7840
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 15746 7828 15752 7880
rect 15804 7868 15810 7880
rect 16393 7871 16451 7877
rect 16393 7868 16405 7871
rect 15804 7840 16405 7868
rect 15804 7828 15810 7840
rect 16393 7837 16405 7840
rect 16439 7837 16451 7871
rect 16393 7831 16451 7837
rect 4893 7803 4951 7809
rect 4893 7769 4905 7803
rect 4939 7800 4951 7803
rect 9766 7800 9772 7812
rect 4939 7772 9772 7800
rect 4939 7769 4951 7772
rect 4893 7763 4951 7769
rect 9766 7760 9772 7772
rect 9824 7760 9830 7812
rect 13265 7803 13323 7809
rect 13265 7769 13277 7803
rect 13311 7800 13323 7803
rect 13630 7800 13636 7812
rect 13311 7772 13636 7800
rect 13311 7769 13323 7772
rect 13265 7763 13323 7769
rect 13630 7760 13636 7772
rect 13688 7760 13694 7812
rect 3234 7732 3240 7744
rect 3195 7704 3240 7732
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 9490 7732 9496 7744
rect 9451 7704 9496 7732
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 9674 7692 9680 7744
rect 9732 7732 9738 7744
rect 9861 7735 9919 7741
rect 9861 7732 9873 7735
rect 9732 7704 9873 7732
rect 9732 7692 9738 7704
rect 9861 7701 9873 7704
rect 9907 7701 9919 7735
rect 9861 7695 9919 7701
rect 11333 7735 11391 7741
rect 11333 7701 11345 7735
rect 11379 7732 11391 7735
rect 12066 7732 12072 7744
rect 11379 7704 12072 7732
rect 11379 7701 11391 7704
rect 11333 7695 11391 7701
rect 12066 7692 12072 7704
rect 12124 7692 12130 7744
rect 16298 7692 16304 7744
rect 16356 7732 16362 7744
rect 16761 7735 16819 7741
rect 16761 7732 16773 7735
rect 16356 7704 16773 7732
rect 16356 7692 16362 7704
rect 16761 7701 16773 7704
rect 16807 7701 16819 7735
rect 16761 7695 16819 7701
rect 1104 7642 19044 7664
rect 1104 7590 3972 7642
rect 4024 7590 4036 7642
rect 4088 7590 4100 7642
rect 4152 7590 4164 7642
rect 4216 7590 9952 7642
rect 10004 7590 10016 7642
rect 10068 7590 10080 7642
rect 10132 7590 10144 7642
rect 10196 7590 15932 7642
rect 15984 7590 15996 7642
rect 16048 7590 16060 7642
rect 16112 7590 16124 7642
rect 16176 7590 19044 7642
rect 1104 7568 19044 7590
rect 13354 7528 13360 7540
rect 13315 7500 13360 7528
rect 13354 7488 13360 7500
rect 13412 7488 13418 7540
rect 16298 7528 16304 7540
rect 16259 7500 16304 7528
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 11057 7463 11115 7469
rect 11057 7429 11069 7463
rect 11103 7460 11115 7463
rect 11790 7460 11796 7472
rect 11103 7432 11796 7460
rect 11103 7429 11115 7432
rect 11057 7423 11115 7429
rect 11790 7420 11796 7432
rect 11848 7420 11854 7472
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7392 5503 7395
rect 5491 7364 7052 7392
rect 5491 7361 5503 7364
rect 5445 7355 5503 7361
rect 1762 7324 1768 7336
rect 1723 7296 1768 7324
rect 1762 7284 1768 7296
rect 1820 7284 1826 7336
rect 2314 7324 2320 7336
rect 2275 7296 2320 7324
rect 2314 7284 2320 7296
rect 2372 7284 2378 7336
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7293 4031 7327
rect 3973 7287 4031 7293
rect 4249 7327 4307 7333
rect 4249 7293 4261 7327
rect 4295 7324 4307 7327
rect 4522 7324 4528 7336
rect 4295 7296 4528 7324
rect 4295 7293 4307 7296
rect 4249 7287 4307 7293
rect 2225 7259 2283 7265
rect 2225 7225 2237 7259
rect 2271 7256 2283 7259
rect 3326 7256 3332 7268
rect 2271 7228 3332 7256
rect 2271 7225 2283 7228
rect 2225 7219 2283 7225
rect 3326 7216 3332 7228
rect 3384 7216 3390 7268
rect 2130 7148 2136 7200
rect 2188 7188 2194 7200
rect 3789 7191 3847 7197
rect 3789 7188 3801 7191
rect 2188 7160 3801 7188
rect 2188 7148 2194 7160
rect 3789 7157 3801 7160
rect 3835 7157 3847 7191
rect 3988 7188 4016 7287
rect 4522 7284 4528 7296
rect 4580 7284 4586 7336
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7324 5779 7327
rect 5994 7324 6000 7336
rect 5767 7296 6000 7324
rect 5767 7293 5779 7296
rect 5721 7287 5779 7293
rect 5994 7284 6000 7296
rect 6052 7284 6058 7336
rect 7024 7333 7052 7364
rect 7009 7327 7067 7333
rect 7009 7293 7021 7327
rect 7055 7324 7067 7327
rect 7374 7324 7380 7336
rect 7055 7296 7380 7324
rect 7055 7293 7067 7296
rect 7009 7287 7067 7293
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 7558 7324 7564 7336
rect 7519 7296 7564 7324
rect 7558 7284 7564 7296
rect 7616 7324 7622 7336
rect 8754 7324 8760 7336
rect 7616 7296 8760 7324
rect 7616 7284 7622 7296
rect 8754 7284 8760 7296
rect 8812 7284 8818 7336
rect 12618 7284 12624 7336
rect 12676 7324 12682 7336
rect 12805 7327 12863 7333
rect 12805 7324 12817 7327
rect 12676 7296 12817 7324
rect 12676 7284 12682 7296
rect 12805 7293 12817 7296
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 13357 7327 13415 7333
rect 13357 7293 13369 7327
rect 13403 7324 13415 7327
rect 13446 7324 13452 7336
rect 13403 7296 13452 7324
rect 13403 7293 13415 7296
rect 13357 7287 13415 7293
rect 13446 7284 13452 7296
rect 13504 7284 13510 7336
rect 14550 7284 14556 7336
rect 14608 7324 14614 7336
rect 15746 7324 15752 7336
rect 14608 7296 15752 7324
rect 14608 7284 14614 7296
rect 15746 7284 15752 7296
rect 15804 7284 15810 7336
rect 16301 7327 16359 7333
rect 16301 7293 16313 7327
rect 16347 7324 16359 7327
rect 16574 7324 16580 7336
rect 16347 7296 16580 7324
rect 16347 7293 16359 7296
rect 16301 7287 16359 7293
rect 16574 7284 16580 7296
rect 16632 7284 16638 7336
rect 4157 7259 4215 7265
rect 4157 7225 4169 7259
rect 4203 7256 4215 7259
rect 5166 7256 5172 7268
rect 4203 7228 5172 7256
rect 4203 7225 4215 7228
rect 4157 7219 4215 7225
rect 5166 7216 5172 7228
rect 5224 7216 5230 7268
rect 5902 7256 5908 7268
rect 5863 7228 5908 7256
rect 5902 7216 5908 7228
rect 5960 7216 5966 7268
rect 9122 7216 9128 7268
rect 9180 7256 9186 7268
rect 10873 7259 10931 7265
rect 10873 7256 10885 7259
rect 9180 7228 10885 7256
rect 9180 7216 9186 7228
rect 10873 7225 10885 7228
rect 10919 7225 10931 7259
rect 10873 7219 10931 7225
rect 6822 7188 6828 7200
rect 3988 7160 6828 7188
rect 3789 7151 3847 7157
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 7926 7188 7932 7200
rect 7887 7160 7932 7188
rect 7926 7148 7932 7160
rect 7984 7148 7990 7200
rect 8570 7148 8576 7200
rect 8628 7188 8634 7200
rect 8665 7191 8723 7197
rect 8665 7188 8677 7191
rect 8628 7160 8677 7188
rect 8628 7148 8634 7160
rect 8665 7157 8677 7160
rect 8711 7157 8723 7191
rect 8665 7151 8723 7157
rect 8754 7148 8760 7200
rect 8812 7188 8818 7200
rect 8812 7160 8857 7188
rect 8812 7148 8818 7160
rect 1104 7098 19044 7120
rect 1104 7046 6962 7098
rect 7014 7046 7026 7098
rect 7078 7046 7090 7098
rect 7142 7046 7154 7098
rect 7206 7046 12942 7098
rect 12994 7046 13006 7098
rect 13058 7046 13070 7098
rect 13122 7046 13134 7098
rect 13186 7046 19044 7098
rect 1104 7024 19044 7046
rect 2130 6984 2136 6996
rect 2091 6956 2136 6984
rect 2130 6944 2136 6956
rect 2188 6944 2194 6996
rect 4338 6944 4344 6996
rect 4396 6984 4402 6996
rect 7558 6984 7564 6996
rect 4396 6956 7564 6984
rect 4396 6944 4402 6956
rect 1578 6876 1584 6928
rect 1636 6916 1642 6928
rect 4356 6916 4384 6944
rect 4724 6925 4752 6956
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 12066 6984 12072 6996
rect 12027 6956 12072 6984
rect 12066 6944 12072 6956
rect 12124 6944 12130 6996
rect 13173 6987 13231 6993
rect 13173 6953 13185 6987
rect 13219 6984 13231 6987
rect 13354 6984 13360 6996
rect 13219 6956 13360 6984
rect 13219 6953 13231 6956
rect 13173 6947 13231 6953
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 13630 6984 13636 6996
rect 13591 6956 13636 6984
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 1636 6888 4384 6916
rect 4709 6919 4767 6925
rect 1636 6876 1642 6888
rect 1578 6740 1584 6792
rect 1636 6780 1642 6792
rect 2424 6789 2452 6888
rect 4709 6885 4721 6919
rect 4755 6885 4767 6919
rect 4709 6879 4767 6885
rect 4801 6919 4859 6925
rect 4801 6885 4813 6919
rect 4847 6885 4859 6919
rect 4982 6916 4988 6928
rect 4943 6888 4988 6916
rect 4801 6879 4859 6885
rect 3234 6808 3240 6860
rect 3292 6848 3298 6860
rect 3329 6851 3387 6857
rect 3329 6848 3341 6851
rect 3292 6820 3341 6848
rect 3292 6808 3298 6820
rect 3329 6817 3341 6820
rect 3375 6817 3387 6851
rect 4816 6848 4844 6879
rect 4982 6876 4988 6888
rect 5040 6876 5046 6928
rect 15105 6919 15163 6925
rect 15105 6885 15117 6919
rect 15151 6916 15163 6919
rect 15470 6916 15476 6928
rect 15151 6888 15476 6916
rect 15151 6885 15163 6888
rect 15105 6879 15163 6885
rect 15470 6876 15476 6888
rect 15528 6876 15534 6928
rect 16298 6876 16304 6928
rect 16356 6916 16362 6928
rect 16485 6919 16543 6925
rect 16485 6916 16497 6919
rect 16356 6888 16497 6916
rect 16356 6876 16362 6888
rect 16485 6885 16497 6888
rect 16531 6885 16543 6919
rect 16485 6879 16543 6885
rect 4890 6848 4896 6860
rect 4816 6820 4896 6848
rect 3329 6811 3387 6817
rect 4890 6808 4896 6820
rect 4948 6808 4954 6860
rect 6181 6851 6239 6857
rect 6181 6817 6193 6851
rect 6227 6848 6239 6851
rect 6641 6851 6699 6857
rect 6641 6848 6653 6851
rect 6227 6820 6653 6848
rect 6227 6817 6239 6820
rect 6181 6811 6239 6817
rect 6641 6817 6653 6820
rect 6687 6817 6699 6851
rect 6641 6811 6699 6817
rect 7374 6808 7380 6860
rect 7432 6848 7438 6860
rect 7561 6851 7619 6857
rect 7561 6848 7573 6851
rect 7432 6820 7573 6848
rect 7432 6808 7438 6820
rect 7561 6817 7573 6820
rect 7607 6817 7619 6851
rect 7561 6811 7619 6817
rect 8021 6851 8079 6857
rect 8021 6817 8033 6851
rect 8067 6848 8079 6851
rect 8110 6848 8116 6860
rect 8067 6820 8116 6848
rect 8067 6817 8079 6820
rect 8021 6811 8079 6817
rect 8110 6808 8116 6820
rect 8168 6808 8174 6860
rect 8573 6851 8631 6857
rect 8573 6817 8585 6851
rect 8619 6848 8631 6851
rect 9306 6848 9312 6860
rect 8619 6820 9312 6848
rect 8619 6817 8631 6820
rect 8573 6811 8631 6817
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 9953 6851 10011 6857
rect 9953 6848 9965 6851
rect 9824 6820 9965 6848
rect 9824 6808 9830 6820
rect 9953 6817 9965 6820
rect 9999 6817 10011 6851
rect 9953 6811 10011 6817
rect 10597 6851 10655 6857
rect 10597 6817 10609 6851
rect 10643 6817 10655 6851
rect 10870 6848 10876 6860
rect 10831 6820 10876 6848
rect 10597 6811 10655 6817
rect 2225 6783 2283 6789
rect 2225 6780 2237 6783
rect 1636 6752 2237 6780
rect 1636 6740 1642 6752
rect 2225 6749 2237 6752
rect 2271 6749 2283 6783
rect 2225 6743 2283 6749
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6749 2467 6783
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2409 6743 2467 6749
rect 2746 6752 2973 6780
rect 1762 6712 1768 6724
rect 1675 6684 1768 6712
rect 1762 6672 1768 6684
rect 1820 6712 1826 6724
rect 2746 6712 2774 6752
rect 2961 6749 2973 6752
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6780 6975 6783
rect 8294 6780 8300 6792
rect 6963 6752 8300 6780
rect 6963 6749 6975 6752
rect 6917 6743 6975 6749
rect 8294 6740 8300 6752
rect 8352 6780 8358 6792
rect 9122 6780 9128 6792
rect 8352 6752 9128 6780
rect 8352 6740 8358 6752
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 9324 6780 9352 6808
rect 10612 6780 10640 6811
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 11900 6820 12434 6848
rect 11790 6780 11796 6792
rect 9324 6752 10640 6780
rect 11751 6752 11796 6780
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 1820 6684 2774 6712
rect 5261 6715 5319 6721
rect 1820 6672 1826 6684
rect 5261 6681 5273 6715
rect 5307 6712 5319 6715
rect 11900 6712 11928 6820
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6749 12035 6783
rect 12406 6780 12434 6820
rect 13446 6808 13452 6860
rect 13504 6848 13510 6860
rect 13817 6851 13875 6857
rect 13817 6848 13829 6851
rect 13504 6820 13829 6848
rect 13504 6808 13510 6820
rect 13817 6817 13829 6820
rect 13863 6848 13875 6851
rect 14826 6848 14832 6860
rect 13863 6820 14832 6848
rect 13863 6817 13875 6820
rect 13817 6811 13875 6817
rect 14826 6808 14832 6820
rect 14884 6808 14890 6860
rect 14918 6808 14924 6860
rect 14976 6848 14982 6860
rect 15197 6851 15255 6857
rect 15197 6848 15209 6851
rect 14976 6820 15209 6848
rect 14976 6808 14982 6820
rect 15197 6817 15209 6820
rect 15243 6817 15255 6851
rect 18322 6848 18328 6860
rect 18283 6820 18328 6848
rect 15197 6811 15255 6817
rect 18322 6808 18328 6820
rect 18380 6808 18386 6860
rect 14550 6780 14556 6792
rect 12406 6752 14556 6780
rect 11977 6743 12035 6749
rect 5307 6684 11928 6712
rect 11992 6712 12020 6743
rect 14550 6740 14556 6752
rect 14608 6740 14614 6792
rect 14642 6740 14648 6792
rect 14700 6780 14706 6792
rect 15289 6783 15347 6789
rect 15289 6780 15301 6783
rect 14700 6752 15301 6780
rect 14700 6740 14706 6752
rect 15289 6749 15301 6752
rect 15335 6749 15347 6783
rect 15289 6743 15347 6749
rect 16546 6752 18184 6780
rect 16546 6712 16574 6752
rect 18156 6721 18184 6752
rect 11992 6684 16574 6712
rect 18141 6715 18199 6721
rect 5307 6681 5319 6684
rect 5261 6675 5319 6681
rect 18141 6681 18153 6715
rect 18187 6681 18199 6715
rect 18141 6675 18199 6681
rect 3326 6644 3332 6656
rect 3287 6616 3332 6644
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 8570 6644 8576 6656
rect 8531 6616 8576 6644
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 12342 6604 12348 6656
rect 12400 6644 12406 6656
rect 12437 6647 12495 6653
rect 12437 6644 12449 6647
rect 12400 6616 12449 6644
rect 12400 6604 12406 6616
rect 12437 6613 12449 6616
rect 12483 6613 12495 6647
rect 12437 6607 12495 6613
rect 12710 6604 12716 6656
rect 12768 6644 12774 6656
rect 13081 6647 13139 6653
rect 13081 6644 13093 6647
rect 12768 6616 13093 6644
rect 12768 6604 12774 6616
rect 13081 6613 13093 6616
rect 13127 6613 13139 6647
rect 14734 6644 14740 6656
rect 14695 6616 14740 6644
rect 13081 6607 13139 6613
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 14826 6604 14832 6656
rect 14884 6644 14890 6656
rect 16393 6647 16451 6653
rect 16393 6644 16405 6647
rect 14884 6616 16405 6644
rect 14884 6604 14890 6616
rect 16393 6613 16405 6616
rect 16439 6613 16451 6647
rect 16393 6607 16451 6613
rect 1104 6554 19044 6576
rect 1104 6502 3972 6554
rect 4024 6502 4036 6554
rect 4088 6502 4100 6554
rect 4152 6502 4164 6554
rect 4216 6502 9952 6554
rect 10004 6502 10016 6554
rect 10068 6502 10080 6554
rect 10132 6502 10144 6554
rect 10196 6502 15932 6554
rect 15984 6502 15996 6554
rect 16048 6502 16060 6554
rect 16112 6502 16124 6554
rect 16176 6502 19044 6554
rect 1104 6480 19044 6502
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 14734 6440 14740 6452
rect 2746 6412 14740 6440
rect 2498 6332 2504 6384
rect 2556 6372 2562 6384
rect 2746 6372 2774 6412
rect 14734 6400 14740 6412
rect 14792 6400 14798 6452
rect 12710 6372 12716 6384
rect 2556 6344 2774 6372
rect 12671 6344 12716 6372
rect 2556 6332 2562 6344
rect 12710 6332 12716 6344
rect 12768 6332 12774 6384
rect 16390 6372 16396 6384
rect 16040 6344 16396 6372
rect 4065 6307 4123 6313
rect 4065 6273 4077 6307
rect 4111 6304 4123 6307
rect 4430 6304 4436 6316
rect 4111 6276 4436 6304
rect 4111 6273 4123 6276
rect 4065 6267 4123 6273
rect 4430 6264 4436 6276
rect 4488 6264 4494 6316
rect 8754 6304 8760 6316
rect 7944 6276 8760 6304
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 6638 6196 6644 6248
rect 6696 6236 6702 6248
rect 7944 6245 7972 6276
rect 8754 6264 8760 6276
rect 8812 6264 8818 6316
rect 10873 6307 10931 6313
rect 10873 6304 10885 6307
rect 9324 6276 10885 6304
rect 9324 6248 9352 6276
rect 10873 6273 10885 6276
rect 10919 6273 10931 6307
rect 14642 6304 14648 6316
rect 14603 6276 14648 6304
rect 10873 6267 10931 6273
rect 14642 6264 14648 6276
rect 14700 6264 14706 6316
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 6696 6208 7021 6236
rect 6696 6196 6702 6208
rect 7009 6205 7021 6208
rect 7055 6205 7067 6239
rect 7009 6199 7067 6205
rect 7929 6239 7987 6245
rect 7929 6205 7941 6239
rect 7975 6205 7987 6239
rect 8386 6236 8392 6248
rect 8347 6208 8392 6236
rect 7929 6199 7987 6205
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 9122 6236 9128 6248
rect 9083 6208 9128 6236
rect 9122 6196 9128 6208
rect 9180 6196 9186 6248
rect 9306 6236 9312 6248
rect 9267 6208 9312 6236
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 9766 6196 9772 6248
rect 9824 6236 9830 6248
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 9824 6208 10241 6236
rect 9824 6196 9830 6208
rect 10229 6205 10241 6208
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 10778 6196 10784 6248
rect 10836 6236 10842 6248
rect 10965 6239 11023 6245
rect 10965 6236 10977 6239
rect 10836 6208 10977 6236
rect 10836 6196 10842 6208
rect 10965 6205 10977 6208
rect 11011 6205 11023 6239
rect 12342 6236 12348 6248
rect 12303 6208 12348 6236
rect 10965 6199 11023 6205
rect 12342 6196 12348 6208
rect 12400 6196 12406 6248
rect 14829 6239 14887 6245
rect 14829 6236 14841 6239
rect 12544 6208 14841 6236
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 4525 6171 4583 6177
rect 4525 6168 4537 6171
rect 4120 6140 4537 6168
rect 4120 6128 4126 6140
rect 4525 6137 4537 6140
rect 4571 6137 4583 6171
rect 4525 6131 4583 6137
rect 4617 6171 4675 6177
rect 4617 6137 4629 6171
rect 4663 6168 4675 6171
rect 5077 6171 5135 6177
rect 5077 6168 5089 6171
rect 4663 6140 5089 6168
rect 4663 6137 4675 6140
rect 4617 6131 4675 6137
rect 5077 6137 5089 6140
rect 5123 6137 5135 6171
rect 5077 6131 5135 6137
rect 7653 6171 7711 6177
rect 7653 6137 7665 6171
rect 7699 6168 7711 6171
rect 9140 6168 9168 6196
rect 7699 6140 9168 6168
rect 7699 6137 7711 6140
rect 7653 6131 7711 6137
rect 5258 6100 5264 6112
rect 5219 6072 5264 6100
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 12544 6100 12572 6208
rect 14829 6205 14841 6208
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 15013 6239 15071 6245
rect 15013 6205 15025 6239
rect 15059 6205 15071 6239
rect 15013 6199 15071 6205
rect 15289 6239 15347 6245
rect 15289 6205 15301 6239
rect 15335 6236 15347 6239
rect 15841 6239 15899 6245
rect 15841 6236 15853 6239
rect 15335 6208 15853 6236
rect 15335 6205 15347 6208
rect 15289 6199 15347 6205
rect 15841 6205 15853 6208
rect 15887 6236 15899 6239
rect 15930 6236 15936 6248
rect 15887 6208 15936 6236
rect 15887 6205 15899 6208
rect 15841 6199 15899 6205
rect 12710 6100 12716 6112
rect 9548 6072 12572 6100
rect 12671 6072 12716 6100
rect 9548 6060 9554 6072
rect 12710 6060 12716 6072
rect 12768 6060 12774 6112
rect 14844 6100 14872 6199
rect 15028 6168 15056 6199
rect 15930 6196 15936 6208
rect 15988 6196 15994 6248
rect 16040 6245 16068 6344
rect 16390 6332 16396 6344
rect 16448 6372 16454 6384
rect 18046 6372 18052 6384
rect 16448 6344 18052 6372
rect 16448 6332 16454 6344
rect 18046 6332 18052 6344
rect 18104 6332 18110 6384
rect 16025 6239 16083 6245
rect 16025 6205 16037 6239
rect 16071 6205 16083 6239
rect 16025 6199 16083 6205
rect 16209 6239 16267 6245
rect 16209 6205 16221 6239
rect 16255 6236 16267 6239
rect 17126 6236 17132 6248
rect 16255 6208 17132 6236
rect 16255 6205 16267 6208
rect 16209 6199 16267 6205
rect 16040 6168 16068 6199
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 15028 6140 16068 6168
rect 15562 6100 15568 6112
rect 14844 6072 15568 6100
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 15838 6100 15844 6112
rect 15799 6072 15844 6100
rect 15838 6060 15844 6072
rect 15896 6060 15902 6112
rect 1104 6010 19044 6032
rect 1104 5958 6962 6010
rect 7014 5958 7026 6010
rect 7078 5958 7090 6010
rect 7142 5958 7154 6010
rect 7206 5958 12942 6010
rect 12994 5958 13006 6010
rect 13058 5958 13070 6010
rect 13122 5958 13134 6010
rect 13186 5958 19044 6010
rect 1104 5936 19044 5958
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 5629 5899 5687 5905
rect 5629 5896 5641 5899
rect 5316 5868 5641 5896
rect 5316 5856 5322 5868
rect 5629 5865 5641 5868
rect 5675 5865 5687 5899
rect 6638 5896 6644 5908
rect 6599 5868 6644 5896
rect 5629 5859 5687 5865
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 6822 5856 6828 5908
rect 6880 5896 6886 5908
rect 7009 5899 7067 5905
rect 7009 5896 7021 5899
rect 6880 5868 7021 5896
rect 6880 5856 6886 5868
rect 7009 5865 7021 5868
rect 7055 5865 7067 5899
rect 8570 5896 8576 5908
rect 8531 5868 8576 5896
rect 7009 5859 7067 5865
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 10778 5896 10784 5908
rect 10739 5868 10784 5896
rect 10778 5856 10784 5868
rect 10836 5856 10842 5908
rect 14185 5899 14243 5905
rect 14185 5865 14197 5899
rect 14231 5896 14243 5899
rect 15013 5899 15071 5905
rect 15013 5896 15025 5899
rect 14231 5868 15025 5896
rect 14231 5865 14243 5868
rect 14185 5859 14243 5865
rect 15013 5865 15025 5868
rect 15059 5865 15071 5899
rect 15470 5896 15476 5908
rect 15431 5868 15476 5896
rect 15013 5859 15071 5865
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 17126 5896 17132 5908
rect 17087 5868 17132 5896
rect 17126 5856 17132 5868
rect 17184 5856 17190 5908
rect 3050 5828 3056 5840
rect 3011 5800 3056 5828
rect 3050 5788 3056 5800
rect 3108 5788 3114 5840
rect 4062 5828 4068 5840
rect 3252 5800 4068 5828
rect 3252 5772 3280 5800
rect 4062 5788 4068 5800
rect 4120 5828 4126 5840
rect 4893 5831 4951 5837
rect 4893 5828 4905 5831
rect 4120 5800 4905 5828
rect 4120 5788 4126 5800
rect 4893 5797 4905 5800
rect 4939 5797 4951 5831
rect 4893 5791 4951 5797
rect 12529 5831 12587 5837
rect 12529 5797 12541 5831
rect 12575 5828 12587 5831
rect 12710 5828 12716 5840
rect 12575 5800 12716 5828
rect 12575 5797 12587 5800
rect 12529 5791 12587 5797
rect 12710 5788 12716 5800
rect 12768 5788 12774 5840
rect 15838 5828 15844 5840
rect 14936 5800 15844 5828
rect 3234 5760 3240 5772
rect 3195 5732 3240 5760
rect 3234 5720 3240 5732
rect 3292 5720 3298 5772
rect 4249 5763 4307 5769
rect 4249 5729 4261 5763
rect 4295 5760 4307 5763
rect 4430 5760 4436 5772
rect 4295 5732 4436 5760
rect 4295 5729 4307 5732
rect 4249 5723 4307 5729
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 5166 5760 5172 5772
rect 5127 5732 5172 5760
rect 5166 5720 5172 5732
rect 5224 5720 5230 5772
rect 5442 5720 5448 5772
rect 5500 5760 5506 5772
rect 5997 5763 6055 5769
rect 5997 5760 6009 5763
rect 5500 5732 6009 5760
rect 5500 5720 5506 5732
rect 5997 5729 6009 5732
rect 6043 5729 6055 5763
rect 5997 5723 6055 5729
rect 7101 5763 7159 5769
rect 7101 5729 7113 5763
rect 7147 5760 7159 5763
rect 7147 5732 8064 5760
rect 7147 5729 7159 5732
rect 7101 5723 7159 5729
rect 5626 5692 5632 5704
rect 5587 5664 5632 5692
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 7285 5695 7343 5701
rect 7285 5661 7297 5695
rect 7331 5692 7343 5695
rect 7558 5692 7564 5704
rect 7331 5664 7564 5692
rect 7331 5661 7343 5664
rect 7285 5655 7343 5661
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 8036 5692 8064 5732
rect 8110 5720 8116 5772
rect 8168 5760 8174 5772
rect 8205 5763 8263 5769
rect 8205 5760 8217 5763
rect 8168 5732 8217 5760
rect 8168 5720 8174 5732
rect 8205 5729 8217 5732
rect 8251 5729 8263 5763
rect 8205 5723 8263 5729
rect 9306 5720 9312 5772
rect 9364 5760 9370 5772
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9364 5732 9689 5760
rect 9364 5720 9370 5732
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 10502 5720 10508 5772
rect 10560 5760 10566 5772
rect 10689 5763 10747 5769
rect 10689 5760 10701 5763
rect 10560 5732 10701 5760
rect 10560 5720 10566 5732
rect 10689 5729 10701 5732
rect 10735 5729 10747 5763
rect 10689 5723 10747 5729
rect 12069 5763 12127 5769
rect 12069 5729 12081 5763
rect 12115 5760 12127 5763
rect 12342 5760 12348 5772
rect 12115 5732 12348 5760
rect 12115 5729 12127 5732
rect 12069 5723 12127 5729
rect 12342 5720 12348 5732
rect 12400 5720 12406 5772
rect 12621 5763 12679 5769
rect 12621 5729 12633 5763
rect 12667 5760 12679 5763
rect 13446 5760 13452 5772
rect 12667 5732 13452 5760
rect 12667 5729 12679 5732
rect 12621 5723 12679 5729
rect 13446 5720 13452 5732
rect 13504 5720 13510 5772
rect 14936 5701 14964 5800
rect 15838 5788 15844 5800
rect 15896 5788 15902 5840
rect 15930 5788 15936 5840
rect 15988 5828 15994 5840
rect 15988 5800 16528 5828
rect 15988 5788 15994 5800
rect 16500 5772 16528 5800
rect 15102 5760 15108 5772
rect 15063 5732 15108 5760
rect 15102 5720 15108 5732
rect 15160 5720 15166 5772
rect 15562 5720 15568 5772
rect 15620 5760 15626 5772
rect 16117 5763 16175 5769
rect 16117 5760 16129 5763
rect 15620 5732 16129 5760
rect 15620 5720 15626 5732
rect 16117 5729 16129 5732
rect 16163 5729 16175 5763
rect 16298 5760 16304 5772
rect 16259 5732 16304 5760
rect 16117 5723 16175 5729
rect 14921 5695 14979 5701
rect 8036 5664 14872 5692
rect 8573 5627 8631 5633
rect 8573 5593 8585 5627
rect 8619 5624 8631 5627
rect 9493 5627 9551 5633
rect 9493 5624 9505 5627
rect 8619 5596 9505 5624
rect 8619 5593 8631 5596
rect 8573 5587 8631 5593
rect 9493 5593 9505 5596
rect 9539 5593 9551 5627
rect 14844 5624 14872 5664
rect 14921 5661 14933 5695
rect 14967 5661 14979 5695
rect 14921 5655 14979 5661
rect 15654 5652 15660 5704
rect 15712 5692 15718 5704
rect 15933 5695 15991 5701
rect 15933 5692 15945 5695
rect 15712 5664 15945 5692
rect 15712 5652 15718 5664
rect 15933 5661 15945 5664
rect 15979 5661 15991 5695
rect 16132 5692 16160 5723
rect 16298 5720 16304 5732
rect 16356 5720 16362 5772
rect 16482 5760 16488 5772
rect 16443 5732 16488 5760
rect 16482 5720 16488 5732
rect 16540 5720 16546 5772
rect 17037 5763 17095 5769
rect 17037 5729 17049 5763
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 17052 5692 17080 5723
rect 16132 5664 17080 5692
rect 15933 5655 15991 5661
rect 14844 5596 16574 5624
rect 9493 5587 9551 5593
rect 5718 5516 5724 5568
rect 5776 5556 5782 5568
rect 14185 5559 14243 5565
rect 14185 5556 14197 5559
rect 5776 5528 14197 5556
rect 5776 5516 5782 5528
rect 14185 5525 14197 5528
rect 14231 5525 14243 5559
rect 16546 5556 16574 5596
rect 18138 5556 18144 5568
rect 16546 5528 18144 5556
rect 14185 5519 14243 5525
rect 18138 5516 18144 5528
rect 18196 5516 18202 5568
rect 1104 5466 19044 5488
rect 1104 5414 3972 5466
rect 4024 5414 4036 5466
rect 4088 5414 4100 5466
rect 4152 5414 4164 5466
rect 4216 5414 9952 5466
rect 10004 5414 10016 5466
rect 10068 5414 10080 5466
rect 10132 5414 10144 5466
rect 10196 5414 15932 5466
rect 15984 5414 15996 5466
rect 16048 5414 16060 5466
rect 16112 5414 16124 5466
rect 16176 5414 19044 5466
rect 1104 5392 19044 5414
rect 15013 5355 15071 5361
rect 15013 5321 15025 5355
rect 15059 5352 15071 5355
rect 15102 5352 15108 5364
rect 15059 5324 15108 5352
rect 15059 5321 15071 5324
rect 15013 5315 15071 5321
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 16298 5352 16304 5364
rect 16259 5324 16304 5352
rect 16298 5312 16304 5324
rect 16356 5352 16362 5364
rect 16356 5324 16574 5352
rect 16356 5312 16362 5324
rect 5442 5284 5448 5296
rect 4908 5256 5448 5284
rect 2742 5151 2800 5157
rect 2742 5117 2754 5151
rect 2788 5148 2800 5151
rect 3234 5148 3240 5160
rect 2788 5120 3240 5148
rect 2788 5117 2800 5120
rect 2742 5111 2800 5117
rect 3234 5108 3240 5120
rect 3292 5108 3298 5160
rect 3326 5108 3332 5160
rect 3384 5148 3390 5160
rect 4908 5157 4936 5256
rect 5442 5244 5448 5256
rect 5500 5244 5506 5296
rect 7193 5287 7251 5293
rect 7193 5253 7205 5287
rect 7239 5284 7251 5287
rect 8386 5284 8392 5296
rect 7239 5256 8392 5284
rect 7239 5253 7251 5256
rect 7193 5247 7251 5253
rect 8386 5244 8392 5256
rect 8444 5244 8450 5296
rect 10505 5287 10563 5293
rect 10505 5253 10517 5287
rect 10551 5284 10563 5287
rect 10965 5287 11023 5293
rect 10965 5284 10977 5287
rect 10551 5256 10977 5284
rect 10551 5253 10563 5256
rect 10505 5247 10563 5253
rect 10965 5253 10977 5256
rect 11011 5253 11023 5287
rect 10965 5247 11023 5253
rect 5258 5216 5264 5228
rect 5219 5188 5264 5216
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 15654 5216 15660 5228
rect 15615 5188 15660 5216
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 16546 5216 16574 5324
rect 17126 5244 17132 5296
rect 17184 5284 17190 5296
rect 17184 5256 17816 5284
rect 17184 5244 17190 5256
rect 17788 5225 17816 5256
rect 17773 5219 17831 5225
rect 16546 5188 17632 5216
rect 4893 5151 4951 5157
rect 3384 5120 3429 5148
rect 3384 5108 3390 5120
rect 4893 5117 4905 5151
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 5166 5108 5172 5160
rect 5224 5148 5230 5160
rect 5445 5151 5503 5157
rect 5445 5148 5457 5151
rect 5224 5120 5457 5148
rect 5224 5108 5230 5120
rect 5445 5117 5457 5120
rect 5491 5117 5503 5151
rect 5445 5111 5503 5117
rect 6638 5108 6644 5160
rect 6696 5148 6702 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6696 5120 6837 5148
rect 6696 5108 6702 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 7009 5151 7067 5157
rect 7009 5117 7021 5151
rect 7055 5148 7067 5151
rect 7374 5148 7380 5160
rect 7055 5120 7380 5148
rect 7055 5117 7067 5120
rect 7009 5111 7067 5117
rect 7374 5108 7380 5120
rect 7432 5108 7438 5160
rect 9766 5108 9772 5160
rect 9824 5148 9830 5160
rect 10137 5151 10195 5157
rect 10137 5148 10149 5151
rect 9824 5120 10149 5148
rect 9824 5108 9830 5120
rect 10137 5117 10149 5120
rect 10183 5117 10195 5151
rect 10137 5111 10195 5117
rect 10870 5108 10876 5160
rect 10928 5148 10934 5160
rect 11149 5151 11207 5157
rect 11149 5148 11161 5151
rect 10928 5120 11161 5148
rect 10928 5108 10934 5120
rect 11149 5117 11161 5120
rect 11195 5148 11207 5151
rect 11514 5148 11520 5160
rect 11195 5120 11520 5148
rect 11195 5117 11207 5120
rect 11149 5111 11207 5117
rect 11514 5108 11520 5120
rect 11572 5108 11578 5160
rect 12621 5151 12679 5157
rect 12621 5117 12633 5151
rect 12667 5148 12679 5151
rect 12710 5148 12716 5160
rect 12667 5120 12716 5148
rect 12667 5117 12679 5120
rect 12621 5111 12679 5117
rect 12710 5108 12716 5120
rect 12768 5108 12774 5160
rect 12802 5108 12808 5160
rect 12860 5148 12866 5160
rect 13357 5151 13415 5157
rect 13357 5148 13369 5151
rect 12860 5120 13369 5148
rect 12860 5108 12866 5120
rect 13357 5117 13369 5120
rect 13403 5117 13415 5151
rect 16390 5148 16396 5160
rect 16351 5120 16396 5148
rect 13357 5111 13415 5117
rect 16390 5108 16396 5120
rect 16448 5108 16454 5160
rect 16482 5108 16488 5160
rect 16540 5148 16546 5160
rect 17604 5157 17632 5188
rect 17773 5185 17785 5219
rect 17819 5185 17831 5219
rect 17773 5179 17831 5185
rect 17313 5151 17371 5157
rect 17313 5148 17325 5151
rect 16540 5120 17325 5148
rect 16540 5108 16546 5120
rect 17313 5117 17325 5120
rect 17359 5117 17371 5151
rect 17313 5111 17371 5117
rect 17589 5151 17647 5157
rect 17589 5117 17601 5151
rect 17635 5117 17647 5151
rect 17589 5111 17647 5117
rect 10686 5040 10692 5092
rect 10744 5080 10750 5092
rect 12437 5083 12495 5089
rect 12437 5080 12449 5083
rect 10744 5052 12449 5080
rect 10744 5040 10750 5052
rect 12437 5049 12449 5052
rect 12483 5049 12495 5083
rect 12437 5043 12495 5049
rect 15381 5083 15439 5089
rect 15381 5049 15393 5083
rect 15427 5080 15439 5083
rect 16022 5080 16028 5092
rect 15427 5052 16028 5080
rect 15427 5049 15439 5052
rect 15381 5043 15439 5049
rect 16022 5040 16028 5052
rect 16080 5040 16086 5092
rect 2406 4972 2412 5024
rect 2464 5012 2470 5024
rect 2639 5015 2697 5021
rect 2639 5012 2651 5015
rect 2464 4984 2651 5012
rect 2464 4972 2470 4984
rect 2639 4981 2651 4984
rect 2685 4981 2697 5015
rect 2639 4975 2697 4981
rect 3421 5015 3479 5021
rect 3421 4981 3433 5015
rect 3467 5012 3479 5015
rect 7926 5012 7932 5024
rect 3467 4984 7932 5012
rect 3467 4981 3479 4984
rect 3421 4975 3479 4981
rect 7926 4972 7932 4984
rect 7984 4972 7990 5024
rect 10502 5012 10508 5024
rect 10463 4984 10508 5012
rect 10502 4972 10508 4984
rect 10560 4972 10566 5024
rect 12618 4972 12624 5024
rect 12676 5012 12682 5024
rect 13173 5015 13231 5021
rect 13173 5012 13185 5015
rect 12676 4984 13185 5012
rect 12676 4972 12682 4984
rect 13173 4981 13185 4984
rect 13219 4981 13231 5015
rect 15470 5012 15476 5024
rect 15431 4984 15476 5012
rect 13173 4975 13231 4981
rect 15470 4972 15476 4984
rect 15528 4972 15534 5024
rect 16666 4972 16672 5024
rect 16724 5012 16730 5024
rect 17405 5015 17463 5021
rect 17405 5012 17417 5015
rect 16724 4984 17417 5012
rect 16724 4972 16730 4984
rect 17405 4981 17417 4984
rect 17451 4981 17463 5015
rect 17405 4975 17463 4981
rect 1104 4922 19044 4944
rect 1104 4870 6962 4922
rect 7014 4870 7026 4922
rect 7078 4870 7090 4922
rect 7142 4870 7154 4922
rect 7206 4870 12942 4922
rect 12994 4870 13006 4922
rect 13058 4870 13070 4922
rect 13122 4870 13134 4922
rect 13186 4870 19044 4922
rect 1104 4848 19044 4870
rect 1486 4808 1492 4820
rect 1447 4780 1492 4808
rect 1486 4768 1492 4780
rect 1544 4768 1550 4820
rect 5626 4808 5632 4820
rect 5587 4780 5632 4808
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 7926 4768 7932 4820
rect 7984 4808 7990 4820
rect 13265 4811 13323 4817
rect 7984 4780 13216 4808
rect 7984 4768 7990 4780
rect 10502 4740 10508 4752
rect 10463 4712 10508 4740
rect 10502 4700 10508 4712
rect 10560 4700 10566 4752
rect 13188 4740 13216 4780
rect 13265 4777 13277 4811
rect 13311 4808 13323 4811
rect 13630 4808 13636 4820
rect 13311 4780 13636 4808
rect 13311 4777 13323 4780
rect 13265 4771 13323 4777
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 16022 4808 16028 4820
rect 15983 4780 16028 4808
rect 16022 4768 16028 4780
rect 16080 4768 16086 4820
rect 18138 4808 18144 4820
rect 18099 4780 18144 4808
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 13538 4740 13544 4752
rect 13188 4712 13544 4740
rect 13538 4700 13544 4712
rect 13596 4700 13602 4752
rect 1581 4675 1639 4681
rect 1581 4641 1593 4675
rect 1627 4641 1639 4675
rect 2406 4672 2412 4684
rect 2367 4644 2412 4672
rect 1581 4635 1639 4641
rect 1596 4604 1624 4635
rect 2406 4632 2412 4644
rect 2464 4632 2470 4684
rect 5166 4632 5172 4684
rect 5224 4672 5230 4684
rect 5813 4675 5871 4681
rect 5813 4672 5825 4675
rect 5224 4644 5825 4672
rect 5224 4632 5230 4644
rect 5813 4641 5825 4644
rect 5859 4672 5871 4675
rect 6273 4675 6331 4681
rect 6273 4672 6285 4675
rect 5859 4644 6285 4672
rect 5859 4641 5871 4644
rect 5813 4635 5871 4641
rect 6273 4641 6285 4644
rect 6319 4641 6331 4675
rect 6273 4635 6331 4641
rect 6457 4675 6515 4681
rect 6457 4641 6469 4675
rect 6503 4641 6515 4675
rect 6457 4635 6515 4641
rect 4338 4604 4344 4616
rect 1596 4576 4344 4604
rect 4338 4564 4344 4576
rect 4396 4564 4402 4616
rect 2314 4468 2320 4480
rect 2275 4440 2320 4468
rect 2314 4428 2320 4440
rect 2372 4428 2378 4480
rect 6472 4468 6500 4635
rect 9766 4632 9772 4684
rect 9824 4672 9830 4684
rect 10045 4675 10103 4681
rect 10045 4672 10057 4675
rect 9824 4644 10057 4672
rect 9824 4632 9830 4644
rect 10045 4641 10057 4644
rect 10091 4641 10103 4675
rect 10045 4635 10103 4641
rect 10597 4675 10655 4681
rect 10597 4641 10609 4675
rect 10643 4672 10655 4675
rect 11514 4672 11520 4684
rect 10643 4644 11520 4672
rect 10643 4641 10655 4644
rect 10597 4635 10655 4641
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 11790 4632 11796 4684
rect 11848 4672 11854 4684
rect 12437 4675 12495 4681
rect 12437 4672 12449 4675
rect 11848 4644 12449 4672
rect 11848 4632 11854 4644
rect 12437 4641 12449 4644
rect 12483 4672 12495 4675
rect 12710 4672 12716 4684
rect 12483 4644 12716 4672
rect 12483 4641 12495 4644
rect 12437 4635 12495 4641
rect 12710 4632 12716 4644
rect 12768 4632 12774 4684
rect 16390 4672 16396 4684
rect 16351 4644 16396 4672
rect 16390 4632 16396 4644
rect 16448 4632 16454 4684
rect 18322 4672 18328 4684
rect 18283 4644 18328 4672
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 7282 4604 7288 4616
rect 7243 4576 7288 4604
rect 7282 4564 7288 4576
rect 7340 4564 7346 4616
rect 7650 4604 7656 4616
rect 7611 4576 7656 4604
rect 7650 4564 7656 4576
rect 7708 4564 7714 4616
rect 11606 4604 11612 4616
rect 11567 4576 11612 4604
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 12894 4604 12900 4616
rect 12855 4576 12900 4604
rect 12894 4564 12900 4576
rect 12952 4564 12958 4616
rect 16485 4607 16543 4613
rect 16485 4573 16497 4607
rect 16531 4573 16543 4607
rect 16666 4604 16672 4616
rect 16627 4576 16672 4604
rect 16485 4567 16543 4573
rect 13262 4536 13268 4548
rect 13223 4508 13268 4536
rect 13262 4496 13268 4508
rect 13320 4496 13326 4548
rect 16500 4536 16528 4567
rect 16666 4564 16672 4576
rect 16724 4564 16730 4616
rect 16574 4536 16580 4548
rect 16500 4508 16580 4536
rect 16574 4496 16580 4508
rect 16632 4536 16638 4548
rect 18414 4536 18420 4548
rect 16632 4508 18420 4536
rect 16632 4496 16638 4508
rect 18414 4496 18420 4508
rect 18472 4496 18478 4548
rect 7285 4471 7343 4477
rect 7285 4468 7297 4471
rect 6472 4440 7297 4468
rect 7285 4437 7297 4440
rect 7331 4468 7343 4471
rect 7374 4468 7380 4480
rect 7331 4440 7380 4468
rect 7331 4437 7343 4440
rect 7285 4431 7343 4437
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 1104 4378 19044 4400
rect 1104 4326 3972 4378
rect 4024 4326 4036 4378
rect 4088 4326 4100 4378
rect 4152 4326 4164 4378
rect 4216 4326 9952 4378
rect 10004 4326 10016 4378
rect 10068 4326 10080 4378
rect 10132 4326 10144 4378
rect 10196 4326 15932 4378
rect 15984 4326 15996 4378
rect 16048 4326 16060 4378
rect 16112 4326 16124 4378
rect 16176 4326 19044 4378
rect 1104 4304 19044 4326
rect 7650 4264 7656 4276
rect 7611 4236 7656 4264
rect 7650 4224 7656 4236
rect 7708 4224 7714 4276
rect 9766 4224 9772 4276
rect 9824 4264 9830 4276
rect 9861 4267 9919 4273
rect 9861 4264 9873 4267
rect 9824 4236 9873 4264
rect 9824 4224 9830 4236
rect 9861 4233 9873 4236
rect 9907 4233 9919 4267
rect 9861 4227 9919 4233
rect 12805 4267 12863 4273
rect 12805 4233 12817 4267
rect 12851 4264 12863 4267
rect 12894 4264 12900 4276
rect 12851 4236 12900 4264
rect 12851 4233 12863 4236
rect 12805 4227 12863 4233
rect 12894 4224 12900 4236
rect 12952 4224 12958 4276
rect 7558 4196 7564 4208
rect 7116 4168 7564 4196
rect 7116 4137 7144 4168
rect 7558 4156 7564 4168
rect 7616 4196 7622 4208
rect 9582 4196 9588 4208
rect 7616 4168 9588 4196
rect 7616 4156 7622 4168
rect 9582 4156 9588 4168
rect 9640 4196 9646 4208
rect 11606 4196 11612 4208
rect 9640 4168 11612 4196
rect 9640 4156 9646 4168
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4097 7159 4131
rect 7101 4091 7159 4097
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 8481 4131 8539 4137
rect 8481 4128 8493 4131
rect 7432 4100 8493 4128
rect 7432 4088 7438 4100
rect 8481 4097 8493 4100
rect 8527 4097 8539 4131
rect 10318 4128 10324 4140
rect 8481 4091 8539 4097
rect 9232 4100 10324 4128
rect 7285 4063 7343 4069
rect 7285 4029 7297 4063
rect 7331 4060 7343 4063
rect 7466 4060 7472 4072
rect 7331 4032 7472 4060
rect 7331 4029 7343 4032
rect 7285 4023 7343 4029
rect 7466 4020 7472 4032
rect 7524 4020 7530 4072
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 8113 4063 8171 4069
rect 8113 4060 8125 4063
rect 7708 4032 8125 4060
rect 7708 4020 7714 4032
rect 8113 4029 8125 4032
rect 8159 4029 8171 4063
rect 8662 4060 8668 4072
rect 8623 4032 8668 4060
rect 8113 4023 8171 4029
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 9232 4069 9260 4100
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 10520 4137 10548 4168
rect 11606 4156 11612 4168
rect 11664 4156 11670 4208
rect 12710 4196 12716 4208
rect 12268 4168 12716 4196
rect 12268 4137 12296 4168
rect 12710 4156 12716 4168
rect 12768 4156 12774 4208
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4097 12311 4131
rect 12253 4091 12311 4097
rect 12345 4131 12403 4137
rect 12345 4097 12357 4131
rect 12391 4128 12403 4131
rect 12618 4128 12624 4140
rect 12391 4100 12624 4128
rect 12391 4097 12403 4100
rect 12345 4091 12403 4097
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 13630 4128 13636 4140
rect 13591 4100 13636 4128
rect 13630 4088 13636 4100
rect 13688 4128 13694 4140
rect 13688 4100 15056 4128
rect 13688 4088 13694 4100
rect 9217 4063 9275 4069
rect 9217 4029 9229 4063
rect 9263 4029 9275 4063
rect 12434 4060 12440 4072
rect 9217 4023 9275 4029
rect 9324 4032 10456 4060
rect 12395 4032 12440 4060
rect 7193 3995 7251 4001
rect 7193 3961 7205 3995
rect 7239 3992 7251 3995
rect 9324 3992 9352 4032
rect 10321 3995 10379 4001
rect 10321 3992 10333 3995
rect 7239 3964 9352 3992
rect 9416 3964 10333 3992
rect 7239 3961 7251 3964
rect 7193 3955 7251 3961
rect 9416 3933 9444 3964
rect 10321 3961 10333 3964
rect 10367 3961 10379 3995
rect 10428 3992 10456 4032
rect 12434 4020 12440 4032
rect 12492 4020 12498 4072
rect 12894 4020 12900 4072
rect 12952 4060 12958 4072
rect 13265 4063 13323 4069
rect 13265 4060 13277 4063
rect 12952 4032 13277 4060
rect 12952 4020 12958 4032
rect 13265 4029 13277 4032
rect 13311 4029 13323 4063
rect 13265 4023 13323 4029
rect 13538 4020 13544 4072
rect 13596 4060 13602 4072
rect 15028 4069 15056 4100
rect 13817 4063 13875 4069
rect 13817 4060 13829 4063
rect 13596 4032 13829 4060
rect 13596 4020 13602 4032
rect 13817 4029 13829 4032
rect 13863 4029 13875 4063
rect 13817 4023 13875 4029
rect 15013 4063 15071 4069
rect 15013 4029 15025 4063
rect 15059 4029 15071 4063
rect 15013 4023 15071 4029
rect 13354 3992 13360 4004
rect 10428 3964 13360 3992
rect 10321 3955 10379 3961
rect 13354 3952 13360 3964
rect 13412 3952 13418 4004
rect 13446 3952 13452 4004
rect 13504 3992 13510 4004
rect 14277 3995 14335 4001
rect 14277 3992 14289 3995
rect 13504 3964 14289 3992
rect 13504 3952 13510 3964
rect 14277 3961 14289 3964
rect 14323 3961 14335 3995
rect 14277 3955 14335 3961
rect 14461 3995 14519 4001
rect 14461 3961 14473 3995
rect 14507 3992 14519 3995
rect 14507 3964 15056 3992
rect 14507 3961 14519 3964
rect 14461 3955 14519 3961
rect 15028 3936 15056 3964
rect 9401 3927 9459 3933
rect 9401 3893 9413 3927
rect 9447 3893 9459 3927
rect 9401 3887 9459 3893
rect 10229 3927 10287 3933
rect 10229 3893 10241 3927
rect 10275 3924 10287 3927
rect 10778 3924 10784 3936
rect 10275 3896 10784 3924
rect 10275 3893 10287 3896
rect 10229 3887 10287 3893
rect 10778 3884 10784 3896
rect 10836 3884 10842 3936
rect 15010 3884 15016 3936
rect 15068 3884 15074 3936
rect 15102 3884 15108 3936
rect 15160 3924 15166 3936
rect 15160 3896 15205 3924
rect 15160 3884 15166 3896
rect 1104 3834 19044 3856
rect 1104 3782 6962 3834
rect 7014 3782 7026 3834
rect 7078 3782 7090 3834
rect 7142 3782 7154 3834
rect 7206 3782 12942 3834
rect 12994 3782 13006 3834
rect 13058 3782 13070 3834
rect 13122 3782 13134 3834
rect 13186 3782 19044 3834
rect 1104 3760 19044 3782
rect 6822 3720 6828 3732
rect 5644 3692 6828 3720
rect 5644 3638 5672 3692
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7469 3723 7527 3729
rect 7469 3689 7481 3723
rect 7515 3720 7527 3723
rect 8297 3723 8355 3729
rect 8297 3720 8309 3723
rect 7515 3692 8309 3720
rect 7515 3689 7527 3692
rect 7469 3683 7527 3689
rect 8297 3689 8309 3692
rect 8343 3720 8355 3723
rect 8386 3720 8392 3732
rect 8343 3692 8392 3720
rect 8343 3689 8355 3692
rect 8297 3683 8355 3689
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 10965 3723 11023 3729
rect 10965 3689 10977 3723
rect 11011 3689 11023 3723
rect 11514 3720 11520 3732
rect 11475 3692 11520 3720
rect 10965 3683 11023 3689
rect 5810 3612 5816 3664
rect 5868 3652 5874 3664
rect 7282 3652 7288 3664
rect 5868 3624 6408 3652
rect 7243 3624 7288 3652
rect 5868 3612 5874 3624
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 4338 3584 4344 3596
rect 4251 3556 4344 3584
rect 4338 3544 4344 3556
rect 4396 3544 4402 3596
rect 6380 3593 6408 3624
rect 7282 3612 7288 3624
rect 7340 3612 7346 3664
rect 10502 3612 10508 3664
rect 10560 3652 10566 3664
rect 10980 3652 11008 3683
rect 11514 3680 11520 3692
rect 11572 3680 11578 3732
rect 13262 3720 13268 3732
rect 13223 3692 13268 3720
rect 13262 3680 13268 3692
rect 13320 3680 13326 3732
rect 13354 3680 13360 3732
rect 13412 3720 13418 3732
rect 18138 3720 18144 3732
rect 13412 3692 18144 3720
rect 13412 3680 13418 3692
rect 18138 3680 18144 3692
rect 18196 3680 18202 3732
rect 11609 3655 11667 3661
rect 11609 3652 11621 3655
rect 10560 3624 11621 3652
rect 10560 3612 10566 3624
rect 11609 3621 11621 3624
rect 11655 3621 11667 3655
rect 11609 3615 11667 3621
rect 12526 3612 12532 3664
rect 12584 3612 12590 3664
rect 15562 3612 15568 3664
rect 15620 3652 15626 3664
rect 15620 3624 16330 3652
rect 15620 3612 15626 3624
rect 6365 3587 6423 3593
rect 6365 3553 6377 3587
rect 6411 3553 6423 3587
rect 6365 3547 6423 3553
rect 8662 3544 8668 3596
rect 8720 3584 8726 3596
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 8720 3556 9689 3584
rect 8720 3544 8726 3556
rect 9677 3553 9689 3556
rect 9723 3584 9735 3587
rect 10686 3584 10692 3596
rect 9723 3556 10692 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 12544 3584 12572 3612
rect 12621 3587 12679 3593
rect 12621 3584 12633 3587
rect 12544 3556 12633 3584
rect 12621 3553 12633 3556
rect 12667 3553 12679 3587
rect 12621 3547 12679 3553
rect 13449 3587 13507 3593
rect 13449 3553 13461 3587
rect 13495 3584 13507 3587
rect 13538 3584 13544 3596
rect 13495 3556 13544 3584
rect 13495 3553 13507 3556
rect 13449 3547 13507 3553
rect 13538 3544 13544 3556
rect 13596 3544 13602 3596
rect 15102 3584 15108 3596
rect 15063 3556 15108 3584
rect 15102 3544 15108 3556
rect 15160 3544 15166 3596
rect 17589 3587 17647 3593
rect 17589 3553 17601 3587
rect 17635 3553 17647 3587
rect 18322 3584 18328 3596
rect 18283 3556 18328 3584
rect 17589 3547 17647 3553
rect 4356 3516 4384 3544
rect 6089 3519 6147 3525
rect 6089 3516 6101 3519
rect 4356 3488 6101 3516
rect 6089 3485 6101 3488
rect 6135 3516 6147 3519
rect 7926 3516 7932 3528
rect 6135 3488 6316 3516
rect 7887 3488 7932 3516
rect 6135 3485 6147 3488
rect 6089 3479 6147 3485
rect 6288 3448 6316 3488
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 10318 3476 10324 3528
rect 10376 3516 10382 3528
rect 10597 3519 10655 3525
rect 10597 3516 10609 3519
rect 10376 3488 10609 3516
rect 10376 3476 10382 3488
rect 10597 3485 10609 3488
rect 10643 3485 10655 3519
rect 10597 3479 10655 3485
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3516 12311 3519
rect 12526 3516 12532 3528
rect 12299 3488 12532 3516
rect 12299 3485 12311 3488
rect 12253 3479 12311 3485
rect 12526 3476 12532 3488
rect 12584 3476 12590 3528
rect 14734 3516 14740 3528
rect 14695 3488 14740 3516
rect 14734 3476 14740 3488
rect 14792 3476 14798 3528
rect 15565 3519 15623 3525
rect 15565 3485 15577 3519
rect 15611 3485 15623 3519
rect 15565 3479 15623 3485
rect 15841 3519 15899 3525
rect 15841 3485 15853 3519
rect 15887 3516 15899 3519
rect 16574 3516 16580 3528
rect 15887 3488 16580 3516
rect 15887 3485 15899 3488
rect 15841 3479 15899 3485
rect 8297 3451 8355 3457
rect 6288 3420 8248 3448
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3380 1639 3383
rect 8110 3380 8116 3392
rect 1627 3352 8116 3380
rect 1627 3349 1639 3352
rect 1581 3343 1639 3349
rect 8110 3340 8116 3352
rect 8168 3340 8174 3392
rect 8220 3380 8248 3420
rect 8297 3417 8309 3451
rect 8343 3448 8355 3451
rect 9493 3451 9551 3457
rect 9493 3448 9505 3451
rect 8343 3420 9505 3448
rect 8343 3417 8355 3420
rect 8297 3411 8355 3417
rect 9493 3417 9505 3420
rect 9539 3417 9551 3451
rect 9493 3411 9551 3417
rect 10965 3451 11023 3457
rect 10965 3417 10977 3451
rect 11011 3448 11023 3451
rect 11054 3448 11060 3460
rect 11011 3420 11060 3448
rect 11011 3417 11023 3420
rect 10965 3411 11023 3417
rect 11054 3408 11060 3420
rect 11112 3408 11118 3460
rect 15470 3448 15476 3460
rect 11164 3420 15476 3448
rect 11164 3380 11192 3420
rect 15470 3408 15476 3420
rect 15528 3448 15534 3460
rect 15580 3448 15608 3479
rect 16574 3476 16580 3488
rect 16632 3516 16638 3528
rect 17604 3516 17632 3547
rect 18322 3544 18328 3556
rect 18380 3544 18386 3596
rect 16632 3488 17632 3516
rect 16632 3476 16638 3488
rect 15528 3420 15608 3448
rect 15528 3408 15534 3420
rect 8220 3352 11192 3380
rect 12066 3340 12072 3392
rect 12124 3380 12130 3392
rect 12253 3383 12311 3389
rect 12253 3380 12265 3383
rect 12124 3352 12265 3380
rect 12124 3340 12130 3352
rect 12253 3349 12265 3352
rect 12299 3349 12311 3383
rect 15102 3380 15108 3392
rect 15063 3352 15108 3380
rect 12253 3343 12311 3349
rect 15102 3340 15108 3352
rect 15160 3340 15166 3392
rect 17310 3340 17316 3392
rect 17368 3380 17374 3392
rect 18141 3383 18199 3389
rect 18141 3380 18153 3383
rect 17368 3352 18153 3380
rect 17368 3340 17374 3352
rect 18141 3349 18153 3352
rect 18187 3349 18199 3383
rect 18141 3343 18199 3349
rect 1104 3290 19044 3312
rect 1104 3238 3972 3290
rect 4024 3238 4036 3290
rect 4088 3238 4100 3290
rect 4152 3238 4164 3290
rect 4216 3238 9952 3290
rect 10004 3238 10016 3290
rect 10068 3238 10080 3290
rect 10132 3238 10144 3290
rect 10196 3238 15932 3290
rect 15984 3238 15996 3290
rect 16048 3238 16060 3290
rect 16112 3238 16124 3290
rect 16176 3238 19044 3290
rect 1104 3216 19044 3238
rect 8386 3176 8392 3188
rect 8347 3148 8392 3176
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 10502 3176 10508 3188
rect 10463 3148 10508 3176
rect 10502 3136 10508 3148
rect 10560 3136 10566 3188
rect 11054 3176 11060 3188
rect 11015 3148 11060 3176
rect 11054 3136 11060 3148
rect 11112 3136 11118 3188
rect 12066 3176 12072 3188
rect 12027 3148 12072 3176
rect 12066 3136 12072 3148
rect 12124 3136 12130 3188
rect 13357 3179 13415 3185
rect 13357 3145 13369 3179
rect 13403 3176 13415 3179
rect 15102 3176 15108 3188
rect 13403 3148 15108 3176
rect 13403 3145 13415 3148
rect 13357 3139 13415 3145
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 16942 3136 16948 3188
rect 17000 3176 17006 3188
rect 17313 3179 17371 3185
rect 17313 3176 17325 3179
rect 17000 3148 17325 3176
rect 17000 3136 17006 3148
rect 17313 3145 17325 3148
rect 17359 3145 17371 3179
rect 18138 3176 18144 3188
rect 18099 3148 18144 3176
rect 17313 3139 17371 3145
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 5718 3108 5724 3120
rect 4356 3080 5724 3108
rect 2314 3000 2320 3052
rect 2372 3040 2378 3052
rect 3053 3043 3111 3049
rect 3053 3040 3065 3043
rect 2372 3012 3065 3040
rect 2372 3000 2378 3012
rect 3053 3009 3065 3012
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3040 3387 3043
rect 4356 3040 4384 3080
rect 5718 3068 5724 3080
rect 5776 3068 5782 3120
rect 8662 3108 8668 3120
rect 8404 3080 8668 3108
rect 6822 3040 6828 3052
rect 3375 3012 4384 3040
rect 4448 3012 6828 3040
rect 3375 3009 3387 3012
rect 3329 3003 3387 3009
rect 474 2932 480 2984
rect 532 2972 538 2984
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 532 2944 1409 2972
rect 532 2932 538 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 4448 2958 4476 3012
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 5077 2975 5135 2981
rect 1397 2935 1455 2941
rect 5077 2941 5089 2975
rect 5123 2972 5135 2975
rect 5718 2972 5724 2984
rect 5123 2944 5724 2972
rect 5123 2941 5135 2944
rect 5077 2935 5135 2941
rect 5718 2932 5724 2944
rect 5776 2932 5782 2984
rect 5902 2932 5908 2984
rect 5960 2972 5966 2984
rect 6917 2975 6975 2981
rect 6917 2972 6929 2975
rect 5960 2944 6929 2972
rect 5960 2932 5966 2944
rect 6917 2941 6929 2944
rect 6963 2941 6975 2975
rect 6917 2935 6975 2941
rect 7837 2975 7895 2981
rect 7837 2941 7849 2975
rect 7883 2972 7895 2975
rect 7926 2972 7932 2984
rect 7883 2944 7932 2972
rect 7883 2941 7895 2944
rect 7837 2935 7895 2941
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 8404 2981 8432 3080
rect 8662 3068 8668 3080
rect 8720 3068 8726 3120
rect 9490 3108 9496 3120
rect 9451 3080 9496 3108
rect 9490 3068 9496 3080
rect 9548 3068 9554 3120
rect 16574 3108 16580 3120
rect 16408 3080 16580 3108
rect 15562 3040 15568 3052
rect 9876 3012 15568 3040
rect 8389 2975 8447 2981
rect 8389 2941 8401 2975
rect 8435 2941 8447 2975
rect 9766 2972 9772 2984
rect 8389 2935 8447 2941
rect 8496 2944 9772 2972
rect 8496 2904 8524 2944
rect 9766 2932 9772 2944
rect 9824 2932 9830 2984
rect 6288 2876 8524 2904
rect 1581 2839 1639 2845
rect 1581 2805 1593 2839
rect 1627 2836 1639 2839
rect 6288 2836 6316 2876
rect 9214 2864 9220 2916
rect 9272 2904 9278 2916
rect 9309 2907 9367 2913
rect 9309 2904 9321 2907
rect 9272 2876 9321 2904
rect 9272 2864 9278 2876
rect 9309 2873 9321 2876
rect 9355 2873 9367 2907
rect 9309 2867 9367 2873
rect 1627 2808 6316 2836
rect 1627 2805 1639 2808
rect 1581 2799 1639 2805
rect 6822 2796 6828 2848
rect 6880 2836 6886 2848
rect 7101 2839 7159 2845
rect 7101 2836 7113 2839
rect 6880 2808 7113 2836
rect 6880 2796 6886 2808
rect 7101 2805 7113 2808
rect 7147 2836 7159 2839
rect 9876 2836 9904 3012
rect 15562 3000 15568 3012
rect 15620 3000 15626 3052
rect 16408 3049 16436 3080
rect 16574 3068 16580 3080
rect 16632 3068 16638 3120
rect 16393 3043 16451 3049
rect 16393 3009 16405 3043
rect 16439 3009 16451 3043
rect 16393 3003 16451 3009
rect 9953 2975 10011 2981
rect 9953 2941 9965 2975
rect 9999 2972 10011 2975
rect 10318 2972 10324 2984
rect 9999 2944 10324 2972
rect 9999 2941 10011 2944
rect 9953 2935 10011 2941
rect 10318 2932 10324 2944
rect 10376 2932 10382 2984
rect 10505 2975 10563 2981
rect 10505 2941 10517 2975
rect 10551 2972 10563 2975
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 10551 2944 12081 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 12069 2941 12081 2944
rect 12115 2972 12127 2975
rect 12434 2972 12440 2984
rect 12115 2944 12440 2972
rect 12115 2941 12127 2944
rect 12069 2935 12127 2941
rect 12434 2932 12440 2944
rect 12492 2932 12498 2984
rect 12618 2972 12624 2984
rect 12579 2944 12624 2972
rect 12618 2932 12624 2944
rect 12676 2932 12682 2984
rect 13357 2975 13415 2981
rect 13357 2941 13369 2975
rect 13403 2972 13415 2975
rect 13538 2972 13544 2984
rect 13403 2944 13544 2972
rect 13403 2941 13415 2944
rect 13357 2935 13415 2941
rect 13538 2932 13544 2944
rect 13596 2932 13602 2984
rect 13909 2975 13967 2981
rect 13909 2941 13921 2975
rect 13955 2972 13967 2975
rect 14734 2972 14740 2984
rect 13955 2944 14740 2972
rect 13955 2941 13967 2944
rect 13909 2935 13967 2941
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 16574 2932 16580 2984
rect 16632 2972 16638 2984
rect 17497 2975 17555 2981
rect 17497 2972 17509 2975
rect 16632 2944 17509 2972
rect 16632 2932 16638 2944
rect 17497 2941 17509 2944
rect 17543 2941 17555 2975
rect 17497 2935 17555 2941
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2972 18383 2975
rect 18414 2972 18420 2984
rect 18371 2944 18420 2972
rect 18371 2941 18383 2944
rect 18325 2935 18383 2941
rect 18414 2932 18420 2944
rect 18472 2932 18478 2984
rect 11149 2907 11207 2913
rect 11149 2873 11161 2907
rect 11195 2904 11207 2907
rect 12158 2904 12164 2916
rect 11195 2876 12164 2904
rect 11195 2873 11207 2876
rect 11149 2867 11207 2873
rect 12158 2864 12164 2876
rect 12216 2864 12222 2916
rect 15562 2864 15568 2916
rect 15620 2864 15626 2916
rect 16117 2907 16175 2913
rect 16117 2873 16129 2907
rect 16163 2904 16175 2907
rect 16390 2904 16396 2916
rect 16163 2876 16396 2904
rect 16163 2873 16175 2876
rect 16117 2867 16175 2873
rect 7147 2808 9904 2836
rect 7147 2805 7159 2808
rect 7101 2799 7159 2805
rect 11974 2796 11980 2848
rect 12032 2836 12038 2848
rect 12802 2836 12808 2848
rect 12032 2808 12808 2836
rect 12032 2796 12038 2808
rect 12802 2796 12808 2808
rect 12860 2796 12866 2848
rect 14369 2839 14427 2845
rect 14369 2805 14381 2839
rect 14415 2836 14427 2839
rect 16132 2836 16160 2867
rect 16390 2864 16396 2876
rect 16448 2864 16454 2916
rect 14415 2808 16160 2836
rect 14415 2805 14427 2808
rect 14369 2799 14427 2805
rect 1104 2746 19044 2768
rect 1104 2694 6962 2746
rect 7014 2694 7026 2746
rect 7078 2694 7090 2746
rect 7142 2694 7154 2746
rect 7206 2694 12942 2746
rect 12994 2694 13006 2746
rect 13058 2694 13070 2746
rect 13122 2694 13134 2746
rect 13186 2694 19044 2746
rect 1104 2672 19044 2694
rect 3329 2635 3387 2641
rect 3329 2601 3341 2635
rect 3375 2632 3387 2635
rect 3510 2632 3516 2644
rect 3375 2604 3516 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 4801 2635 4859 2641
rect 4801 2601 4813 2635
rect 4847 2632 4859 2635
rect 4890 2632 4896 2644
rect 4847 2604 4896 2632
rect 4847 2601 4859 2604
rect 4801 2595 4859 2601
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 5813 2635 5871 2641
rect 5813 2601 5825 2635
rect 5859 2632 5871 2635
rect 5902 2632 5908 2644
rect 5859 2604 5908 2632
rect 5859 2601 5871 2604
rect 5813 2595 5871 2601
rect 5902 2592 5908 2604
rect 5960 2592 5966 2644
rect 7653 2635 7711 2641
rect 7653 2601 7665 2635
rect 7699 2632 7711 2635
rect 7834 2632 7840 2644
rect 7699 2604 7840 2632
rect 7699 2601 7711 2604
rect 7653 2595 7711 2601
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8110 2632 8116 2644
rect 8071 2604 8116 2632
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 9953 2635 10011 2641
rect 9953 2632 9965 2635
rect 9732 2604 9965 2632
rect 9732 2592 9738 2604
rect 9953 2601 9965 2604
rect 9999 2601 10011 2635
rect 10318 2632 10324 2644
rect 10279 2604 10324 2632
rect 9953 2595 10011 2601
rect 10318 2592 10324 2604
rect 10376 2592 10382 2644
rect 10870 2632 10876 2644
rect 10831 2604 10876 2632
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 12526 2592 12532 2644
rect 12584 2632 12590 2644
rect 12621 2635 12679 2641
rect 12621 2632 12633 2635
rect 12584 2604 12633 2632
rect 12584 2592 12590 2604
rect 12621 2601 12633 2604
rect 12667 2601 12679 2635
rect 12621 2595 12679 2601
rect 14734 2592 14740 2644
rect 14792 2632 14798 2644
rect 14921 2635 14979 2641
rect 14921 2632 14933 2635
rect 14792 2604 14933 2632
rect 14792 2592 14798 2604
rect 14921 2601 14933 2604
rect 14967 2601 14979 2635
rect 14921 2595 14979 2601
rect 15381 2635 15439 2641
rect 15381 2601 15393 2635
rect 15427 2632 15439 2635
rect 17310 2632 17316 2644
rect 15427 2604 17316 2632
rect 15427 2601 15439 2604
rect 15381 2595 15439 2601
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 2041 2567 2099 2573
rect 2041 2533 2053 2567
rect 2087 2564 2099 2567
rect 2314 2564 2320 2576
rect 2087 2536 2320 2564
rect 2087 2533 2099 2536
rect 2041 2527 2099 2533
rect 2314 2524 2320 2536
rect 2372 2524 2378 2576
rect 6546 2524 6552 2576
rect 6604 2564 6610 2576
rect 6604 2536 14044 2564
rect 6604 2524 6610 2536
rect 3145 2499 3203 2505
rect 3145 2465 3157 2499
rect 3191 2496 3203 2499
rect 3234 2496 3240 2508
rect 3191 2468 3240 2496
rect 3191 2465 3203 2468
rect 3145 2459 3203 2465
rect 3234 2456 3240 2468
rect 3292 2456 3298 2508
rect 4614 2496 4620 2508
rect 4575 2468 4620 2496
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 5994 2496 6000 2508
rect 5955 2468 6000 2496
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2496 7067 2499
rect 7834 2496 7840 2508
rect 7055 2468 7840 2496
rect 7055 2465 7067 2468
rect 7009 2459 7067 2465
rect 7834 2456 7840 2468
rect 7892 2456 7898 2508
rect 8018 2496 8024 2508
rect 7979 2468 8024 2496
rect 8018 2456 8024 2468
rect 8076 2456 8082 2508
rect 9766 2456 9772 2508
rect 9824 2496 9830 2508
rect 10781 2499 10839 2505
rect 10781 2496 10793 2499
rect 9824 2468 10793 2496
rect 9824 2456 9830 2468
rect 10781 2465 10793 2468
rect 10827 2465 10839 2499
rect 10781 2459 10839 2465
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 12805 2499 12863 2505
rect 12805 2496 12817 2499
rect 12492 2468 12817 2496
rect 12492 2456 12498 2468
rect 12805 2465 12817 2468
rect 12851 2496 12863 2499
rect 13446 2496 13452 2508
rect 12851 2468 13452 2496
rect 12851 2465 12863 2468
rect 12805 2459 12863 2465
rect 13446 2456 13452 2468
rect 13504 2456 13510 2508
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 13909 2499 13967 2505
rect 13909 2496 13921 2499
rect 13872 2468 13921 2496
rect 13872 2456 13878 2468
rect 13909 2465 13921 2468
rect 13955 2465 13967 2499
rect 14016 2496 14044 2536
rect 15194 2524 15200 2576
rect 15252 2564 15258 2576
rect 16209 2567 16267 2573
rect 16209 2564 16221 2567
rect 15252 2536 16221 2564
rect 15252 2524 15258 2536
rect 16209 2533 16221 2536
rect 16255 2533 16267 2567
rect 16209 2527 16267 2533
rect 16390 2524 16396 2576
rect 16448 2564 16454 2576
rect 18141 2567 18199 2573
rect 18141 2564 18153 2567
rect 16448 2536 18153 2564
rect 16448 2524 16454 2536
rect 18141 2533 18153 2536
rect 18187 2533 18199 2567
rect 18141 2527 18199 2533
rect 15289 2499 15347 2505
rect 15289 2496 15301 2499
rect 14016 2468 15301 2496
rect 13909 2459 13967 2465
rect 15289 2465 15301 2468
rect 15335 2465 15347 2499
rect 15289 2459 15347 2465
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2428 8355 2431
rect 9582 2428 9588 2440
rect 8343 2400 9588 2428
rect 8343 2397 8355 2400
rect 8297 2391 8355 2397
rect 9582 2388 9588 2400
rect 9640 2428 9646 2440
rect 9677 2431 9735 2437
rect 9677 2428 9689 2431
rect 9640 2400 9689 2428
rect 9640 2388 9646 2400
rect 9677 2397 9689 2400
rect 9723 2397 9735 2431
rect 9677 2391 9735 2397
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 1854 2360 1860 2372
rect 1815 2332 1860 2360
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 7193 2363 7251 2369
rect 7193 2329 7205 2363
rect 7239 2360 7251 2363
rect 9876 2360 9904 2391
rect 12710 2388 12716 2440
rect 12768 2428 12774 2440
rect 13633 2431 13691 2437
rect 13633 2428 13645 2431
rect 12768 2400 13645 2428
rect 12768 2388 12774 2400
rect 13633 2397 13645 2400
rect 13679 2428 13691 2431
rect 15473 2431 15531 2437
rect 15473 2428 15485 2431
rect 13679 2400 15485 2428
rect 13679 2397 13691 2400
rect 13633 2391 13691 2397
rect 15473 2397 15485 2400
rect 15519 2397 15531 2431
rect 15473 2391 15531 2397
rect 16393 2431 16451 2437
rect 16393 2397 16405 2431
rect 16439 2428 16451 2431
rect 16482 2428 16488 2440
rect 16439 2400 16488 2428
rect 16439 2397 16451 2400
rect 16393 2391 16451 2397
rect 16482 2388 16488 2400
rect 16540 2388 16546 2440
rect 17954 2360 17960 2372
rect 7239 2332 9904 2360
rect 17915 2332 17960 2360
rect 7239 2329 7251 2332
rect 7193 2323 7251 2329
rect 17954 2320 17960 2332
rect 18012 2320 18018 2372
rect 1104 2202 19044 2224
rect 1104 2150 3972 2202
rect 4024 2150 4036 2202
rect 4088 2150 4100 2202
rect 4152 2150 4164 2202
rect 4216 2150 9952 2202
rect 10004 2150 10016 2202
rect 10068 2150 10080 2202
rect 10132 2150 10144 2202
rect 10196 2150 15932 2202
rect 15984 2150 15996 2202
rect 16048 2150 16060 2202
rect 16112 2150 16124 2202
rect 16176 2150 19044 2202
rect 1104 2128 19044 2150
<< via1 >>
rect 6962 20102 7014 20154
rect 7026 20102 7078 20154
rect 7090 20102 7142 20154
rect 7154 20102 7206 20154
rect 12942 20102 12994 20154
rect 13006 20102 13058 20154
rect 13070 20102 13122 20154
rect 13134 20102 13186 20154
rect 1492 20043 1544 20052
rect 1492 20009 1501 20043
rect 1501 20009 1535 20043
rect 1535 20009 1544 20043
rect 1492 20000 1544 20009
rect 7104 19932 7156 19984
rect 8300 19932 8352 19984
rect 1584 19907 1636 19916
rect 1584 19873 1593 19907
rect 1593 19873 1627 19907
rect 1627 19873 1636 19907
rect 1584 19864 1636 19873
rect 2320 19907 2372 19916
rect 2320 19873 2329 19907
rect 2329 19873 2363 19907
rect 2363 19873 2372 19907
rect 2320 19864 2372 19873
rect 2964 19864 3016 19916
rect 3700 19864 3752 19916
rect 5540 19907 5592 19916
rect 5540 19873 5549 19907
rect 5549 19873 5583 19907
rect 5583 19873 5592 19907
rect 5540 19864 5592 19873
rect 6920 19907 6972 19916
rect 6920 19873 6929 19907
rect 6929 19873 6963 19907
rect 6963 19873 6972 19907
rect 6920 19864 6972 19873
rect 7380 19864 7432 19916
rect 7840 19907 7892 19916
rect 7840 19873 7849 19907
rect 7849 19873 7883 19907
rect 7883 19873 7892 19907
rect 7840 19864 7892 19873
rect 8208 19864 8260 19916
rect 9680 19864 9732 19916
rect 18880 19932 18932 19984
rect 11520 19864 11572 19916
rect 12808 19864 12860 19916
rect 14280 19864 14332 19916
rect 15660 19864 15712 19916
rect 16488 19864 16540 19916
rect 8576 19728 8628 19780
rect 10692 19728 10744 19780
rect 18052 19771 18104 19780
rect 18052 19737 18061 19771
rect 18061 19737 18095 19771
rect 18095 19737 18104 19771
rect 18052 19728 18104 19737
rect 2688 19660 2740 19712
rect 3148 19660 3200 19712
rect 4804 19660 4856 19712
rect 5632 19660 5684 19712
rect 8024 19660 8076 19712
rect 10324 19703 10376 19712
rect 10324 19669 10333 19703
rect 10333 19669 10367 19703
rect 10367 19669 10376 19703
rect 10324 19660 10376 19669
rect 11244 19660 11296 19712
rect 12716 19660 12768 19712
rect 14372 19660 14424 19712
rect 15292 19660 15344 19712
rect 16488 19703 16540 19712
rect 16488 19669 16497 19703
rect 16497 19669 16531 19703
rect 16531 19669 16540 19703
rect 16488 19660 16540 19669
rect 3972 19558 4024 19610
rect 4036 19558 4088 19610
rect 4100 19558 4152 19610
rect 4164 19558 4216 19610
rect 9952 19558 10004 19610
rect 10016 19558 10068 19610
rect 10080 19558 10132 19610
rect 10144 19558 10196 19610
rect 15932 19558 15984 19610
rect 15996 19558 16048 19610
rect 16060 19558 16112 19610
rect 16124 19558 16176 19610
rect 1584 19456 1636 19508
rect 3700 19320 3752 19372
rect 8024 19363 8076 19372
rect 1860 19295 1912 19304
rect 1860 19261 1869 19295
rect 1869 19261 1903 19295
rect 1903 19261 1912 19295
rect 2412 19295 2464 19304
rect 1860 19252 1912 19261
rect 2412 19261 2421 19295
rect 2421 19261 2455 19295
rect 2455 19261 2464 19295
rect 2412 19252 2464 19261
rect 3976 19252 4028 19304
rect 940 19184 992 19236
rect 2964 19184 3016 19236
rect 3332 19184 3384 19236
rect 4528 19116 4580 19168
rect 5908 19159 5960 19168
rect 5908 19125 5917 19159
rect 5917 19125 5951 19159
rect 5951 19125 5960 19159
rect 5908 19116 5960 19125
rect 6000 19116 6052 19168
rect 7104 19295 7156 19304
rect 7104 19261 7113 19295
rect 7113 19261 7147 19295
rect 7147 19261 7156 19295
rect 7104 19252 7156 19261
rect 7564 19252 7616 19304
rect 8024 19329 8033 19363
rect 8033 19329 8067 19363
rect 8067 19329 8076 19363
rect 8024 19320 8076 19329
rect 12808 19295 12860 19304
rect 12808 19261 12817 19295
rect 12817 19261 12851 19295
rect 12851 19261 12860 19295
rect 12808 19252 12860 19261
rect 14924 19252 14976 19304
rect 17592 19252 17644 19304
rect 7380 19184 7432 19236
rect 7472 19116 7524 19168
rect 9036 19184 9088 19236
rect 9680 19184 9732 19236
rect 7748 19116 7800 19168
rect 7840 19116 7892 19168
rect 10600 19159 10652 19168
rect 10600 19125 10609 19159
rect 10609 19125 10643 19159
rect 10643 19125 10652 19159
rect 10600 19116 10652 19125
rect 13820 19184 13872 19236
rect 15752 19184 15804 19236
rect 17776 19184 17828 19236
rect 13268 19116 13320 19168
rect 13452 19116 13504 19168
rect 15476 19159 15528 19168
rect 15476 19125 15485 19159
rect 15485 19125 15519 19159
rect 15519 19125 15528 19159
rect 15476 19116 15528 19125
rect 17316 19159 17368 19168
rect 17316 19125 17325 19159
rect 17325 19125 17359 19159
rect 17359 19125 17368 19159
rect 17316 19116 17368 19125
rect 6962 19014 7014 19066
rect 7026 19014 7078 19066
rect 7090 19014 7142 19066
rect 7154 19014 7206 19066
rect 12942 19014 12994 19066
rect 13006 19014 13058 19066
rect 13070 19014 13122 19066
rect 13134 19014 13186 19066
rect 3332 18955 3384 18964
rect 3332 18921 3341 18955
rect 3341 18921 3375 18955
rect 3375 18921 3384 18955
rect 3332 18912 3384 18921
rect 6000 18912 6052 18964
rect 7288 18912 7340 18964
rect 7840 18912 7892 18964
rect 5908 18844 5960 18896
rect 2780 18776 2832 18828
rect 3976 18776 4028 18828
rect 4528 18776 4580 18828
rect 7748 18776 7800 18828
rect 8208 18912 8260 18964
rect 10600 18844 10652 18896
rect 8024 18819 8076 18828
rect 8024 18785 8033 18819
rect 8033 18785 8067 18819
rect 8067 18785 8076 18819
rect 8208 18819 8260 18828
rect 8024 18776 8076 18785
rect 8208 18785 8217 18819
rect 8217 18785 8251 18819
rect 8251 18785 8260 18819
rect 8208 18776 8260 18785
rect 9680 18819 9732 18828
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 13452 18912 13504 18964
rect 13820 18955 13872 18964
rect 13820 18921 13829 18955
rect 13829 18921 13863 18955
rect 13863 18921 13872 18955
rect 13820 18912 13872 18921
rect 13544 18844 13596 18896
rect 2412 18708 2464 18760
rect 4988 18751 5040 18760
rect 4988 18717 4997 18751
rect 4997 18717 5031 18751
rect 5031 18717 5040 18751
rect 4988 18708 5040 18717
rect 6552 18640 6604 18692
rect 7564 18640 7616 18692
rect 12164 18819 12216 18828
rect 12164 18785 12173 18819
rect 12173 18785 12207 18819
rect 12207 18785 12216 18819
rect 12164 18776 12216 18785
rect 12440 18819 12492 18828
rect 12440 18785 12449 18819
rect 12449 18785 12483 18819
rect 12483 18785 12492 18819
rect 12440 18776 12492 18785
rect 12348 18708 12400 18760
rect 12532 18708 12584 18760
rect 13176 18819 13228 18828
rect 13176 18785 13185 18819
rect 13185 18785 13219 18819
rect 13219 18785 13228 18819
rect 13176 18776 13228 18785
rect 14924 18844 14976 18896
rect 15292 18844 15344 18896
rect 15476 18844 15528 18896
rect 17132 18819 17184 18828
rect 17132 18785 17141 18819
rect 17141 18785 17175 18819
rect 17175 18785 17184 18819
rect 17132 18776 17184 18785
rect 12808 18708 12860 18760
rect 14648 18708 14700 18760
rect 16948 18751 17000 18760
rect 16948 18717 16957 18751
rect 16957 18717 16991 18751
rect 16991 18717 17000 18751
rect 16948 18708 17000 18717
rect 13268 18640 13320 18692
rect 4344 18615 4396 18624
rect 4344 18581 4353 18615
rect 4353 18581 4387 18615
rect 4387 18581 4396 18615
rect 4344 18572 4396 18581
rect 7656 18615 7708 18624
rect 7656 18581 7665 18615
rect 7665 18581 7699 18615
rect 7699 18581 7708 18615
rect 7656 18572 7708 18581
rect 12164 18572 12216 18624
rect 16304 18572 16356 18624
rect 18236 18572 18288 18624
rect 3972 18470 4024 18522
rect 4036 18470 4088 18522
rect 4100 18470 4152 18522
rect 4164 18470 4216 18522
rect 9952 18470 10004 18522
rect 10016 18470 10068 18522
rect 10080 18470 10132 18522
rect 10144 18470 10196 18522
rect 15932 18470 15984 18522
rect 15996 18470 16048 18522
rect 16060 18470 16112 18522
rect 16124 18470 16176 18522
rect 3700 18411 3752 18420
rect 3700 18377 3709 18411
rect 3709 18377 3743 18411
rect 3743 18377 3752 18411
rect 3700 18368 3752 18377
rect 9036 18411 9088 18420
rect 9036 18377 9045 18411
rect 9045 18377 9079 18411
rect 9079 18377 9088 18411
rect 9036 18368 9088 18377
rect 4344 18300 4396 18352
rect 4160 18275 4212 18284
rect 4160 18241 4169 18275
rect 4169 18241 4203 18275
rect 4203 18241 4212 18275
rect 4160 18232 4212 18241
rect 7288 18232 7340 18284
rect 4528 18164 4580 18216
rect 4620 18164 4672 18216
rect 7472 18164 7524 18216
rect 7840 18232 7892 18284
rect 12440 18368 12492 18420
rect 13176 18368 13228 18420
rect 17132 18368 17184 18420
rect 11704 18300 11756 18352
rect 18328 18343 18380 18352
rect 7932 18207 7984 18216
rect 7932 18173 7941 18207
rect 7941 18173 7975 18207
rect 7975 18173 7984 18207
rect 7932 18164 7984 18173
rect 8484 18207 8536 18216
rect 7840 18096 7892 18148
rect 8484 18173 8493 18207
rect 8493 18173 8527 18207
rect 8527 18173 8536 18207
rect 8484 18164 8536 18173
rect 12164 18232 12216 18284
rect 18328 18309 18337 18343
rect 18337 18309 18371 18343
rect 18371 18309 18380 18343
rect 18328 18300 18380 18309
rect 16948 18232 17000 18284
rect 4344 18028 4396 18080
rect 6828 18071 6880 18080
rect 6828 18037 6837 18071
rect 6837 18037 6871 18071
rect 6871 18037 6880 18071
rect 6828 18028 6880 18037
rect 7472 18028 7524 18080
rect 12164 18096 12216 18148
rect 14188 18164 14240 18216
rect 14648 18207 14700 18216
rect 14648 18173 14657 18207
rect 14657 18173 14691 18207
rect 14691 18173 14700 18207
rect 14648 18164 14700 18173
rect 13452 18139 13504 18148
rect 13452 18105 13461 18139
rect 13461 18105 13495 18139
rect 13495 18105 13504 18139
rect 13452 18096 13504 18105
rect 13544 18139 13596 18148
rect 13544 18105 13553 18139
rect 13553 18105 13587 18139
rect 13587 18105 13596 18139
rect 13544 18096 13596 18105
rect 17960 18096 18012 18148
rect 18420 18096 18472 18148
rect 11796 18028 11848 18080
rect 12624 18028 12676 18080
rect 12808 18028 12860 18080
rect 6962 17926 7014 17978
rect 7026 17926 7078 17978
rect 7090 17926 7142 17978
rect 7154 17926 7206 17978
rect 12942 17926 12994 17978
rect 13006 17926 13058 17978
rect 13070 17926 13122 17978
rect 13134 17926 13186 17978
rect 4988 17824 5040 17876
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 2780 17688 2832 17697
rect 4528 17688 4580 17740
rect 5448 17688 5500 17740
rect 6552 17824 6604 17876
rect 6828 17824 6880 17876
rect 7932 17824 7984 17876
rect 11796 17731 11848 17740
rect 7656 17620 7708 17672
rect 9680 17620 9732 17672
rect 11796 17697 11805 17731
rect 11805 17697 11839 17731
rect 11839 17697 11848 17731
rect 11796 17688 11848 17697
rect 12624 17824 12676 17876
rect 16948 17824 17000 17876
rect 17960 17867 18012 17876
rect 17960 17833 17969 17867
rect 17969 17833 18003 17867
rect 18003 17833 18012 17867
rect 17960 17824 18012 17833
rect 12808 17756 12860 17808
rect 16304 17756 16356 17808
rect 17316 17756 17368 17808
rect 11704 17663 11756 17672
rect 11704 17629 11713 17663
rect 11713 17629 11747 17663
rect 11747 17629 11756 17663
rect 11704 17620 11756 17629
rect 12164 17688 12216 17740
rect 13452 17688 13504 17740
rect 14740 17688 14792 17740
rect 14924 17731 14976 17740
rect 14924 17697 14933 17731
rect 14933 17697 14967 17731
rect 14967 17697 14976 17731
rect 14924 17688 14976 17697
rect 18512 17688 18564 17740
rect 12716 17620 12768 17672
rect 14188 17620 14240 17672
rect 2596 17527 2648 17536
rect 2596 17493 2605 17527
rect 2605 17493 2639 17527
rect 2639 17493 2648 17527
rect 2596 17484 2648 17493
rect 3700 17484 3752 17536
rect 13544 17552 13596 17604
rect 6000 17484 6052 17536
rect 9772 17484 9824 17536
rect 10416 17484 10468 17536
rect 14832 17484 14884 17536
rect 3972 17382 4024 17434
rect 4036 17382 4088 17434
rect 4100 17382 4152 17434
rect 4164 17382 4216 17434
rect 9952 17382 10004 17434
rect 10016 17382 10068 17434
rect 10080 17382 10132 17434
rect 10144 17382 10196 17434
rect 15932 17382 15984 17434
rect 15996 17382 16048 17434
rect 16060 17382 16112 17434
rect 16124 17382 16176 17434
rect 5448 17323 5500 17332
rect 5448 17289 5457 17323
rect 5457 17289 5491 17323
rect 5491 17289 5500 17323
rect 5448 17280 5500 17289
rect 3700 17076 3752 17128
rect 1860 17008 1912 17060
rect 2596 17008 2648 17060
rect 4068 17051 4120 17060
rect 4068 17017 4077 17051
rect 4077 17017 4111 17051
rect 4111 17017 4120 17051
rect 4068 17008 4120 17017
rect 4160 17051 4212 17060
rect 4160 17017 4169 17051
rect 4169 17017 4203 17051
rect 4203 17017 4212 17051
rect 4988 17187 5040 17196
rect 4988 17153 4997 17187
rect 4997 17153 5031 17187
rect 5031 17153 5040 17187
rect 4988 17144 5040 17153
rect 4620 17076 4672 17128
rect 4896 17119 4948 17128
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 5172 17119 5224 17128
rect 5172 17085 5181 17119
rect 5181 17085 5215 17119
rect 5215 17085 5224 17119
rect 5172 17076 5224 17085
rect 9680 17187 9732 17196
rect 5448 17076 5500 17128
rect 9680 17153 9689 17187
rect 9689 17153 9723 17187
rect 9723 17153 9732 17187
rect 9680 17144 9732 17153
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 10416 17144 10468 17196
rect 7472 17119 7524 17128
rect 7472 17085 7481 17119
rect 7481 17085 7515 17119
rect 7515 17085 7524 17119
rect 7472 17076 7524 17085
rect 7748 17076 7800 17128
rect 8484 17076 8536 17128
rect 4160 17008 4212 17017
rect 8300 17008 8352 17060
rect 10784 17119 10836 17128
rect 10784 17085 10793 17119
rect 10793 17085 10827 17119
rect 10827 17085 10836 17119
rect 12348 17119 12400 17128
rect 10784 17076 10836 17085
rect 12348 17085 12357 17119
rect 12357 17085 12391 17119
rect 12391 17085 12400 17119
rect 12348 17076 12400 17085
rect 13452 17212 13504 17264
rect 16120 17212 16172 17264
rect 16856 17212 16908 17264
rect 12808 17144 12860 17196
rect 14464 17144 14516 17196
rect 12716 17119 12768 17128
rect 12716 17085 12725 17119
rect 12725 17085 12759 17119
rect 12759 17085 12768 17119
rect 12716 17076 12768 17085
rect 13360 17076 13412 17128
rect 13544 17119 13596 17128
rect 13544 17085 13553 17119
rect 13553 17085 13587 17119
rect 13587 17085 13596 17119
rect 13544 17076 13596 17085
rect 17224 17144 17276 17196
rect 4528 16940 4580 16992
rect 6368 16940 6420 16992
rect 7564 16940 7616 16992
rect 10784 16940 10836 16992
rect 14832 17008 14884 17060
rect 16396 17076 16448 17128
rect 17776 17076 17828 17128
rect 17684 17008 17736 17060
rect 6962 16838 7014 16890
rect 7026 16838 7078 16890
rect 7090 16838 7142 16890
rect 7154 16838 7206 16890
rect 12942 16838 12994 16890
rect 13006 16838 13058 16890
rect 13070 16838 13122 16890
rect 13134 16838 13186 16890
rect 5172 16736 5224 16788
rect 5816 16736 5868 16788
rect 6828 16736 6880 16788
rect 4896 16668 4948 16720
rect 7564 16668 7616 16720
rect 12808 16736 12860 16788
rect 13544 16736 13596 16788
rect 14188 16736 14240 16788
rect 15384 16779 15436 16788
rect 15384 16745 15393 16779
rect 15393 16745 15427 16779
rect 15427 16745 15436 16779
rect 15384 16736 15436 16745
rect 5448 16643 5500 16652
rect 5448 16609 5457 16643
rect 5457 16609 5491 16643
rect 5491 16609 5500 16643
rect 5448 16600 5500 16609
rect 9772 16600 9824 16652
rect 10416 16668 10468 16720
rect 12716 16668 12768 16720
rect 16396 16736 16448 16788
rect 10508 16643 10560 16652
rect 4068 16532 4120 16584
rect 6368 16532 6420 16584
rect 6552 16575 6604 16584
rect 6552 16541 6561 16575
rect 6561 16541 6595 16575
rect 6595 16541 6604 16575
rect 6552 16532 6604 16541
rect 6920 16532 6972 16584
rect 10508 16609 10517 16643
rect 10517 16609 10551 16643
rect 10551 16609 10560 16643
rect 10508 16600 10560 16609
rect 10784 16643 10836 16652
rect 10784 16609 10793 16643
rect 10793 16609 10827 16643
rect 10827 16609 10836 16643
rect 10784 16600 10836 16609
rect 10416 16532 10468 16584
rect 12348 16600 12400 16652
rect 13360 16643 13412 16652
rect 13360 16609 13369 16643
rect 13369 16609 13403 16643
rect 13403 16609 13412 16643
rect 13360 16600 13412 16609
rect 14648 16600 14700 16652
rect 18144 16668 18196 16720
rect 15752 16600 15804 16652
rect 16120 16643 16172 16652
rect 16120 16609 16129 16643
rect 16129 16609 16163 16643
rect 16163 16609 16172 16643
rect 16120 16600 16172 16609
rect 12164 16532 12216 16584
rect 14464 16532 14516 16584
rect 5080 16464 5132 16516
rect 14188 16464 14240 16516
rect 16948 16532 17000 16584
rect 4988 16396 5040 16448
rect 5724 16396 5776 16448
rect 7840 16396 7892 16448
rect 12256 16439 12308 16448
rect 12256 16405 12265 16439
rect 12265 16405 12299 16439
rect 12299 16405 12308 16439
rect 12256 16396 12308 16405
rect 18328 16439 18380 16448
rect 18328 16405 18337 16439
rect 18337 16405 18371 16439
rect 18371 16405 18380 16439
rect 18328 16396 18380 16405
rect 3972 16294 4024 16346
rect 4036 16294 4088 16346
rect 4100 16294 4152 16346
rect 4164 16294 4216 16346
rect 9952 16294 10004 16346
rect 10016 16294 10068 16346
rect 10080 16294 10132 16346
rect 10144 16294 10196 16346
rect 15932 16294 15984 16346
rect 15996 16294 16048 16346
rect 16060 16294 16112 16346
rect 16124 16294 16176 16346
rect 5816 16235 5868 16244
rect 5816 16201 5825 16235
rect 5825 16201 5859 16235
rect 5859 16201 5868 16235
rect 5816 16192 5868 16201
rect 6920 16235 6972 16244
rect 6920 16201 6929 16235
rect 6929 16201 6963 16235
rect 6963 16201 6972 16235
rect 6920 16192 6972 16201
rect 8576 16192 8628 16244
rect 9588 16192 9640 16244
rect 1860 16099 1912 16108
rect 1860 16065 1869 16099
rect 1869 16065 1903 16099
rect 1903 16065 1912 16099
rect 1860 16056 1912 16065
rect 4712 16056 4764 16108
rect 5080 15988 5132 16040
rect 5724 16031 5776 16040
rect 5724 15997 5733 16031
rect 5733 15997 5767 16031
rect 5767 15997 5776 16031
rect 5724 15988 5776 15997
rect 6828 15988 6880 16040
rect 8208 16056 8260 16108
rect 9496 16099 9548 16108
rect 9496 16065 9505 16099
rect 9505 16065 9539 16099
rect 9539 16065 9548 16099
rect 9496 16056 9548 16065
rect 9864 16056 9916 16108
rect 2872 15920 2924 15972
rect 4988 15963 5040 15972
rect 4988 15929 4997 15963
rect 4997 15929 5031 15963
rect 5031 15929 5040 15963
rect 4988 15920 5040 15929
rect 3516 15852 3568 15904
rect 4436 15852 4488 15904
rect 8300 15988 8352 16040
rect 8576 16031 8628 16040
rect 8576 15997 8585 16031
rect 8585 15997 8619 16031
rect 8619 15997 8628 16031
rect 8576 15988 8628 15997
rect 9404 16031 9456 16040
rect 9404 15997 9413 16031
rect 9413 15997 9447 16031
rect 9447 15997 9456 16031
rect 9404 15988 9456 15997
rect 9588 15988 9640 16040
rect 10232 16031 10284 16040
rect 7196 15963 7248 15972
rect 7196 15929 7205 15963
rect 7205 15929 7239 15963
rect 7239 15929 7248 15963
rect 7196 15920 7248 15929
rect 7840 15920 7892 15972
rect 10232 15997 10241 16031
rect 10241 15997 10275 16031
rect 10275 15997 10284 16031
rect 10232 15988 10284 15997
rect 11152 15988 11204 16040
rect 12532 16056 12584 16108
rect 12164 15988 12216 16040
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 13544 15988 13596 16040
rect 15752 16124 15804 16176
rect 17224 16192 17276 16244
rect 17776 16124 17828 16176
rect 14464 15988 14516 16040
rect 14832 15988 14884 16040
rect 14924 15988 14976 16040
rect 16212 16031 16264 16040
rect 16212 15997 16221 16031
rect 16221 15997 16255 16031
rect 16255 15997 16264 16031
rect 16212 15988 16264 15997
rect 17500 16031 17552 16040
rect 17500 15997 17509 16031
rect 17509 15997 17543 16031
rect 17543 15997 17552 16031
rect 17500 15988 17552 15997
rect 17592 15988 17644 16040
rect 12348 15963 12400 15972
rect 12348 15929 12357 15963
rect 12357 15929 12391 15963
rect 12391 15929 12400 15963
rect 12348 15920 12400 15929
rect 14004 15920 14056 15972
rect 14648 15963 14700 15972
rect 14648 15929 14657 15963
rect 14657 15929 14691 15963
rect 14691 15929 14700 15963
rect 14648 15920 14700 15929
rect 7564 15852 7616 15904
rect 11980 15852 12032 15904
rect 13452 15852 13504 15904
rect 15016 15852 15068 15904
rect 15568 15895 15620 15904
rect 15568 15861 15577 15895
rect 15577 15861 15611 15895
rect 15611 15861 15620 15895
rect 15568 15852 15620 15861
rect 17040 15852 17092 15904
rect 17408 15852 17460 15904
rect 6962 15750 7014 15802
rect 7026 15750 7078 15802
rect 7090 15750 7142 15802
rect 7154 15750 7206 15802
rect 12942 15750 12994 15802
rect 13006 15750 13058 15802
rect 13070 15750 13122 15802
rect 13134 15750 13186 15802
rect 2872 15648 2924 15700
rect 3516 15648 3568 15700
rect 7564 15691 7616 15700
rect 7564 15657 7573 15691
rect 7573 15657 7607 15691
rect 7607 15657 7616 15691
rect 7564 15648 7616 15657
rect 10508 15648 10560 15700
rect 11980 15648 12032 15700
rect 4528 15623 4580 15632
rect 4528 15589 4537 15623
rect 4537 15589 4571 15623
rect 4571 15589 4580 15623
rect 4528 15580 4580 15589
rect 5540 15623 5592 15632
rect 5540 15589 5549 15623
rect 5549 15589 5583 15623
rect 5583 15589 5592 15623
rect 5540 15580 5592 15589
rect 10232 15580 10284 15632
rect 14096 15648 14148 15700
rect 14924 15648 14976 15700
rect 16948 15691 17000 15700
rect 16948 15657 16957 15691
rect 16957 15657 16991 15691
rect 16991 15657 17000 15691
rect 16948 15648 17000 15657
rect 13452 15623 13504 15632
rect 13452 15589 13461 15623
rect 13461 15589 13495 15623
rect 13495 15589 13504 15623
rect 13452 15580 13504 15589
rect 15016 15623 15068 15632
rect 15016 15589 15025 15623
rect 15025 15589 15059 15623
rect 15059 15589 15068 15623
rect 15016 15580 15068 15589
rect 15568 15580 15620 15632
rect 18236 15648 18288 15700
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 2780 15555 2832 15564
rect 2780 15521 2789 15555
rect 2789 15521 2823 15555
rect 2823 15521 2832 15555
rect 4436 15555 4488 15564
rect 2780 15512 2832 15521
rect 4436 15521 4445 15555
rect 4445 15521 4479 15555
rect 4479 15521 4488 15555
rect 4436 15512 4488 15521
rect 4344 15444 4396 15496
rect 4712 15555 4764 15564
rect 4712 15521 4747 15555
rect 4747 15521 4764 15555
rect 4712 15512 4764 15521
rect 4620 15376 4672 15428
rect 5172 15512 5224 15564
rect 5724 15555 5776 15564
rect 5724 15521 5733 15555
rect 5733 15521 5767 15555
rect 5767 15521 5776 15555
rect 5724 15512 5776 15521
rect 7656 15555 7708 15564
rect 5080 15444 5132 15496
rect 7656 15521 7665 15555
rect 7665 15521 7699 15555
rect 7699 15521 7708 15555
rect 7656 15512 7708 15521
rect 9680 15555 9732 15564
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 12164 15512 12216 15564
rect 17132 15555 17184 15564
rect 17132 15521 17141 15555
rect 17141 15521 17175 15555
rect 17175 15521 17184 15555
rect 17132 15512 17184 15521
rect 7932 15444 7984 15496
rect 9404 15444 9456 15496
rect 12256 15444 12308 15496
rect 14188 15444 14240 15496
rect 17776 15512 17828 15564
rect 18328 15512 18380 15564
rect 12072 15376 12124 15428
rect 1768 15308 1820 15360
rect 9496 15308 9548 15360
rect 11060 15308 11112 15360
rect 11980 15351 12032 15360
rect 11980 15317 11989 15351
rect 11989 15317 12023 15351
rect 12023 15317 12032 15351
rect 11980 15308 12032 15317
rect 16304 15308 16356 15360
rect 17592 15308 17644 15360
rect 3972 15206 4024 15258
rect 4036 15206 4088 15258
rect 4100 15206 4152 15258
rect 4164 15206 4216 15258
rect 9952 15206 10004 15258
rect 10016 15206 10068 15258
rect 10080 15206 10132 15258
rect 10144 15206 10196 15258
rect 15932 15206 15984 15258
rect 15996 15206 16048 15258
rect 16060 15206 16112 15258
rect 16124 15206 16176 15258
rect 4988 15104 5040 15156
rect 5264 15104 5316 15156
rect 5724 15104 5776 15156
rect 7656 15104 7708 15156
rect 9680 15147 9732 15156
rect 4712 14900 4764 14952
rect 5080 14900 5132 14952
rect 5816 14968 5868 15020
rect 6828 14900 6880 14952
rect 9680 15113 9689 15147
rect 9689 15113 9723 15147
rect 9723 15113 9732 15147
rect 9680 15104 9732 15113
rect 18144 15147 18196 15156
rect 18144 15113 18153 15147
rect 18153 15113 18187 15147
rect 18187 15113 18196 15147
rect 18144 15104 18196 15113
rect 14464 15079 14516 15088
rect 14464 15045 14473 15079
rect 14473 15045 14507 15079
rect 14507 15045 14516 15079
rect 14464 15036 14516 15045
rect 17500 15036 17552 15088
rect 8116 14900 8168 14952
rect 10416 14968 10468 15020
rect 11980 14968 12032 15020
rect 5816 14832 5868 14884
rect 7472 14875 7524 14884
rect 7472 14841 7481 14875
rect 7481 14841 7515 14875
rect 7515 14841 7524 14875
rect 7472 14832 7524 14841
rect 7840 14832 7892 14884
rect 7932 14832 7984 14884
rect 10876 14900 10928 14952
rect 12256 14943 12308 14952
rect 12256 14909 12265 14943
rect 12265 14909 12299 14943
rect 12299 14909 12308 14943
rect 12256 14900 12308 14909
rect 14648 14943 14700 14952
rect 14648 14909 14657 14943
rect 14657 14909 14691 14943
rect 14691 14909 14700 14943
rect 14648 14900 14700 14909
rect 14832 14968 14884 15020
rect 16212 14900 16264 14952
rect 17408 14943 17460 14952
rect 17408 14909 17417 14943
rect 17417 14909 17451 14943
rect 17451 14909 17460 14943
rect 17408 14900 17460 14909
rect 17592 14943 17644 14952
rect 17592 14909 17601 14943
rect 17601 14909 17635 14943
rect 17635 14909 17644 14943
rect 17592 14900 17644 14909
rect 18512 14900 18564 14952
rect 10968 14875 11020 14884
rect 10968 14841 10977 14875
rect 10977 14841 11011 14875
rect 11011 14841 11020 14875
rect 10968 14832 11020 14841
rect 14464 14832 14516 14884
rect 15108 14832 15160 14884
rect 7288 14764 7340 14816
rect 11520 14764 11572 14816
rect 15200 14764 15252 14816
rect 6962 14662 7014 14714
rect 7026 14662 7078 14714
rect 7090 14662 7142 14714
rect 7154 14662 7206 14714
rect 12942 14662 12994 14714
rect 13006 14662 13058 14714
rect 13070 14662 13122 14714
rect 13134 14662 13186 14714
rect 10876 14560 10928 14612
rect 11520 14560 11572 14612
rect 14648 14560 14700 14612
rect 15752 14560 15804 14612
rect 16212 14603 16264 14612
rect 16212 14569 16221 14603
rect 16221 14569 16255 14603
rect 16255 14569 16264 14603
rect 16212 14560 16264 14569
rect 16856 14560 16908 14612
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 2688 14424 2740 14476
rect 3056 14467 3108 14476
rect 3056 14433 3065 14467
rect 3065 14433 3099 14467
rect 3099 14433 3108 14467
rect 3056 14424 3108 14433
rect 5080 14424 5132 14476
rect 5264 14424 5316 14476
rect 5540 14424 5592 14476
rect 5724 14424 5776 14476
rect 7472 14424 7524 14476
rect 7932 14467 7984 14476
rect 4528 14356 4580 14408
rect 2872 14288 2924 14340
rect 2596 14220 2648 14272
rect 4528 14263 4580 14272
rect 4528 14229 4537 14263
rect 4537 14229 4571 14263
rect 4571 14229 4580 14263
rect 4528 14220 4580 14229
rect 5816 14356 5868 14408
rect 6828 14356 6880 14408
rect 5540 14331 5592 14340
rect 5540 14297 5549 14331
rect 5549 14297 5583 14331
rect 5583 14297 5592 14331
rect 5540 14288 5592 14297
rect 7288 14356 7340 14408
rect 7932 14433 7941 14467
rect 7941 14433 7975 14467
rect 7975 14433 7984 14467
rect 7932 14424 7984 14433
rect 8116 14467 8168 14476
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 8116 14424 8168 14433
rect 9220 14424 9272 14476
rect 11060 14424 11112 14476
rect 11520 14467 11572 14476
rect 11520 14433 11529 14467
rect 11529 14433 11563 14467
rect 11563 14433 11572 14467
rect 11520 14424 11572 14433
rect 13360 14467 13412 14476
rect 13360 14433 13369 14467
rect 13369 14433 13403 14467
rect 13403 14433 13412 14467
rect 13360 14424 13412 14433
rect 15016 14467 15068 14476
rect 15016 14433 15025 14467
rect 15025 14433 15059 14467
rect 15059 14433 15068 14467
rect 15016 14424 15068 14433
rect 16304 14424 16356 14476
rect 17316 14560 17368 14612
rect 17684 14560 17736 14612
rect 5448 14220 5500 14272
rect 7656 14288 7708 14340
rect 7104 14263 7156 14272
rect 7104 14229 7113 14263
rect 7113 14229 7147 14263
rect 7147 14229 7156 14263
rect 11704 14356 11756 14408
rect 17500 14424 17552 14476
rect 17868 14424 17920 14476
rect 8024 14331 8076 14340
rect 8024 14297 8033 14331
rect 8033 14297 8067 14331
rect 8067 14297 8076 14331
rect 8024 14288 8076 14297
rect 7104 14220 7156 14229
rect 8392 14220 8444 14272
rect 9312 14220 9364 14272
rect 13268 14263 13320 14272
rect 13268 14229 13277 14263
rect 13277 14229 13311 14263
rect 13311 14229 13320 14263
rect 13268 14220 13320 14229
rect 3972 14118 4024 14170
rect 4036 14118 4088 14170
rect 4100 14118 4152 14170
rect 4164 14118 4216 14170
rect 9952 14118 10004 14170
rect 10016 14118 10068 14170
rect 10080 14118 10132 14170
rect 10144 14118 10196 14170
rect 15932 14118 15984 14170
rect 15996 14118 16048 14170
rect 16060 14118 16112 14170
rect 16124 14118 16176 14170
rect 3056 14059 3108 14068
rect 3056 14025 3065 14059
rect 3065 14025 3099 14059
rect 3099 14025 3108 14059
rect 3056 14016 3108 14025
rect 7472 14016 7524 14068
rect 8116 14016 8168 14068
rect 8208 14016 8260 14068
rect 11152 14016 11204 14068
rect 1676 13948 1728 14000
rect 5172 13948 5224 14000
rect 2596 13923 2648 13932
rect 2596 13889 2605 13923
rect 2605 13889 2639 13923
rect 2639 13889 2648 13923
rect 2596 13880 2648 13889
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 1492 13812 1544 13864
rect 2872 13812 2924 13864
rect 3056 13855 3108 13864
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3056 13812 3108 13821
rect 3240 13812 3292 13864
rect 4528 13812 4580 13864
rect 7104 13812 7156 13864
rect 7748 13880 7800 13932
rect 7564 13855 7616 13864
rect 7564 13821 7572 13855
rect 7572 13821 7606 13855
rect 7606 13821 7616 13855
rect 7564 13812 7616 13821
rect 8300 13880 8352 13932
rect 8024 13812 8076 13864
rect 9128 13855 9180 13864
rect 9128 13821 9135 13855
rect 9135 13821 9180 13855
rect 9128 13812 9180 13821
rect 9312 13855 9364 13864
rect 9312 13821 9321 13855
rect 9321 13821 9355 13855
rect 9355 13821 9364 13855
rect 9312 13812 9364 13821
rect 9496 13812 9548 13864
rect 10784 13812 10836 13864
rect 13360 13880 13412 13932
rect 14464 13880 14516 13932
rect 15108 13923 15160 13932
rect 15108 13889 15117 13923
rect 15117 13889 15151 13923
rect 15151 13889 15160 13923
rect 15108 13880 15160 13889
rect 4988 13787 5040 13796
rect 4988 13753 4997 13787
rect 4997 13753 5031 13787
rect 5031 13753 5040 13787
rect 4988 13744 5040 13753
rect 5540 13744 5592 13796
rect 9220 13787 9272 13796
rect 4804 13676 4856 13728
rect 6828 13676 6880 13728
rect 9220 13753 9229 13787
rect 9229 13753 9263 13787
rect 9263 13753 9272 13787
rect 9220 13744 9272 13753
rect 13912 13812 13964 13864
rect 14924 13855 14976 13864
rect 14924 13821 14933 13855
rect 14933 13821 14967 13855
rect 14967 13821 14976 13855
rect 14924 13812 14976 13821
rect 15016 13855 15068 13864
rect 15016 13821 15025 13855
rect 15025 13821 15059 13855
rect 15059 13821 15068 13855
rect 15200 13855 15252 13864
rect 15016 13812 15068 13821
rect 15200 13821 15209 13855
rect 15209 13821 15243 13855
rect 15243 13821 15252 13855
rect 15200 13812 15252 13821
rect 16396 13812 16448 13864
rect 17316 13855 17368 13864
rect 17316 13821 17325 13855
rect 17325 13821 17359 13855
rect 17359 13821 17368 13855
rect 17316 13812 17368 13821
rect 17500 13855 17552 13864
rect 17500 13821 17509 13855
rect 17509 13821 17543 13855
rect 17543 13821 17552 13855
rect 17500 13812 17552 13821
rect 17684 13855 17736 13864
rect 17684 13821 17693 13855
rect 17693 13821 17727 13855
rect 17727 13821 17736 13855
rect 17684 13812 17736 13821
rect 13728 13787 13780 13796
rect 13728 13753 13737 13787
rect 13737 13753 13771 13787
rect 13771 13753 13780 13787
rect 13728 13744 13780 13753
rect 15936 13787 15988 13796
rect 15936 13753 15945 13787
rect 15945 13753 15979 13787
rect 15979 13753 15988 13787
rect 15936 13744 15988 13753
rect 17592 13787 17644 13796
rect 17592 13753 17601 13787
rect 17601 13753 17635 13787
rect 17635 13753 17644 13787
rect 17592 13744 17644 13753
rect 10048 13719 10100 13728
rect 10048 13685 10057 13719
rect 10057 13685 10091 13719
rect 10091 13685 10100 13719
rect 10048 13676 10100 13685
rect 13820 13676 13872 13728
rect 14004 13676 14056 13728
rect 15108 13676 15160 13728
rect 17132 13676 17184 13728
rect 6962 13574 7014 13626
rect 7026 13574 7078 13626
rect 7090 13574 7142 13626
rect 7154 13574 7206 13626
rect 12942 13574 12994 13626
rect 13006 13574 13058 13626
rect 13070 13574 13122 13626
rect 13134 13574 13186 13626
rect 1492 13515 1544 13524
rect 1492 13481 1501 13515
rect 1501 13481 1535 13515
rect 1535 13481 1544 13515
rect 1492 13472 1544 13481
rect 3148 13472 3200 13524
rect 4988 13472 5040 13524
rect 7564 13472 7616 13524
rect 9128 13472 9180 13524
rect 11704 13472 11756 13524
rect 13728 13515 13780 13524
rect 2964 13404 3016 13456
rect 10048 13404 10100 13456
rect 11428 13404 11480 13456
rect 13728 13481 13737 13515
rect 13737 13481 13771 13515
rect 13771 13481 13780 13515
rect 13728 13472 13780 13481
rect 15016 13472 15068 13524
rect 15936 13472 15988 13524
rect 17316 13472 17368 13524
rect 17684 13515 17736 13524
rect 17684 13481 17693 13515
rect 17693 13481 17727 13515
rect 17727 13481 17736 13515
rect 17684 13472 17736 13481
rect 18328 13472 18380 13524
rect 2688 13379 2740 13388
rect 1584 13268 1636 13320
rect 2688 13345 2697 13379
rect 2697 13345 2731 13379
rect 2731 13345 2740 13379
rect 2688 13336 2740 13345
rect 3240 13379 3292 13388
rect 3240 13345 3249 13379
rect 3249 13345 3283 13379
rect 3283 13345 3292 13379
rect 3240 13336 3292 13345
rect 5540 13379 5592 13388
rect 4436 13268 4488 13320
rect 4804 13311 4856 13320
rect 4804 13277 4813 13311
rect 4813 13277 4847 13311
rect 4847 13277 4856 13311
rect 4804 13268 4856 13277
rect 5540 13345 5549 13379
rect 5549 13345 5583 13379
rect 5583 13345 5592 13379
rect 5540 13336 5592 13345
rect 7472 13336 7524 13388
rect 7748 13379 7800 13388
rect 7748 13345 7757 13379
rect 7757 13345 7791 13379
rect 7791 13345 7800 13379
rect 7748 13336 7800 13345
rect 9496 13379 9548 13388
rect 9496 13345 9505 13379
rect 9505 13345 9539 13379
rect 9539 13345 9548 13379
rect 9496 13336 9548 13345
rect 5724 13268 5776 13320
rect 6828 13268 6880 13320
rect 4344 13200 4396 13252
rect 4528 13132 4580 13184
rect 7288 13200 7340 13252
rect 8208 13268 8260 13320
rect 10416 13268 10468 13320
rect 13268 13336 13320 13388
rect 13912 13404 13964 13456
rect 13820 13379 13872 13388
rect 13820 13345 13829 13379
rect 13829 13345 13863 13379
rect 13863 13345 13872 13379
rect 13820 13336 13872 13345
rect 15108 13379 15160 13388
rect 15108 13345 15117 13379
rect 15117 13345 15151 13379
rect 15151 13345 15160 13379
rect 15108 13336 15160 13345
rect 13728 13268 13780 13320
rect 15016 13311 15068 13320
rect 15016 13277 15025 13311
rect 15025 13277 15059 13311
rect 15059 13277 15068 13311
rect 15844 13336 15896 13388
rect 15016 13268 15068 13277
rect 15752 13200 15804 13252
rect 7840 13132 7892 13184
rect 8208 13132 8260 13184
rect 11060 13132 11112 13184
rect 15292 13132 15344 13184
rect 17684 13379 17736 13388
rect 16304 13200 16356 13252
rect 17132 13268 17184 13320
rect 17684 13345 17690 13379
rect 17690 13345 17724 13379
rect 17724 13345 17736 13379
rect 17684 13336 17736 13345
rect 18328 13132 18380 13184
rect 3972 13030 4024 13082
rect 4036 13030 4088 13082
rect 4100 13030 4152 13082
rect 4164 13030 4216 13082
rect 9952 13030 10004 13082
rect 10016 13030 10068 13082
rect 10080 13030 10132 13082
rect 10144 13030 10196 13082
rect 15932 13030 15984 13082
rect 15996 13030 16048 13082
rect 16060 13030 16112 13082
rect 16124 13030 16176 13082
rect 3056 12928 3108 12980
rect 5540 12928 5592 12980
rect 5908 12928 5960 12980
rect 7564 12971 7616 12980
rect 7564 12937 7573 12971
rect 7573 12937 7607 12971
rect 7607 12937 7616 12971
rect 7564 12928 7616 12937
rect 8024 12971 8076 12980
rect 8024 12937 8033 12971
rect 8033 12937 8067 12971
rect 8067 12937 8076 12971
rect 8024 12928 8076 12937
rect 14924 12971 14976 12980
rect 14924 12937 14933 12971
rect 14933 12937 14967 12971
rect 14967 12937 14976 12971
rect 14924 12928 14976 12937
rect 15292 12928 15344 12980
rect 3240 12860 3292 12912
rect 13544 12860 13596 12912
rect 15108 12860 15160 12912
rect 9772 12792 9824 12844
rect 2688 12724 2740 12776
rect 3148 12724 3200 12776
rect 5356 12767 5408 12776
rect 5356 12733 5365 12767
rect 5365 12733 5399 12767
rect 5399 12733 5408 12767
rect 5356 12724 5408 12733
rect 5448 12767 5500 12776
rect 5448 12733 5457 12767
rect 5457 12733 5491 12767
rect 5491 12733 5500 12767
rect 5724 12767 5776 12776
rect 5448 12724 5500 12733
rect 5724 12733 5733 12767
rect 5733 12733 5767 12767
rect 5767 12733 5776 12767
rect 5724 12724 5776 12733
rect 7472 12767 7524 12776
rect 7472 12733 7481 12767
rect 7481 12733 7515 12767
rect 7515 12733 7524 12767
rect 7472 12724 7524 12733
rect 7656 12724 7708 12776
rect 7840 12767 7892 12776
rect 7840 12733 7849 12767
rect 7849 12733 7883 12767
rect 7883 12733 7892 12767
rect 13912 12792 13964 12844
rect 7840 12724 7892 12733
rect 11520 12656 11572 12708
rect 10692 12588 10744 12640
rect 12440 12588 12492 12640
rect 13544 12724 13596 12776
rect 15016 12724 15068 12776
rect 15752 12767 15804 12776
rect 15752 12733 15761 12767
rect 15761 12733 15795 12767
rect 15795 12733 15804 12767
rect 15752 12724 15804 12733
rect 17132 12724 17184 12776
rect 17776 12724 17828 12776
rect 13820 12656 13872 12708
rect 14004 12588 14056 12640
rect 16856 12588 16908 12640
rect 17684 12699 17736 12708
rect 17684 12665 17693 12699
rect 17693 12665 17727 12699
rect 17727 12665 17736 12699
rect 17684 12656 17736 12665
rect 18328 12588 18380 12640
rect 6962 12486 7014 12538
rect 7026 12486 7078 12538
rect 7090 12486 7142 12538
rect 7154 12486 7206 12538
rect 12942 12486 12994 12538
rect 13006 12486 13058 12538
rect 13070 12486 13122 12538
rect 13134 12486 13186 12538
rect 8208 12384 8260 12436
rect 3148 12359 3200 12368
rect 3148 12325 3157 12359
rect 3157 12325 3191 12359
rect 3191 12325 3200 12359
rect 3148 12316 3200 12325
rect 4528 12359 4580 12368
rect 4528 12325 4537 12359
rect 4537 12325 4571 12359
rect 4571 12325 4580 12359
rect 4528 12316 4580 12325
rect 7656 12316 7708 12368
rect 2136 12248 2188 12300
rect 2964 12291 3016 12300
rect 2964 12257 2973 12291
rect 2973 12257 3007 12291
rect 3007 12257 3016 12291
rect 2964 12248 3016 12257
rect 5540 12248 5592 12300
rect 3148 12180 3200 12232
rect 5724 12180 5776 12232
rect 6276 12180 6328 12232
rect 5908 12112 5960 12164
rect 6920 12248 6972 12300
rect 8024 12248 8076 12300
rect 8208 12248 8260 12300
rect 8760 12248 8812 12300
rect 9404 12248 9456 12300
rect 11428 12384 11480 12436
rect 13912 12384 13964 12436
rect 18328 12427 18380 12436
rect 18328 12393 18337 12427
rect 18337 12393 18371 12427
rect 18371 12393 18380 12427
rect 18328 12384 18380 12393
rect 12440 12316 12492 12368
rect 13360 12316 13412 12368
rect 14924 12316 14976 12368
rect 16856 12359 16908 12368
rect 11152 12291 11204 12300
rect 7564 12180 7616 12232
rect 5264 12044 5316 12096
rect 8484 12112 8536 12164
rect 9588 12112 9640 12164
rect 9680 12112 9732 12164
rect 11152 12257 11161 12291
rect 11161 12257 11195 12291
rect 11195 12257 11204 12291
rect 11152 12248 11204 12257
rect 14004 12248 14056 12300
rect 16856 12325 16865 12359
rect 16865 12325 16899 12359
rect 16899 12325 16908 12359
rect 16856 12316 16908 12325
rect 17960 12248 18012 12300
rect 10416 12180 10468 12232
rect 14188 12180 14240 12232
rect 11060 12112 11112 12164
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 8300 12044 8352 12096
rect 9404 12044 9456 12096
rect 10784 12044 10836 12096
rect 15200 12044 15252 12096
rect 3972 11942 4024 11994
rect 4036 11942 4088 11994
rect 4100 11942 4152 11994
rect 4164 11942 4216 11994
rect 9952 11942 10004 11994
rect 10016 11942 10068 11994
rect 10080 11942 10132 11994
rect 10144 11942 10196 11994
rect 15932 11942 15984 11994
rect 15996 11942 16048 11994
rect 16060 11942 16112 11994
rect 16124 11942 16176 11994
rect 2136 11840 2188 11892
rect 1584 11747 1636 11756
rect 1584 11713 1593 11747
rect 1593 11713 1627 11747
rect 1627 11713 1636 11747
rect 1584 11704 1636 11713
rect 1768 11747 1820 11756
rect 1768 11713 1777 11747
rect 1777 11713 1811 11747
rect 1811 11713 1820 11747
rect 1768 11704 1820 11713
rect 2964 11840 3016 11892
rect 4436 11840 4488 11892
rect 5356 11840 5408 11892
rect 5540 11883 5592 11892
rect 5540 11849 5549 11883
rect 5549 11849 5583 11883
rect 5583 11849 5592 11883
rect 5540 11840 5592 11849
rect 6920 11840 6972 11892
rect 7196 11840 7248 11892
rect 7288 11840 7340 11892
rect 7840 11840 7892 11892
rect 9772 11840 9824 11892
rect 13360 11883 13412 11892
rect 13360 11849 13369 11883
rect 13369 11849 13403 11883
rect 13403 11849 13412 11883
rect 13360 11840 13412 11849
rect 17960 11883 18012 11892
rect 17960 11849 17969 11883
rect 17969 11849 18003 11883
rect 18003 11849 18012 11883
rect 17960 11840 18012 11849
rect 4988 11772 5040 11824
rect 3056 11679 3108 11688
rect 3056 11645 3065 11679
rect 3065 11645 3099 11679
rect 3099 11645 3108 11679
rect 3056 11636 3108 11645
rect 4620 11636 4672 11688
rect 8484 11772 8536 11824
rect 9496 11815 9548 11824
rect 9496 11781 9505 11815
rect 9505 11781 9539 11815
rect 9539 11781 9548 11815
rect 9496 11772 9548 11781
rect 5908 11704 5960 11756
rect 6552 11704 6604 11756
rect 7748 11704 7800 11756
rect 7840 11704 7892 11756
rect 9404 11747 9456 11756
rect 9128 11679 9180 11688
rect 4252 11568 4304 11620
rect 9128 11645 9137 11679
rect 9137 11645 9171 11679
rect 9171 11645 9180 11679
rect 9128 11636 9180 11645
rect 9404 11713 9413 11747
rect 9413 11713 9447 11747
rect 9447 11713 9456 11747
rect 9404 11704 9456 11713
rect 14464 11747 14516 11756
rect 14464 11713 14473 11747
rect 14473 11713 14507 11747
rect 14507 11713 14516 11747
rect 14464 11704 14516 11713
rect 15752 11704 15804 11756
rect 10324 11636 10376 11688
rect 10600 11679 10652 11688
rect 10600 11645 10609 11679
rect 10609 11645 10643 11679
rect 10643 11645 10652 11679
rect 10600 11636 10652 11645
rect 10784 11679 10836 11688
rect 10784 11645 10793 11679
rect 10793 11645 10827 11679
rect 10827 11645 10836 11679
rect 10784 11636 10836 11645
rect 11152 11636 11204 11688
rect 14004 11636 14056 11688
rect 14188 11679 14240 11688
rect 14188 11645 14197 11679
rect 14197 11645 14231 11679
rect 14231 11645 14240 11679
rect 14188 11636 14240 11645
rect 7380 11568 7432 11620
rect 7656 11568 7708 11620
rect 4896 11500 4948 11552
rect 11336 11568 11388 11620
rect 11152 11500 11204 11552
rect 15200 11568 15252 11620
rect 18512 11636 18564 11688
rect 17408 11500 17460 11552
rect 6962 11398 7014 11450
rect 7026 11398 7078 11450
rect 7090 11398 7142 11450
rect 7154 11398 7206 11450
rect 12942 11398 12994 11450
rect 13006 11398 13058 11450
rect 13070 11398 13122 11450
rect 13134 11398 13186 11450
rect 1492 11339 1544 11348
rect 1492 11305 1501 11339
rect 1501 11305 1535 11339
rect 1535 11305 1544 11339
rect 1492 11296 1544 11305
rect 3056 11296 3108 11348
rect 4252 11339 4304 11348
rect 4252 11305 4261 11339
rect 4261 11305 4295 11339
rect 4295 11305 4304 11339
rect 4252 11296 4304 11305
rect 5080 11296 5132 11348
rect 4528 11228 4580 11280
rect 7472 11296 7524 11348
rect 6276 11271 6328 11280
rect 6276 11237 6285 11271
rect 6285 11237 6319 11271
rect 6319 11237 6328 11271
rect 6276 11228 6328 11237
rect 10600 11296 10652 11348
rect 11336 11339 11388 11348
rect 11336 11305 11345 11339
rect 11345 11305 11379 11339
rect 11379 11305 11388 11339
rect 11336 11296 11388 11305
rect 12624 11296 12676 11348
rect 17684 11296 17736 11348
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 2780 11160 2832 11169
rect 4712 11160 4764 11212
rect 5080 11160 5132 11212
rect 5356 11160 5408 11212
rect 7196 11160 7248 11212
rect 7380 11160 7432 11212
rect 8208 11203 8260 11212
rect 8208 11169 8217 11203
rect 8217 11169 8251 11203
rect 8251 11169 8260 11203
rect 8208 11160 8260 11169
rect 9128 11228 9180 11280
rect 11060 11228 11112 11280
rect 16396 11271 16448 11280
rect 16396 11237 16405 11271
rect 16405 11237 16439 11271
rect 16439 11237 16448 11271
rect 16396 11228 16448 11237
rect 17408 11228 17460 11280
rect 11428 11203 11480 11212
rect 11428 11169 11437 11203
rect 11437 11169 11471 11203
rect 11471 11169 11480 11203
rect 11428 11160 11480 11169
rect 11520 11160 11572 11212
rect 12256 11160 12308 11212
rect 4896 11092 4948 11144
rect 9312 11092 9364 11144
rect 9680 11092 9732 11144
rect 11704 11092 11756 11144
rect 14188 11092 14240 11144
rect 14924 11092 14976 11144
rect 5724 11024 5776 11076
rect 5264 10956 5316 11008
rect 7196 11024 7248 11076
rect 7932 11024 7984 11076
rect 7288 10956 7340 11008
rect 8116 10956 8168 11008
rect 11520 10956 11572 11008
rect 12808 10999 12860 11008
rect 12808 10965 12817 10999
rect 12817 10965 12851 10999
rect 12851 10965 12860 10999
rect 12808 10956 12860 10965
rect 3972 10854 4024 10906
rect 4036 10854 4088 10906
rect 4100 10854 4152 10906
rect 4164 10854 4216 10906
rect 9952 10854 10004 10906
rect 10016 10854 10068 10906
rect 10080 10854 10132 10906
rect 10144 10854 10196 10906
rect 15932 10854 15984 10906
rect 15996 10854 16048 10906
rect 16060 10854 16112 10906
rect 16124 10854 16176 10906
rect 4620 10752 4672 10804
rect 5816 10795 5868 10804
rect 5816 10761 5825 10795
rect 5825 10761 5859 10795
rect 5859 10761 5868 10795
rect 5816 10752 5868 10761
rect 7932 10752 7984 10804
rect 11060 10795 11112 10804
rect 11060 10761 11069 10795
rect 11069 10761 11103 10795
rect 11103 10761 11112 10795
rect 11060 10752 11112 10761
rect 11428 10752 11480 10804
rect 4804 10684 4856 10736
rect 2412 10591 2464 10600
rect 2412 10557 2421 10591
rect 2421 10557 2455 10591
rect 2455 10557 2464 10591
rect 2412 10548 2464 10557
rect 3056 10548 3108 10600
rect 5080 10548 5132 10600
rect 5264 10480 5316 10532
rect 5356 10480 5408 10532
rect 7380 10548 7432 10600
rect 8116 10548 8168 10600
rect 8484 10548 8536 10600
rect 9404 10616 9456 10668
rect 11152 10616 11204 10668
rect 9128 10548 9180 10600
rect 11520 10616 11572 10668
rect 13544 10659 13596 10668
rect 13544 10625 13553 10659
rect 13553 10625 13587 10659
rect 13587 10625 13596 10659
rect 13544 10616 13596 10625
rect 9036 10523 9088 10532
rect 2780 10455 2832 10464
rect 2780 10421 2789 10455
rect 2789 10421 2823 10455
rect 2823 10421 2832 10455
rect 2780 10412 2832 10421
rect 4528 10412 4580 10464
rect 8760 10412 8812 10464
rect 9036 10489 9045 10523
rect 9045 10489 9079 10523
rect 9079 10489 9088 10523
rect 9036 10480 9088 10489
rect 9496 10412 9548 10464
rect 10324 10480 10376 10532
rect 10692 10523 10744 10532
rect 10692 10489 10701 10523
rect 10701 10489 10735 10523
rect 10735 10489 10744 10523
rect 10692 10480 10744 10489
rect 12808 10548 12860 10600
rect 14372 10548 14424 10600
rect 15108 10548 15160 10600
rect 15384 10591 15436 10600
rect 15384 10557 15393 10591
rect 15393 10557 15427 10591
rect 15427 10557 15436 10591
rect 15384 10548 15436 10557
rect 18328 10591 18380 10600
rect 18328 10557 18337 10591
rect 18337 10557 18371 10591
rect 18371 10557 18380 10591
rect 18328 10548 18380 10557
rect 15016 10480 15068 10532
rect 15292 10523 15344 10532
rect 15292 10489 15301 10523
rect 15301 10489 15335 10523
rect 15335 10489 15344 10523
rect 15292 10480 15344 10489
rect 13268 10412 13320 10464
rect 13452 10412 13504 10464
rect 16488 10412 16540 10464
rect 6962 10310 7014 10362
rect 7026 10310 7078 10362
rect 7090 10310 7142 10362
rect 7154 10310 7206 10362
rect 12942 10310 12994 10362
rect 13006 10310 13058 10362
rect 13070 10310 13122 10362
rect 13134 10310 13186 10362
rect 2412 10208 2464 10260
rect 17040 10251 17092 10260
rect 4804 10183 4856 10192
rect 4804 10149 4813 10183
rect 4813 10149 4847 10183
rect 4847 10149 4856 10183
rect 4804 10140 4856 10149
rect 5264 10140 5316 10192
rect 11152 10183 11204 10192
rect 3056 10072 3108 10124
rect 4712 10072 4764 10124
rect 5540 10072 5592 10124
rect 2780 9979 2832 9988
rect 2780 9945 2789 9979
rect 2789 9945 2823 9979
rect 2823 9945 2832 9979
rect 5356 10004 5408 10056
rect 6276 10072 6328 10124
rect 7196 10072 7248 10124
rect 8300 10115 8352 10124
rect 8300 10081 8309 10115
rect 8309 10081 8343 10115
rect 8343 10081 8352 10115
rect 8300 10072 8352 10081
rect 8392 10115 8444 10124
rect 8392 10081 8401 10115
rect 8401 10081 8435 10115
rect 8435 10081 8444 10115
rect 8392 10072 8444 10081
rect 9036 10072 9088 10124
rect 9588 10115 9640 10124
rect 9588 10081 9597 10115
rect 9597 10081 9631 10115
rect 9631 10081 9640 10115
rect 9588 10072 9640 10081
rect 11152 10149 11161 10183
rect 11161 10149 11195 10183
rect 11195 10149 11204 10183
rect 11152 10140 11204 10149
rect 12256 10115 12308 10124
rect 12256 10081 12265 10115
rect 12265 10081 12299 10115
rect 12299 10081 12308 10115
rect 12256 10072 12308 10081
rect 2780 9936 2832 9945
rect 4436 9868 4488 9920
rect 5080 9868 5132 9920
rect 6644 10004 6696 10056
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 9496 10047 9548 10056
rect 9496 10013 9505 10047
rect 9505 10013 9539 10047
rect 9539 10013 9548 10047
rect 9496 10004 9548 10013
rect 11704 10004 11756 10056
rect 13452 10183 13504 10192
rect 13452 10149 13461 10183
rect 13461 10149 13495 10183
rect 13495 10149 13504 10183
rect 13452 10140 13504 10149
rect 15016 10140 15068 10192
rect 17040 10217 17049 10251
rect 17049 10217 17083 10251
rect 17083 10217 17092 10251
rect 17040 10208 17092 10217
rect 18144 10140 18196 10192
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 12532 10004 12584 10056
rect 16948 10072 17000 10124
rect 6828 9868 6880 9920
rect 7472 9911 7524 9920
rect 7472 9877 7481 9911
rect 7481 9877 7515 9911
rect 7515 9877 7524 9911
rect 15108 9979 15160 9988
rect 15108 9945 15117 9979
rect 15117 9945 15151 9979
rect 15151 9945 15160 9979
rect 15108 9936 15160 9945
rect 17500 9911 17552 9920
rect 7472 9868 7524 9877
rect 17500 9877 17509 9911
rect 17509 9877 17543 9911
rect 17543 9877 17552 9911
rect 17500 9868 17552 9877
rect 3972 9766 4024 9818
rect 4036 9766 4088 9818
rect 4100 9766 4152 9818
rect 4164 9766 4216 9818
rect 9952 9766 10004 9818
rect 10016 9766 10068 9818
rect 10080 9766 10132 9818
rect 10144 9766 10196 9818
rect 15932 9766 15984 9818
rect 15996 9766 16048 9818
rect 16060 9766 16112 9818
rect 16124 9766 16176 9818
rect 7564 9664 7616 9716
rect 4988 9596 5040 9648
rect 5540 9596 5592 9648
rect 7288 9596 7340 9648
rect 1584 9528 1636 9580
rect 18144 9639 18196 9648
rect 18144 9605 18153 9639
rect 18153 9605 18187 9639
rect 18187 9605 18196 9639
rect 18144 9596 18196 9605
rect 2872 9503 2924 9512
rect 2872 9469 2881 9503
rect 2881 9469 2915 9503
rect 2915 9469 2924 9503
rect 2872 9460 2924 9469
rect 3332 9460 3384 9512
rect 1676 9392 1728 9444
rect 2320 9392 2372 9444
rect 1860 9367 1912 9376
rect 1860 9333 1869 9367
rect 1869 9333 1903 9367
rect 1903 9333 1912 9367
rect 1860 9324 1912 9333
rect 1952 9324 2004 9376
rect 4344 9324 4396 9376
rect 4896 9503 4948 9512
rect 4896 9469 4905 9503
rect 4905 9469 4939 9503
rect 4939 9469 4948 9503
rect 8208 9528 8260 9580
rect 13268 9571 13320 9580
rect 4896 9460 4948 9469
rect 5356 9392 5408 9444
rect 6644 9460 6696 9512
rect 7288 9503 7340 9512
rect 7288 9469 7297 9503
rect 7297 9469 7331 9503
rect 7331 9469 7340 9503
rect 7288 9460 7340 9469
rect 8392 9460 8444 9512
rect 8668 9503 8720 9512
rect 8668 9469 8677 9503
rect 8677 9469 8711 9503
rect 8711 9469 8720 9503
rect 8668 9460 8720 9469
rect 5264 9324 5316 9376
rect 8484 9367 8536 9376
rect 8484 9333 8493 9367
rect 8493 9333 8527 9367
rect 8527 9333 8536 9367
rect 8484 9324 8536 9333
rect 8944 9503 8996 9512
rect 8944 9469 8953 9503
rect 8953 9469 8987 9503
rect 8987 9469 8996 9503
rect 13268 9537 13277 9571
rect 13277 9537 13311 9571
rect 13311 9537 13320 9571
rect 13268 9528 13320 9537
rect 15108 9528 15160 9580
rect 8944 9460 8996 9469
rect 12808 9460 12860 9512
rect 15384 9460 15436 9512
rect 18328 9503 18380 9512
rect 18328 9469 18337 9503
rect 18337 9469 18371 9503
rect 18371 9469 18380 9503
rect 18328 9460 18380 9469
rect 9680 9392 9732 9444
rect 10692 9392 10744 9444
rect 9496 9367 9548 9376
rect 9496 9333 9505 9367
rect 9505 9333 9539 9367
rect 9539 9333 9548 9367
rect 9496 9324 9548 9333
rect 12716 9324 12768 9376
rect 15292 9324 15344 9376
rect 6962 9222 7014 9274
rect 7026 9222 7078 9274
rect 7090 9222 7142 9274
rect 7154 9222 7206 9274
rect 12942 9222 12994 9274
rect 13006 9222 13058 9274
rect 13070 9222 13122 9274
rect 13134 9222 13186 9274
rect 1860 9120 1912 9172
rect 9588 9120 9640 9172
rect 11244 9163 11296 9172
rect 11244 9129 11253 9163
rect 11253 9129 11287 9163
rect 11287 9129 11296 9163
rect 11244 9120 11296 9129
rect 15292 9120 15344 9172
rect 17684 9120 17736 9172
rect 5816 9052 5868 9104
rect 2504 8984 2556 9036
rect 4896 8984 4948 9036
rect 5172 9027 5224 9036
rect 5172 8993 5204 9027
rect 5204 8993 5224 9027
rect 5172 8984 5224 8993
rect 5540 8984 5592 9036
rect 8668 9052 8720 9104
rect 9312 9052 9364 9104
rect 12716 9052 12768 9104
rect 15384 9052 15436 9104
rect 3332 8959 3384 8968
rect 3332 8925 3341 8959
rect 3341 8925 3375 8959
rect 3375 8925 3384 8959
rect 3332 8916 3384 8925
rect 4988 8916 5040 8968
rect 5264 8959 5316 8968
rect 5264 8925 5273 8959
rect 5273 8925 5307 8959
rect 5307 8925 5316 8959
rect 5264 8916 5316 8925
rect 6644 8959 6696 8968
rect 1400 8891 1452 8900
rect 1400 8857 1409 8891
rect 1409 8857 1443 8891
rect 1443 8857 1452 8891
rect 1400 8848 1452 8857
rect 4528 8780 4580 8832
rect 4620 8780 4672 8832
rect 6644 8925 6653 8959
rect 6653 8925 6687 8959
rect 6687 8925 6696 8959
rect 6644 8916 6696 8925
rect 7564 8984 7616 9036
rect 8208 8984 8260 9036
rect 11796 8984 11848 9036
rect 13268 8984 13320 9036
rect 16488 9027 16540 9036
rect 16488 8993 16497 9027
rect 16497 8993 16531 9027
rect 16531 8993 16540 9027
rect 16488 8984 16540 8993
rect 17500 8984 17552 9036
rect 17868 8984 17920 9036
rect 6552 8848 6604 8900
rect 9496 8916 9548 8968
rect 11704 8916 11756 8968
rect 9588 8848 9640 8900
rect 8024 8780 8076 8832
rect 9680 8823 9732 8832
rect 9680 8789 9689 8823
rect 9689 8789 9723 8823
rect 9723 8789 9732 8823
rect 9680 8780 9732 8789
rect 10324 8780 10376 8832
rect 10692 8780 10744 8832
rect 14464 8780 14516 8832
rect 15660 8823 15712 8832
rect 15660 8789 15669 8823
rect 15669 8789 15703 8823
rect 15703 8789 15712 8823
rect 15660 8780 15712 8789
rect 16580 8823 16632 8832
rect 16580 8789 16589 8823
rect 16589 8789 16623 8823
rect 16623 8789 16632 8823
rect 16580 8780 16632 8789
rect 3972 8678 4024 8730
rect 4036 8678 4088 8730
rect 4100 8678 4152 8730
rect 4164 8678 4216 8730
rect 9952 8678 10004 8730
rect 10016 8678 10068 8730
rect 10080 8678 10132 8730
rect 10144 8678 10196 8730
rect 15932 8678 15984 8730
rect 15996 8678 16048 8730
rect 16060 8678 16112 8730
rect 16124 8678 16176 8730
rect 2596 8576 2648 8628
rect 5448 8576 5500 8628
rect 9588 8576 9640 8628
rect 4344 8440 4396 8492
rect 5632 8483 5684 8492
rect 5632 8449 5641 8483
rect 5641 8449 5675 8483
rect 5675 8449 5684 8483
rect 5632 8440 5684 8449
rect 7564 8440 7616 8492
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 1952 8372 2004 8424
rect 2320 8372 2372 8424
rect 2688 8415 2740 8424
rect 2688 8381 2697 8415
rect 2697 8381 2731 8415
rect 2731 8381 2740 8415
rect 2688 8372 2740 8381
rect 3516 8372 3568 8424
rect 8300 8372 8352 8424
rect 8208 8304 8260 8356
rect 9404 8372 9456 8424
rect 12440 8508 12492 8560
rect 11796 8372 11848 8424
rect 12072 8415 12124 8424
rect 12072 8381 12081 8415
rect 12081 8381 12115 8415
rect 12115 8381 12124 8415
rect 12072 8372 12124 8381
rect 12808 8576 12860 8628
rect 15660 8508 15712 8560
rect 17684 8483 17736 8492
rect 17684 8449 17693 8483
rect 17693 8449 17727 8483
rect 17727 8449 17736 8483
rect 17684 8440 17736 8449
rect 14464 8415 14516 8424
rect 14464 8381 14473 8415
rect 14473 8381 14507 8415
rect 14507 8381 14516 8415
rect 14464 8372 14516 8381
rect 15384 8372 15436 8424
rect 17500 8372 17552 8424
rect 17868 8415 17920 8424
rect 17868 8381 17877 8415
rect 17877 8381 17911 8415
rect 17911 8381 17920 8415
rect 17868 8372 17920 8381
rect 10416 8304 10468 8356
rect 4344 8236 4396 8288
rect 4712 8236 4764 8288
rect 7288 8236 7340 8288
rect 8116 8279 8168 8288
rect 8116 8245 8125 8279
rect 8125 8245 8159 8279
rect 8159 8245 8168 8279
rect 8116 8236 8168 8245
rect 8484 8279 8536 8288
rect 8484 8245 8493 8279
rect 8493 8245 8527 8279
rect 8527 8245 8536 8279
rect 8484 8236 8536 8245
rect 16488 8304 16540 8356
rect 16580 8304 16632 8356
rect 6962 8134 7014 8186
rect 7026 8134 7078 8186
rect 7090 8134 7142 8186
rect 7154 8134 7206 8186
rect 12942 8134 12994 8186
rect 13006 8134 13058 8186
rect 13070 8134 13122 8186
rect 13134 8134 13186 8186
rect 2688 8075 2740 8084
rect 2688 8041 2697 8075
rect 2697 8041 2731 8075
rect 2731 8041 2740 8075
rect 2688 8032 2740 8041
rect 12072 8032 12124 8084
rect 13360 8032 13412 8084
rect 17684 8032 17736 8084
rect 2596 7964 2648 8016
rect 4620 8007 4672 8016
rect 2320 7896 2372 7948
rect 4620 7973 4629 8007
rect 4629 7973 4663 8007
rect 4663 7973 4672 8007
rect 4620 7964 4672 7973
rect 7748 7964 7800 8016
rect 7288 7939 7340 7948
rect 2412 7828 2464 7880
rect 7288 7905 7297 7939
rect 7297 7905 7331 7939
rect 7331 7905 7340 7939
rect 7288 7896 7340 7905
rect 9312 7896 9364 7948
rect 12256 7964 12308 8016
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 11796 7939 11848 7948
rect 11796 7905 11805 7939
rect 11805 7905 11839 7939
rect 11839 7905 11848 7939
rect 11796 7896 11848 7905
rect 12624 7896 12676 7948
rect 4344 7871 4396 7880
rect 4344 7837 4353 7871
rect 4353 7837 4387 7871
rect 4387 7837 4396 7871
rect 4344 7828 4396 7837
rect 15752 7828 15804 7880
rect 9772 7760 9824 7812
rect 13636 7760 13688 7812
rect 3240 7735 3292 7744
rect 3240 7701 3249 7735
rect 3249 7701 3283 7735
rect 3283 7701 3292 7735
rect 3240 7692 3292 7701
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 9680 7692 9732 7744
rect 12072 7692 12124 7744
rect 16304 7692 16356 7744
rect 3972 7590 4024 7642
rect 4036 7590 4088 7642
rect 4100 7590 4152 7642
rect 4164 7590 4216 7642
rect 9952 7590 10004 7642
rect 10016 7590 10068 7642
rect 10080 7590 10132 7642
rect 10144 7590 10196 7642
rect 15932 7590 15984 7642
rect 15996 7590 16048 7642
rect 16060 7590 16112 7642
rect 16124 7590 16176 7642
rect 13360 7531 13412 7540
rect 13360 7497 13369 7531
rect 13369 7497 13403 7531
rect 13403 7497 13412 7531
rect 13360 7488 13412 7497
rect 16304 7531 16356 7540
rect 16304 7497 16313 7531
rect 16313 7497 16347 7531
rect 16347 7497 16356 7531
rect 16304 7488 16356 7497
rect 11796 7420 11848 7472
rect 1768 7327 1820 7336
rect 1768 7293 1777 7327
rect 1777 7293 1811 7327
rect 1811 7293 1820 7327
rect 1768 7284 1820 7293
rect 2320 7327 2372 7336
rect 2320 7293 2329 7327
rect 2329 7293 2363 7327
rect 2363 7293 2372 7327
rect 2320 7284 2372 7293
rect 3332 7216 3384 7268
rect 2136 7148 2188 7200
rect 4528 7284 4580 7336
rect 6000 7284 6052 7336
rect 7380 7284 7432 7336
rect 7564 7327 7616 7336
rect 7564 7293 7573 7327
rect 7573 7293 7607 7327
rect 7607 7293 7616 7327
rect 7564 7284 7616 7293
rect 8760 7284 8812 7336
rect 12624 7284 12676 7336
rect 13452 7284 13504 7336
rect 14556 7284 14608 7336
rect 15752 7327 15804 7336
rect 15752 7293 15761 7327
rect 15761 7293 15795 7327
rect 15795 7293 15804 7327
rect 15752 7284 15804 7293
rect 16580 7284 16632 7336
rect 5172 7216 5224 7268
rect 5908 7259 5960 7268
rect 5908 7225 5917 7259
rect 5917 7225 5951 7259
rect 5951 7225 5960 7259
rect 5908 7216 5960 7225
rect 9128 7216 9180 7268
rect 6828 7148 6880 7200
rect 7932 7191 7984 7200
rect 7932 7157 7941 7191
rect 7941 7157 7975 7191
rect 7975 7157 7984 7191
rect 7932 7148 7984 7157
rect 8576 7148 8628 7200
rect 8760 7191 8812 7200
rect 8760 7157 8769 7191
rect 8769 7157 8803 7191
rect 8803 7157 8812 7191
rect 8760 7148 8812 7157
rect 6962 7046 7014 7098
rect 7026 7046 7078 7098
rect 7090 7046 7142 7098
rect 7154 7046 7206 7098
rect 12942 7046 12994 7098
rect 13006 7046 13058 7098
rect 13070 7046 13122 7098
rect 13134 7046 13186 7098
rect 2136 6987 2188 6996
rect 2136 6953 2145 6987
rect 2145 6953 2179 6987
rect 2179 6953 2188 6987
rect 2136 6944 2188 6953
rect 4344 6944 4396 6996
rect 1584 6876 1636 6928
rect 7564 6944 7616 6996
rect 12072 6987 12124 6996
rect 12072 6953 12081 6987
rect 12081 6953 12115 6987
rect 12115 6953 12124 6987
rect 12072 6944 12124 6953
rect 13360 6944 13412 6996
rect 13636 6987 13688 6996
rect 13636 6953 13645 6987
rect 13645 6953 13679 6987
rect 13679 6953 13688 6987
rect 13636 6944 13688 6953
rect 1584 6740 1636 6792
rect 4988 6919 5040 6928
rect 3240 6808 3292 6860
rect 4988 6885 4997 6919
rect 4997 6885 5031 6919
rect 5031 6885 5040 6919
rect 4988 6876 5040 6885
rect 15476 6876 15528 6928
rect 16304 6876 16356 6928
rect 4896 6808 4948 6860
rect 7380 6808 7432 6860
rect 8116 6808 8168 6860
rect 9312 6808 9364 6860
rect 9772 6808 9824 6860
rect 10876 6851 10928 6860
rect 1768 6715 1820 6724
rect 1768 6681 1777 6715
rect 1777 6681 1811 6715
rect 1811 6681 1820 6715
rect 8300 6740 8352 6792
rect 9128 6740 9180 6792
rect 10876 6817 10885 6851
rect 10885 6817 10919 6851
rect 10919 6817 10928 6851
rect 10876 6808 10928 6817
rect 11796 6783 11848 6792
rect 11796 6749 11805 6783
rect 11805 6749 11839 6783
rect 11839 6749 11848 6783
rect 11796 6740 11848 6749
rect 1768 6672 1820 6681
rect 13452 6808 13504 6860
rect 14832 6808 14884 6860
rect 14924 6808 14976 6860
rect 18328 6851 18380 6860
rect 18328 6817 18337 6851
rect 18337 6817 18371 6851
rect 18371 6817 18380 6851
rect 18328 6808 18380 6817
rect 14556 6740 14608 6792
rect 14648 6740 14700 6792
rect 3332 6647 3384 6656
rect 3332 6613 3341 6647
rect 3341 6613 3375 6647
rect 3375 6613 3384 6647
rect 3332 6604 3384 6613
rect 8576 6647 8628 6656
rect 8576 6613 8585 6647
rect 8585 6613 8619 6647
rect 8619 6613 8628 6647
rect 8576 6604 8628 6613
rect 12348 6604 12400 6656
rect 12716 6604 12768 6656
rect 14740 6647 14792 6656
rect 14740 6613 14749 6647
rect 14749 6613 14783 6647
rect 14783 6613 14792 6647
rect 14740 6604 14792 6613
rect 14832 6604 14884 6656
rect 3972 6502 4024 6554
rect 4036 6502 4088 6554
rect 4100 6502 4152 6554
rect 4164 6502 4216 6554
rect 9952 6502 10004 6554
rect 10016 6502 10068 6554
rect 10080 6502 10132 6554
rect 10144 6502 10196 6554
rect 15932 6502 15984 6554
rect 15996 6502 16048 6554
rect 16060 6502 16112 6554
rect 16124 6502 16176 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 2504 6332 2556 6384
rect 14740 6400 14792 6452
rect 12716 6375 12768 6384
rect 12716 6341 12725 6375
rect 12725 6341 12759 6375
rect 12759 6341 12768 6375
rect 12716 6332 12768 6341
rect 4436 6264 4488 6316
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 6644 6196 6696 6248
rect 8760 6264 8812 6316
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 8392 6239 8444 6248
rect 8392 6205 8401 6239
rect 8401 6205 8435 6239
rect 8435 6205 8444 6239
rect 8392 6196 8444 6205
rect 9128 6239 9180 6248
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 9312 6239 9364 6248
rect 9312 6205 9321 6239
rect 9321 6205 9355 6239
rect 9355 6205 9364 6239
rect 9312 6196 9364 6205
rect 9772 6196 9824 6248
rect 10784 6196 10836 6248
rect 12348 6239 12400 6248
rect 12348 6205 12357 6239
rect 12357 6205 12391 6239
rect 12391 6205 12400 6239
rect 12348 6196 12400 6205
rect 4068 6128 4120 6180
rect 5264 6103 5316 6112
rect 5264 6069 5273 6103
rect 5273 6069 5307 6103
rect 5307 6069 5316 6103
rect 5264 6060 5316 6069
rect 9496 6060 9548 6112
rect 12716 6103 12768 6112
rect 12716 6069 12725 6103
rect 12725 6069 12759 6103
rect 12759 6069 12768 6103
rect 12716 6060 12768 6069
rect 15936 6196 15988 6248
rect 16396 6332 16448 6384
rect 18052 6332 18104 6384
rect 17132 6196 17184 6248
rect 15568 6060 15620 6112
rect 15844 6103 15896 6112
rect 15844 6069 15853 6103
rect 15853 6069 15887 6103
rect 15887 6069 15896 6103
rect 15844 6060 15896 6069
rect 6962 5958 7014 6010
rect 7026 5958 7078 6010
rect 7090 5958 7142 6010
rect 7154 5958 7206 6010
rect 12942 5958 12994 6010
rect 13006 5958 13058 6010
rect 13070 5958 13122 6010
rect 13134 5958 13186 6010
rect 5264 5856 5316 5908
rect 6644 5899 6696 5908
rect 6644 5865 6653 5899
rect 6653 5865 6687 5899
rect 6687 5865 6696 5899
rect 6644 5856 6696 5865
rect 6828 5856 6880 5908
rect 8576 5899 8628 5908
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 10784 5899 10836 5908
rect 10784 5865 10793 5899
rect 10793 5865 10827 5899
rect 10827 5865 10836 5899
rect 10784 5856 10836 5865
rect 15476 5899 15528 5908
rect 15476 5865 15485 5899
rect 15485 5865 15519 5899
rect 15519 5865 15528 5899
rect 15476 5856 15528 5865
rect 17132 5899 17184 5908
rect 17132 5865 17141 5899
rect 17141 5865 17175 5899
rect 17175 5865 17184 5899
rect 17132 5856 17184 5865
rect 3056 5831 3108 5840
rect 3056 5797 3065 5831
rect 3065 5797 3099 5831
rect 3099 5797 3108 5831
rect 3056 5788 3108 5797
rect 4068 5788 4120 5840
rect 12716 5788 12768 5840
rect 3240 5763 3292 5772
rect 3240 5729 3249 5763
rect 3249 5729 3283 5763
rect 3283 5729 3292 5763
rect 3240 5720 3292 5729
rect 4436 5720 4488 5772
rect 5172 5763 5224 5772
rect 5172 5729 5181 5763
rect 5181 5729 5215 5763
rect 5215 5729 5224 5763
rect 5172 5720 5224 5729
rect 5448 5720 5500 5772
rect 5632 5695 5684 5704
rect 5632 5661 5641 5695
rect 5641 5661 5675 5695
rect 5675 5661 5684 5695
rect 5632 5652 5684 5661
rect 7564 5652 7616 5704
rect 8116 5720 8168 5772
rect 9312 5720 9364 5772
rect 10508 5720 10560 5772
rect 12348 5720 12400 5772
rect 13452 5720 13504 5772
rect 15844 5788 15896 5840
rect 15936 5788 15988 5840
rect 15108 5763 15160 5772
rect 15108 5729 15117 5763
rect 15117 5729 15151 5763
rect 15151 5729 15160 5763
rect 15108 5720 15160 5729
rect 15568 5720 15620 5772
rect 16304 5763 16356 5772
rect 15660 5652 15712 5704
rect 16304 5729 16313 5763
rect 16313 5729 16347 5763
rect 16347 5729 16356 5763
rect 16304 5720 16356 5729
rect 16488 5763 16540 5772
rect 16488 5729 16497 5763
rect 16497 5729 16531 5763
rect 16531 5729 16540 5763
rect 16488 5720 16540 5729
rect 5724 5516 5776 5568
rect 18144 5516 18196 5568
rect 3972 5414 4024 5466
rect 4036 5414 4088 5466
rect 4100 5414 4152 5466
rect 4164 5414 4216 5466
rect 9952 5414 10004 5466
rect 10016 5414 10068 5466
rect 10080 5414 10132 5466
rect 10144 5414 10196 5466
rect 15932 5414 15984 5466
rect 15996 5414 16048 5466
rect 16060 5414 16112 5466
rect 16124 5414 16176 5466
rect 15108 5312 15160 5364
rect 16304 5355 16356 5364
rect 16304 5321 16313 5355
rect 16313 5321 16347 5355
rect 16347 5321 16356 5355
rect 16304 5312 16356 5321
rect 3240 5108 3292 5160
rect 3332 5151 3384 5160
rect 3332 5117 3341 5151
rect 3341 5117 3375 5151
rect 3375 5117 3384 5151
rect 5448 5244 5500 5296
rect 8392 5244 8444 5296
rect 5264 5219 5316 5228
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 17132 5244 17184 5296
rect 3332 5108 3384 5117
rect 5172 5108 5224 5160
rect 6644 5108 6696 5160
rect 7380 5108 7432 5160
rect 9772 5108 9824 5160
rect 10876 5108 10928 5160
rect 11520 5108 11572 5160
rect 12716 5108 12768 5160
rect 12808 5108 12860 5160
rect 16396 5151 16448 5160
rect 16396 5117 16405 5151
rect 16405 5117 16439 5151
rect 16439 5117 16448 5151
rect 16396 5108 16448 5117
rect 16488 5108 16540 5160
rect 10692 5040 10744 5092
rect 16028 5040 16080 5092
rect 2412 4972 2464 5024
rect 7932 4972 7984 5024
rect 10508 5015 10560 5024
rect 10508 4981 10517 5015
rect 10517 4981 10551 5015
rect 10551 4981 10560 5015
rect 10508 4972 10560 4981
rect 12624 4972 12676 5024
rect 15476 5015 15528 5024
rect 15476 4981 15485 5015
rect 15485 4981 15519 5015
rect 15519 4981 15528 5015
rect 15476 4972 15528 4981
rect 16672 4972 16724 5024
rect 6962 4870 7014 4922
rect 7026 4870 7078 4922
rect 7090 4870 7142 4922
rect 7154 4870 7206 4922
rect 12942 4870 12994 4922
rect 13006 4870 13058 4922
rect 13070 4870 13122 4922
rect 13134 4870 13186 4922
rect 1492 4811 1544 4820
rect 1492 4777 1501 4811
rect 1501 4777 1535 4811
rect 1535 4777 1544 4811
rect 1492 4768 1544 4777
rect 5632 4811 5684 4820
rect 5632 4777 5641 4811
rect 5641 4777 5675 4811
rect 5675 4777 5684 4811
rect 5632 4768 5684 4777
rect 7932 4768 7984 4820
rect 10508 4743 10560 4752
rect 10508 4709 10517 4743
rect 10517 4709 10551 4743
rect 10551 4709 10560 4743
rect 10508 4700 10560 4709
rect 13636 4768 13688 4820
rect 16028 4811 16080 4820
rect 16028 4777 16037 4811
rect 16037 4777 16071 4811
rect 16071 4777 16080 4811
rect 16028 4768 16080 4777
rect 18144 4811 18196 4820
rect 18144 4777 18153 4811
rect 18153 4777 18187 4811
rect 18187 4777 18196 4811
rect 18144 4768 18196 4777
rect 13544 4700 13596 4752
rect 2412 4675 2464 4684
rect 2412 4641 2421 4675
rect 2421 4641 2455 4675
rect 2455 4641 2464 4675
rect 2412 4632 2464 4641
rect 5172 4632 5224 4684
rect 4344 4564 4396 4616
rect 2320 4471 2372 4480
rect 2320 4437 2329 4471
rect 2329 4437 2363 4471
rect 2363 4437 2372 4471
rect 2320 4428 2372 4437
rect 9772 4632 9824 4684
rect 11520 4632 11572 4684
rect 11796 4632 11848 4684
rect 12716 4632 12768 4684
rect 16396 4675 16448 4684
rect 16396 4641 16405 4675
rect 16405 4641 16439 4675
rect 16439 4641 16448 4675
rect 16396 4632 16448 4641
rect 18328 4675 18380 4684
rect 18328 4641 18337 4675
rect 18337 4641 18371 4675
rect 18371 4641 18380 4675
rect 18328 4632 18380 4641
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 7288 4564 7340 4573
rect 7656 4607 7708 4616
rect 7656 4573 7665 4607
rect 7665 4573 7699 4607
rect 7699 4573 7708 4607
rect 7656 4564 7708 4573
rect 11612 4607 11664 4616
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 12900 4607 12952 4616
rect 12900 4573 12909 4607
rect 12909 4573 12943 4607
rect 12943 4573 12952 4607
rect 12900 4564 12952 4573
rect 16672 4607 16724 4616
rect 13268 4539 13320 4548
rect 13268 4505 13277 4539
rect 13277 4505 13311 4539
rect 13311 4505 13320 4539
rect 13268 4496 13320 4505
rect 16672 4573 16681 4607
rect 16681 4573 16715 4607
rect 16715 4573 16724 4607
rect 16672 4564 16724 4573
rect 16580 4496 16632 4548
rect 18420 4496 18472 4548
rect 7380 4428 7432 4480
rect 3972 4326 4024 4378
rect 4036 4326 4088 4378
rect 4100 4326 4152 4378
rect 4164 4326 4216 4378
rect 9952 4326 10004 4378
rect 10016 4326 10068 4378
rect 10080 4326 10132 4378
rect 10144 4326 10196 4378
rect 15932 4326 15984 4378
rect 15996 4326 16048 4378
rect 16060 4326 16112 4378
rect 16124 4326 16176 4378
rect 7656 4267 7708 4276
rect 7656 4233 7665 4267
rect 7665 4233 7699 4267
rect 7699 4233 7708 4267
rect 7656 4224 7708 4233
rect 9772 4224 9824 4276
rect 12900 4224 12952 4276
rect 7564 4156 7616 4208
rect 9588 4156 9640 4208
rect 7380 4088 7432 4140
rect 7472 4020 7524 4072
rect 7656 4020 7708 4072
rect 8668 4063 8720 4072
rect 8668 4029 8677 4063
rect 8677 4029 8711 4063
rect 8711 4029 8720 4063
rect 8668 4020 8720 4029
rect 10324 4088 10376 4140
rect 11612 4156 11664 4208
rect 12716 4156 12768 4208
rect 12624 4088 12676 4140
rect 13636 4131 13688 4140
rect 13636 4097 13645 4131
rect 13645 4097 13679 4131
rect 13679 4097 13688 4131
rect 13636 4088 13688 4097
rect 12440 4063 12492 4072
rect 12440 4029 12449 4063
rect 12449 4029 12483 4063
rect 12483 4029 12492 4063
rect 12440 4020 12492 4029
rect 12900 4020 12952 4072
rect 13544 4020 13596 4072
rect 13360 3952 13412 4004
rect 13452 3952 13504 4004
rect 10784 3884 10836 3936
rect 15016 3884 15068 3936
rect 15108 3927 15160 3936
rect 15108 3893 15117 3927
rect 15117 3893 15151 3927
rect 15151 3893 15160 3927
rect 15108 3884 15160 3893
rect 6962 3782 7014 3834
rect 7026 3782 7078 3834
rect 7090 3782 7142 3834
rect 7154 3782 7206 3834
rect 12942 3782 12994 3834
rect 13006 3782 13058 3834
rect 13070 3782 13122 3834
rect 13134 3782 13186 3834
rect 6828 3680 6880 3732
rect 8392 3680 8444 3732
rect 11520 3723 11572 3732
rect 5816 3612 5868 3664
rect 7288 3655 7340 3664
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 4344 3587 4396 3596
rect 4344 3553 4353 3587
rect 4353 3553 4387 3587
rect 4387 3553 4396 3587
rect 4344 3544 4396 3553
rect 7288 3621 7297 3655
rect 7297 3621 7331 3655
rect 7331 3621 7340 3655
rect 7288 3612 7340 3621
rect 10508 3612 10560 3664
rect 11520 3689 11529 3723
rect 11529 3689 11563 3723
rect 11563 3689 11572 3723
rect 11520 3680 11572 3689
rect 13268 3723 13320 3732
rect 13268 3689 13277 3723
rect 13277 3689 13311 3723
rect 13311 3689 13320 3723
rect 13268 3680 13320 3689
rect 13360 3680 13412 3732
rect 18144 3680 18196 3732
rect 12532 3612 12584 3664
rect 15568 3612 15620 3664
rect 8668 3544 8720 3596
rect 10692 3544 10744 3596
rect 13544 3544 13596 3596
rect 15108 3587 15160 3596
rect 15108 3553 15117 3587
rect 15117 3553 15151 3587
rect 15151 3553 15160 3587
rect 15108 3544 15160 3553
rect 18328 3587 18380 3596
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 10324 3476 10376 3528
rect 12532 3476 12584 3528
rect 14740 3519 14792 3528
rect 14740 3485 14749 3519
rect 14749 3485 14783 3519
rect 14783 3485 14792 3519
rect 14740 3476 14792 3485
rect 8116 3340 8168 3392
rect 11060 3408 11112 3460
rect 15476 3408 15528 3460
rect 16580 3476 16632 3528
rect 18328 3553 18337 3587
rect 18337 3553 18371 3587
rect 18371 3553 18380 3587
rect 18328 3544 18380 3553
rect 12072 3340 12124 3392
rect 15108 3383 15160 3392
rect 15108 3349 15117 3383
rect 15117 3349 15151 3383
rect 15151 3349 15160 3383
rect 15108 3340 15160 3349
rect 17316 3340 17368 3392
rect 3972 3238 4024 3290
rect 4036 3238 4088 3290
rect 4100 3238 4152 3290
rect 4164 3238 4216 3290
rect 9952 3238 10004 3290
rect 10016 3238 10068 3290
rect 10080 3238 10132 3290
rect 10144 3238 10196 3290
rect 15932 3238 15984 3290
rect 15996 3238 16048 3290
rect 16060 3238 16112 3290
rect 16124 3238 16176 3290
rect 8392 3179 8444 3188
rect 8392 3145 8401 3179
rect 8401 3145 8435 3179
rect 8435 3145 8444 3179
rect 8392 3136 8444 3145
rect 10508 3179 10560 3188
rect 10508 3145 10517 3179
rect 10517 3145 10551 3179
rect 10551 3145 10560 3179
rect 10508 3136 10560 3145
rect 11060 3179 11112 3188
rect 11060 3145 11069 3179
rect 11069 3145 11103 3179
rect 11103 3145 11112 3179
rect 11060 3136 11112 3145
rect 12072 3179 12124 3188
rect 12072 3145 12081 3179
rect 12081 3145 12115 3179
rect 12115 3145 12124 3179
rect 12072 3136 12124 3145
rect 15108 3136 15160 3188
rect 16948 3136 17000 3188
rect 18144 3179 18196 3188
rect 18144 3145 18153 3179
rect 18153 3145 18187 3179
rect 18187 3145 18196 3179
rect 18144 3136 18196 3145
rect 2320 3000 2372 3052
rect 5724 3068 5776 3120
rect 480 2932 532 2984
rect 6828 3000 6880 3052
rect 5724 2932 5776 2984
rect 5908 2932 5960 2984
rect 7932 2932 7984 2984
rect 8668 3068 8720 3120
rect 9496 3111 9548 3120
rect 9496 3077 9505 3111
rect 9505 3077 9539 3111
rect 9539 3077 9548 3111
rect 9496 3068 9548 3077
rect 9772 2932 9824 2984
rect 9220 2864 9272 2916
rect 6828 2796 6880 2848
rect 15568 3000 15620 3052
rect 16580 3068 16632 3120
rect 10324 2932 10376 2984
rect 12440 2932 12492 2984
rect 12624 2975 12676 2984
rect 12624 2941 12633 2975
rect 12633 2941 12667 2975
rect 12667 2941 12676 2975
rect 12624 2932 12676 2941
rect 13544 2932 13596 2984
rect 14740 2932 14792 2984
rect 16580 2932 16632 2984
rect 18420 2932 18472 2984
rect 12164 2864 12216 2916
rect 15568 2864 15620 2916
rect 11980 2796 12032 2848
rect 12808 2796 12860 2848
rect 16396 2864 16448 2916
rect 6962 2694 7014 2746
rect 7026 2694 7078 2746
rect 7090 2694 7142 2746
rect 7154 2694 7206 2746
rect 12942 2694 12994 2746
rect 13006 2694 13058 2746
rect 13070 2694 13122 2746
rect 13134 2694 13186 2746
rect 3516 2592 3568 2644
rect 4896 2592 4948 2644
rect 5908 2592 5960 2644
rect 7840 2592 7892 2644
rect 8116 2635 8168 2644
rect 8116 2601 8125 2635
rect 8125 2601 8159 2635
rect 8159 2601 8168 2635
rect 8116 2592 8168 2601
rect 9680 2592 9732 2644
rect 10324 2635 10376 2644
rect 10324 2601 10333 2635
rect 10333 2601 10367 2635
rect 10367 2601 10376 2635
rect 10324 2592 10376 2601
rect 10876 2635 10928 2644
rect 10876 2601 10885 2635
rect 10885 2601 10919 2635
rect 10919 2601 10928 2635
rect 10876 2592 10928 2601
rect 12532 2592 12584 2644
rect 14740 2592 14792 2644
rect 17316 2592 17368 2644
rect 2320 2524 2372 2576
rect 6552 2524 6604 2576
rect 3240 2456 3292 2508
rect 4620 2499 4672 2508
rect 4620 2465 4629 2499
rect 4629 2465 4663 2499
rect 4663 2465 4672 2499
rect 4620 2456 4672 2465
rect 6000 2499 6052 2508
rect 6000 2465 6009 2499
rect 6009 2465 6043 2499
rect 6043 2465 6052 2499
rect 6000 2456 6052 2465
rect 7840 2456 7892 2508
rect 8024 2499 8076 2508
rect 8024 2465 8033 2499
rect 8033 2465 8067 2499
rect 8067 2465 8076 2499
rect 8024 2456 8076 2465
rect 9772 2456 9824 2508
rect 12440 2456 12492 2508
rect 13452 2456 13504 2508
rect 13820 2456 13872 2508
rect 15200 2524 15252 2576
rect 16396 2524 16448 2576
rect 9588 2388 9640 2440
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 12716 2388 12768 2440
rect 16488 2388 16540 2440
rect 17960 2363 18012 2372
rect 17960 2329 17969 2363
rect 17969 2329 18003 2363
rect 18003 2329 18012 2363
rect 17960 2320 18012 2329
rect 3972 2150 4024 2202
rect 4036 2150 4088 2202
rect 4100 2150 4152 2202
rect 4164 2150 4216 2202
rect 9952 2150 10004 2202
rect 10016 2150 10068 2202
rect 10080 2150 10132 2202
rect 10144 2150 10196 2202
rect 15932 2150 15984 2202
rect 15996 2150 16048 2202
rect 16060 2150 16112 2202
rect 16124 2150 16176 2202
<< metal2 >>
rect 938 21540 994 22340
rect 2318 21540 2374 22340
rect 3698 21540 3754 22340
rect 5538 21540 5594 22340
rect 6918 21540 6974 22340
rect 8298 21540 8354 22340
rect 9678 21540 9734 22340
rect 11518 21540 11574 22340
rect 12898 21540 12954 22340
rect 14278 21540 14334 22340
rect 15658 21540 15714 22340
rect 17498 21540 17554 22340
rect 18878 21540 18934 22340
rect 952 19242 980 21540
rect 1490 20496 1546 20505
rect 1490 20431 1546 20440
rect 1504 20058 1532 20431
rect 1492 20052 1544 20058
rect 1492 19994 1544 20000
rect 2332 19922 2360 21540
rect 3712 19922 3740 21540
rect 5552 19922 5580 21540
rect 6932 20346 6960 21540
rect 6840 20318 6960 20346
rect 6840 19938 6868 20318
rect 6936 20156 7232 20176
rect 6992 20154 7016 20156
rect 7072 20154 7096 20156
rect 7152 20154 7176 20156
rect 7014 20102 7016 20154
rect 7078 20102 7090 20154
rect 7152 20102 7154 20154
rect 6992 20100 7016 20102
rect 7072 20100 7096 20102
rect 7152 20100 7176 20102
rect 6936 20080 7232 20100
rect 8312 19990 8340 21540
rect 7104 19984 7156 19990
rect 6840 19922 6960 19938
rect 7104 19926 7156 19932
rect 8300 19984 8352 19990
rect 8300 19926 8352 19932
rect 1584 19916 1636 19922
rect 1584 19858 1636 19864
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 2964 19916 3016 19922
rect 2964 19858 3016 19864
rect 3700 19916 3752 19922
rect 3700 19858 3752 19864
rect 5540 19916 5592 19922
rect 6840 19916 6972 19922
rect 6840 19910 6920 19916
rect 5540 19858 5592 19864
rect 6920 19858 6972 19864
rect 1596 19514 1624 19858
rect 2688 19712 2740 19718
rect 2688 19654 2740 19660
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 2412 19304 2464 19310
rect 2412 19246 2464 19252
rect 940 19236 992 19242
rect 940 19178 992 19184
rect 1398 17776 1454 17785
rect 1398 17711 1400 17720
rect 1452 17711 1454 17720
rect 1400 17682 1452 17688
rect 1872 17066 1900 19246
rect 2424 18766 2452 19246
rect 2412 18760 2464 18766
rect 2412 18702 2464 18708
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2608 17066 2636 17478
rect 1860 17060 1912 17066
rect 1860 17002 1912 17008
rect 2596 17060 2648 17066
rect 2596 17002 2648 17008
rect 1872 16114 1900 17002
rect 2700 16574 2728 19654
rect 2976 19242 3004 19858
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 2964 19236 3016 19242
rect 2964 19178 3016 19184
rect 2780 18828 2832 18834
rect 2780 18770 2832 18776
rect 2792 17746 2820 18770
rect 2780 17740 2832 17746
rect 2780 17682 2832 17688
rect 2516 16546 2728 16574
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1398 15736 1454 15745
rect 1398 15671 1454 15680
rect 1412 15570 1440 15671
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1768 15360 1820 15366
rect 1768 15302 1820 15308
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1504 13870 1532 14418
rect 1676 14000 1728 14006
rect 1676 13942 1728 13948
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1412 13705 1440 13806
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 1504 13530 1532 13806
rect 1492 13524 1544 13530
rect 1492 13466 1544 13472
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1596 11762 1624 13262
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1490 11656 1546 11665
rect 1490 11591 1546 11600
rect 1504 11354 1532 11591
rect 1492 11348 1544 11354
rect 1492 11290 1544 11296
rect 1596 9586 1624 11698
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1398 8936 1454 8945
rect 1398 8871 1400 8880
rect 1452 8871 1454 8880
rect 1400 8842 1452 8848
rect 1596 6934 1624 9522
rect 1688 9450 1716 13942
rect 1780 11762 1808 15302
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2148 11898 2176 12242
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2424 10266 2452 10542
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2516 10146 2544 16546
rect 2792 15570 2820 17682
rect 2872 15972 2924 15978
rect 2872 15914 2924 15920
rect 2884 15706 2912 15914
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 2608 13938 2636 14214
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2700 13394 2728 14418
rect 2872 14340 2924 14346
rect 2872 14282 2924 14288
rect 2884 13870 2912 14282
rect 3068 14074 3096 14418
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3068 13954 3096 14010
rect 2976 13926 3096 13954
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2700 12782 2728 13330
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2792 10470 2820 11154
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2424 10118 2544 10146
rect 1676 9444 1728 9450
rect 1676 9386 1728 9392
rect 2320 9444 2372 9450
rect 2320 9386 2372 9392
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1872 9178 1900 9318
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1964 8430 1992 9318
rect 2332 8430 2360 9386
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2332 7954 2360 8366
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2332 7342 2360 7890
rect 2424 7886 2452 10118
rect 2792 9994 2820 10406
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2884 9518 2912 13806
rect 2976 13462 3004 13926
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 2964 13456 3016 13462
rect 2964 13398 3016 13404
rect 3068 12986 3096 13806
rect 3160 13530 3188 19654
rect 3946 19612 4242 19632
rect 4002 19610 4026 19612
rect 4082 19610 4106 19612
rect 4162 19610 4186 19612
rect 4024 19558 4026 19610
rect 4088 19558 4100 19610
rect 4162 19558 4164 19610
rect 4002 19556 4026 19558
rect 4082 19556 4106 19558
rect 4162 19556 4186 19558
rect 3946 19536 4242 19556
rect 3700 19372 3752 19378
rect 3700 19314 3752 19320
rect 3332 19236 3384 19242
rect 3332 19178 3384 19184
rect 3344 18970 3372 19178
rect 3332 18964 3384 18970
rect 3332 18906 3384 18912
rect 3712 18426 3740 19314
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3988 18834 4016 19246
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4540 18834 4568 19110
rect 3976 18828 4028 18834
rect 3976 18770 4028 18776
rect 4528 18828 4580 18834
rect 4528 18770 4580 18776
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 3946 18524 4242 18544
rect 4002 18522 4026 18524
rect 4082 18522 4106 18524
rect 4162 18522 4186 18524
rect 4024 18470 4026 18522
rect 4088 18470 4100 18522
rect 4162 18470 4164 18522
rect 4002 18468 4026 18470
rect 4082 18468 4106 18470
rect 4162 18468 4186 18470
rect 3946 18448 4242 18468
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 4356 18358 4384 18566
rect 4344 18352 4396 18358
rect 4344 18294 4396 18300
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 4172 18068 4200 18226
rect 4540 18222 4568 18770
rect 4528 18216 4580 18222
rect 4528 18158 4580 18164
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 4344 18080 4396 18086
rect 4172 18040 4344 18068
rect 4344 18022 4396 18028
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 3712 17134 3740 17478
rect 3946 17436 4242 17456
rect 4002 17434 4026 17436
rect 4082 17434 4106 17436
rect 4162 17434 4186 17436
rect 4024 17382 4026 17434
rect 4088 17382 4100 17434
rect 4162 17382 4164 17434
rect 4002 17380 4026 17382
rect 4082 17380 4106 17382
rect 4162 17380 4186 17382
rect 3946 17360 4242 17380
rect 3700 17128 3752 17134
rect 3700 17070 3752 17076
rect 4068 17060 4120 17066
rect 4068 17002 4120 17008
rect 4160 17060 4212 17066
rect 4356 17048 4384 18022
rect 4540 17746 4568 18158
rect 4528 17740 4580 17746
rect 4528 17682 4580 17688
rect 4212 17020 4384 17048
rect 4160 17002 4212 17008
rect 4080 16590 4108 17002
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 3946 16348 4242 16368
rect 4002 16346 4026 16348
rect 4082 16346 4106 16348
rect 4162 16346 4186 16348
rect 4024 16294 4026 16346
rect 4088 16294 4100 16346
rect 4162 16294 4164 16346
rect 4002 16292 4026 16294
rect 4082 16292 4106 16294
rect 4162 16292 4186 16294
rect 3946 16272 4242 16292
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3528 15706 3556 15846
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 4356 15502 4384 17020
rect 4540 16998 4568 17682
rect 4632 17134 4660 18158
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4436 15904 4488 15910
rect 4436 15846 4488 15852
rect 4448 15570 4476 15846
rect 4528 15632 4580 15638
rect 4528 15574 4580 15580
rect 4436 15564 4488 15570
rect 4436 15506 4488 15512
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 3946 15260 4242 15280
rect 4002 15258 4026 15260
rect 4082 15258 4106 15260
rect 4162 15258 4186 15260
rect 4024 15206 4026 15258
rect 4088 15206 4100 15258
rect 4162 15206 4164 15258
rect 4002 15204 4026 15206
rect 4082 15204 4106 15206
rect 4162 15204 4186 15206
rect 3946 15184 4242 15204
rect 3946 14172 4242 14192
rect 4002 14170 4026 14172
rect 4082 14170 4106 14172
rect 4162 14170 4186 14172
rect 4024 14118 4026 14170
rect 4088 14118 4100 14170
rect 4162 14118 4164 14170
rect 4002 14116 4026 14118
rect 4082 14116 4106 14118
rect 4162 14116 4186 14118
rect 3946 14096 4242 14116
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 3252 13394 3280 13806
rect 3240 13388 3292 13394
rect 3240 13330 3292 13336
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3252 12918 3280 13330
rect 4356 13258 4384 15438
rect 4540 14414 4568 15574
rect 4632 15434 4660 17070
rect 4712 16108 4764 16114
rect 4816 16096 4844 19654
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 5000 17882 5028 18702
rect 4988 17876 5040 17882
rect 4988 17818 5040 17824
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5460 17338 5488 17682
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4908 16726 4936 17070
rect 4896 16720 4948 16726
rect 4896 16662 4948 16668
rect 5000 16454 5028 17138
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 5184 16794 5212 17070
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 5460 16658 5488 17070
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5080 16516 5132 16522
rect 5080 16458 5132 16464
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 4816 16068 4936 16096
rect 4712 16050 4764 16056
rect 4724 15570 4752 16050
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4620 15428 4672 15434
rect 4620 15370 4672 15376
rect 4724 14958 4752 15506
rect 4712 14952 4764 14958
rect 4712 14894 4764 14900
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4540 13870 4568 14214
rect 4528 13864 4580 13870
rect 4528 13806 4580 13812
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 3946 13084 4242 13104
rect 4002 13082 4026 13084
rect 4082 13082 4106 13084
rect 4162 13082 4186 13084
rect 4024 13030 4026 13082
rect 4088 13030 4100 13082
rect 4162 13030 4164 13082
rect 4002 13028 4026 13030
rect 4082 13028 4106 13030
rect 4162 13028 4186 13030
rect 3946 13008 4242 13028
rect 3240 12912 3292 12918
rect 3240 12854 3292 12860
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3160 12374 3188 12718
rect 3148 12368 3200 12374
rect 3148 12310 3200 12316
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 2976 11898 3004 12242
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 3068 11354 3096 11630
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 3056 10600 3108 10606
rect 3160 10588 3188 12174
rect 3946 11996 4242 12016
rect 4002 11994 4026 11996
rect 4082 11994 4106 11996
rect 4162 11994 4186 11996
rect 4024 11942 4026 11994
rect 4088 11942 4100 11994
rect 4162 11942 4164 11994
rect 4002 11940 4026 11942
rect 4082 11940 4106 11942
rect 4162 11940 4186 11942
rect 3946 11920 4242 11940
rect 4448 11898 4476 13262
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4540 12374 4568 13126
rect 4528 12368 4580 12374
rect 4528 12310 4580 12316
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4264 11354 4292 11562
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4528 11280 4580 11286
rect 4528 11222 4580 11228
rect 3946 10908 4242 10928
rect 4002 10906 4026 10908
rect 4082 10906 4106 10908
rect 4162 10906 4186 10908
rect 4024 10854 4026 10906
rect 4088 10854 4100 10906
rect 4162 10854 4164 10906
rect 4002 10852 4026 10854
rect 4082 10852 4106 10854
rect 4162 10852 4186 10854
rect 3946 10832 4242 10852
rect 3108 10560 3188 10588
rect 3056 10542 3108 10548
rect 3068 10130 3096 10542
rect 4540 10470 4568 11222
rect 4632 10810 4660 11630
rect 4724 11218 4752 14894
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4816 13326 4844 13670
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4908 11558 4936 16068
rect 5092 16046 5120 16458
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 4988 15972 5040 15978
rect 4988 15914 5040 15920
rect 5000 15162 5028 15914
rect 5092 15502 5120 15982
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5172 15564 5224 15570
rect 5172 15506 5224 15512
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 4988 15156 5040 15162
rect 4988 15098 5040 15104
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5092 14482 5120 14894
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 4988 13796 5040 13802
rect 4988 13738 5040 13744
rect 5000 13530 5028 13738
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 4988 11824 5040 11830
rect 4988 11766 5040 11772
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 5000 11336 5028 11766
rect 5092 11354 5120 14418
rect 5184 14006 5212 15506
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5276 14482 5304 15098
rect 5552 14482 5580 15574
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 5460 12782 5488 14214
rect 5552 13802 5580 14282
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5552 13394 5580 13738
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5552 12986 5580 13330
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5368 12434 5396 12718
rect 5276 12406 5396 12434
rect 5276 12102 5304 12406
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 4908 11308 5028 11336
rect 5080 11348 5132 11354
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4908 11150 4936 11308
rect 5080 11290 5132 11296
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4804 10736 4856 10742
rect 4804 10678 4856 10684
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 1584 6928 1636 6934
rect 1398 6896 1454 6905
rect 1584 6870 1636 6876
rect 1398 6831 1454 6840
rect 1412 6254 1440 6831
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1596 6458 1624 6734
rect 1780 6730 1808 7278
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 2148 7002 2176 7142
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 1768 6724 1820 6730
rect 1768 6666 1820 6672
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 2516 6390 2544 8978
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2608 8022 2636 8570
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2700 8090 2728 8366
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2596 8016 2648 8022
rect 2596 7958 2648 7964
rect 2504 6384 2556 6390
rect 2504 6326 2556 6332
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 3068 5846 3096 10066
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 3946 9820 4242 9840
rect 4002 9818 4026 9820
rect 4082 9818 4106 9820
rect 4162 9818 4186 9820
rect 4024 9766 4026 9818
rect 4088 9766 4100 9818
rect 4162 9766 4164 9818
rect 4002 9764 4026 9766
rect 4082 9764 4106 9766
rect 4162 9764 4186 9766
rect 3946 9744 4242 9764
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3344 8974 3372 9454
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3946 8732 4242 8752
rect 4002 8730 4026 8732
rect 4082 8730 4106 8732
rect 4162 8730 4186 8732
rect 4024 8678 4026 8730
rect 4088 8678 4100 8730
rect 4162 8678 4164 8730
rect 4002 8676 4026 8678
rect 4082 8676 4106 8678
rect 4162 8676 4186 8678
rect 3946 8656 4242 8676
rect 4356 8498 4384 9318
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 6866 3280 7686
rect 3332 7268 3384 7274
rect 3332 7210 3384 7216
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3344 6662 3372 7210
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3056 5840 3108 5846
rect 3056 5782 3108 5788
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3252 5166 3280 5714
rect 3344 5166 3372 6598
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 1490 4856 1546 4865
rect 1490 4791 1492 4800
rect 1544 4791 1546 4800
rect 1492 4762 1544 4768
rect 2424 4690 2452 4966
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 480 2984 532 2990
rect 480 2926 532 2932
rect 492 800 520 2926
rect 1412 2825 1440 3538
rect 2332 3058 2360 4422
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 1398 2816 1454 2825
rect 1398 2751 1454 2760
rect 2332 2582 2360 2994
rect 3528 2650 3556 8366
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4356 7886 4384 8230
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 3946 7644 4242 7664
rect 4002 7642 4026 7644
rect 4082 7642 4106 7644
rect 4162 7642 4186 7644
rect 4024 7590 4026 7642
rect 4088 7590 4100 7642
rect 4162 7590 4164 7642
rect 4002 7588 4026 7590
rect 4082 7588 4106 7590
rect 4162 7588 4186 7590
rect 3946 7568 4242 7588
rect 4356 7002 4384 7822
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 3946 6556 4242 6576
rect 4002 6554 4026 6556
rect 4082 6554 4106 6556
rect 4162 6554 4186 6556
rect 4024 6502 4026 6554
rect 4088 6502 4100 6554
rect 4162 6502 4164 6554
rect 4002 6500 4026 6502
rect 4082 6500 4106 6502
rect 4162 6500 4186 6502
rect 3946 6480 4242 6500
rect 4448 6322 4476 9862
rect 4540 8838 4568 10406
rect 4816 10198 4844 10678
rect 4804 10192 4856 10198
rect 4804 10134 4856 10140
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4540 7342 4568 8774
rect 4632 8022 4660 8774
rect 4724 8294 4752 10066
rect 4908 9518 4936 11086
rect 5092 10606 5120 11154
rect 5276 11014 5304 12038
rect 5552 11898 5580 12242
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5368 11218 5396 11834
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5092 9926 5120 10542
rect 5276 10538 5304 10950
rect 5368 10538 5396 11154
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5276 10198 5304 10474
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 5092 9674 5120 9862
rect 4988 9648 5040 9654
rect 5092 9646 5212 9674
rect 4988 9590 5040 9596
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4908 9042 4936 9454
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 5000 8974 5028 9590
rect 5184 9042 5212 9646
rect 5276 9382 5304 10134
rect 5368 10062 5396 10474
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5368 9450 5396 9998
rect 5552 9654 5580 10066
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 5000 6934 5028 8910
rect 5184 7274 5212 8978
rect 5276 8974 5304 9318
rect 5552 9042 5580 9590
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5172 7268 5224 7274
rect 5172 7210 5224 7216
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 4080 5846 4108 6122
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4448 5778 4476 6258
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 3946 5468 4242 5488
rect 4002 5466 4026 5468
rect 4082 5466 4106 5468
rect 4162 5466 4186 5468
rect 4024 5414 4026 5466
rect 4088 5414 4100 5466
rect 4162 5414 4164 5466
rect 4002 5412 4026 5414
rect 4082 5412 4106 5414
rect 4162 5412 4186 5414
rect 3946 5392 4242 5412
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 3946 4380 4242 4400
rect 4002 4378 4026 4380
rect 4082 4378 4106 4380
rect 4162 4378 4186 4380
rect 4024 4326 4026 4378
rect 4088 4326 4100 4378
rect 4162 4326 4164 4378
rect 4002 4324 4026 4326
rect 4082 4324 4106 4326
rect 4162 4324 4186 4326
rect 3946 4304 4242 4324
rect 4356 3602 4384 4558
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 3946 3292 4242 3312
rect 4002 3290 4026 3292
rect 4082 3290 4106 3292
rect 4162 3290 4186 3292
rect 4024 3238 4026 3290
rect 4088 3238 4100 3290
rect 4162 3238 4164 3290
rect 4002 3236 4026 3238
rect 4082 3236 4106 3238
rect 4162 3236 4186 3238
rect 3946 3216 4242 3236
rect 4908 2650 4936 6802
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5276 5914 5304 6054
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5184 5166 5212 5714
rect 5276 5234 5304 5850
rect 5460 5778 5488 8570
rect 5644 8498 5672 19654
rect 7116 19310 7144 19926
rect 9692 19922 9720 21540
rect 11532 19922 11560 21540
rect 12912 20346 12940 21540
rect 12820 20318 12940 20346
rect 12820 19922 12848 20318
rect 12916 20156 13212 20176
rect 12972 20154 12996 20156
rect 13052 20154 13076 20156
rect 13132 20154 13156 20156
rect 12994 20102 12996 20154
rect 13058 20102 13070 20154
rect 13132 20102 13134 20154
rect 12972 20100 12996 20102
rect 13052 20100 13076 20102
rect 13132 20100 13156 20102
rect 12916 20080 13212 20100
rect 14292 19922 14320 21540
rect 15672 19922 15700 21540
rect 16486 20496 16542 20505
rect 16486 20431 16542 20440
rect 16500 19922 16528 20431
rect 7380 19916 7432 19922
rect 7380 19858 7432 19864
rect 7840 19916 7892 19922
rect 7840 19858 7892 19864
rect 8208 19916 8260 19922
rect 8208 19858 8260 19864
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 16488 19916 16540 19922
rect 16488 19858 16540 19864
rect 7104 19304 7156 19310
rect 7156 19264 7328 19292
rect 7104 19246 7156 19252
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 5920 18902 5948 19110
rect 6012 18970 6040 19110
rect 6936 19068 7232 19088
rect 6992 19066 7016 19068
rect 7072 19066 7096 19068
rect 7152 19066 7176 19068
rect 7014 19014 7016 19066
rect 7078 19014 7090 19066
rect 7152 19014 7154 19066
rect 6992 19012 7016 19014
rect 7072 19012 7096 19014
rect 7152 19012 7176 19014
rect 6936 18992 7232 19012
rect 7300 18970 7328 19264
rect 7392 19242 7420 19858
rect 7564 19304 7616 19310
rect 7564 19246 7616 19252
rect 7380 19236 7432 19242
rect 7380 19178 7432 19184
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 6000 18964 6052 18970
rect 6000 18906 6052 18912
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 5908 18896 5960 18902
rect 5908 18838 5960 18844
rect 6552 18692 6604 18698
rect 6552 18634 6604 18640
rect 6564 17882 6592 18634
rect 7300 18290 7328 18906
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7484 18222 7512 19110
rect 7576 18698 7604 19246
rect 7852 19174 7880 19858
rect 8024 19712 8076 19718
rect 8024 19654 8076 19660
rect 8036 19378 8064 19654
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7760 18834 7788 19110
rect 7852 18970 7880 19110
rect 8220 18970 8248 19858
rect 8576 19780 8628 19786
rect 8576 19722 8628 19728
rect 10692 19780 10744 19786
rect 10692 19722 10744 19728
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7484 18086 7512 18158
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 6840 17882 6868 18022
rect 6936 17980 7232 18000
rect 6992 17978 7016 17980
rect 7072 17978 7096 17980
rect 7152 17978 7176 17980
rect 7014 17926 7016 17978
rect 7078 17926 7090 17978
rect 7152 17926 7154 17978
rect 6992 17924 7016 17926
rect 7072 17924 7096 17926
rect 7152 17924 7176 17926
rect 6936 17904 7232 17924
rect 6552 17876 6604 17882
rect 6552 17818 6604 17824
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5736 16046 5764 16390
rect 5828 16250 5856 16730
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5724 15564 5776 15570
rect 5724 15506 5776 15512
rect 5736 15162 5764 15506
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5736 14482 5764 15098
rect 5828 15026 5856 16186
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5828 14890 5856 14962
rect 5816 14884 5868 14890
rect 5816 14826 5868 14832
rect 5828 14498 5856 14826
rect 5724 14476 5776 14482
rect 5828 14470 5948 14498
rect 5724 14418 5776 14424
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5736 12782 5764 13262
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5736 12238 5764 12718
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5460 5302 5488 5714
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 5184 4690 5212 5102
rect 5644 4826 5672 5646
rect 5736 5574 5764 11018
rect 5828 10810 5856 14350
rect 5920 12986 5948 14470
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 5908 12164 5960 12170
rect 5908 12106 5960 12112
rect 5920 11762 5948 12106
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5828 9110 5856 10746
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 6012 7342 6040 17478
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 6380 16590 6408 16934
rect 6564 16590 6592 17818
rect 7484 17134 7512 18022
rect 7668 17678 7696 18566
rect 7760 18170 7788 18770
rect 7852 18290 7880 18906
rect 8220 18834 8248 18906
rect 8024 18828 8076 18834
rect 7944 18788 8024 18816
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7944 18222 7972 18788
rect 8024 18770 8076 18776
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 7932 18216 7984 18222
rect 7760 18154 7880 18170
rect 7932 18158 7984 18164
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 7760 18148 7892 18154
rect 7760 18142 7840 18148
rect 7840 18090 7892 18096
rect 7944 17882 7972 18158
rect 7932 17876 7984 17882
rect 7932 17818 7984 17824
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 8496 17134 8524 18158
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 6936 16892 7232 16912
rect 6992 16890 7016 16892
rect 7072 16890 7096 16892
rect 7152 16890 7176 16892
rect 7014 16838 7016 16890
rect 7078 16838 7090 16890
rect 7152 16838 7154 16890
rect 6992 16836 7016 16838
rect 7072 16836 7096 16838
rect 7152 16836 7176 16838
rect 6936 16816 7232 16836
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6288 11286 6316 12174
rect 6564 11762 6592 16526
rect 6840 16046 6868 16730
rect 7576 16726 7604 16934
rect 7564 16720 7616 16726
rect 7564 16662 7616 16668
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 6932 16250 6960 16526
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6840 14958 6868 15982
rect 7208 15978 7328 15994
rect 7196 15972 7328 15978
rect 7248 15966 7328 15972
rect 7196 15914 7248 15920
rect 6936 15804 7232 15824
rect 6992 15802 7016 15804
rect 7072 15802 7096 15804
rect 7152 15802 7176 15804
rect 7014 15750 7016 15802
rect 7078 15750 7090 15802
rect 7152 15750 7154 15802
rect 6992 15748 7016 15750
rect 7072 15748 7096 15750
rect 7152 15748 7176 15750
rect 6936 15728 7232 15748
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6840 14414 6868 14894
rect 7300 14822 7328 15966
rect 7564 15904 7616 15910
rect 7564 15846 7616 15852
rect 7576 15706 7604 15846
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7668 15162 7696 15506
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7472 14884 7524 14890
rect 7472 14826 7524 14832
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 6936 14716 7232 14736
rect 6992 14714 7016 14716
rect 7072 14714 7096 14716
rect 7152 14714 7176 14716
rect 7014 14662 7016 14714
rect 7078 14662 7090 14714
rect 7152 14662 7154 14714
rect 6992 14660 7016 14662
rect 7072 14660 7096 14662
rect 7152 14660 7176 14662
rect 6936 14640 7232 14660
rect 7300 14414 7328 14758
rect 7484 14482 7512 14826
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 7116 13870 7144 14214
rect 7484 14074 7512 14418
rect 7656 14340 7708 14346
rect 7656 14282 7708 14288
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 13326 6868 13670
rect 6936 13628 7232 13648
rect 6992 13626 7016 13628
rect 7072 13626 7096 13628
rect 7152 13626 7176 13628
rect 7014 13574 7016 13626
rect 7078 13574 7090 13626
rect 7152 13574 7154 13626
rect 6992 13572 7016 13574
rect 7072 13572 7096 13574
rect 7152 13572 7176 13574
rect 6936 13552 7232 13572
rect 7576 13530 7604 13806
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 6936 12540 7232 12560
rect 6992 12538 7016 12540
rect 7072 12538 7096 12540
rect 7152 12538 7176 12540
rect 7014 12486 7016 12538
rect 7078 12486 7090 12538
rect 7152 12486 7154 12538
rect 6992 12484 7016 12486
rect 7072 12484 7096 12486
rect 7152 12484 7176 12486
rect 6936 12464 7232 12484
rect 7300 12434 7328 13194
rect 7484 12782 7512 13330
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7208 12406 7328 12434
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6932 11898 6960 12242
rect 7208 11898 7236 12406
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7300 11778 7328 11834
rect 6552 11756 6604 11762
rect 7300 11750 7420 11778
rect 6552 11698 6604 11704
rect 7392 11626 7420 11750
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 6936 11452 7232 11472
rect 6992 11450 7016 11452
rect 7072 11450 7096 11452
rect 7152 11450 7176 11452
rect 7014 11398 7016 11450
rect 7078 11398 7090 11450
rect 7152 11398 7154 11450
rect 6992 11396 7016 11398
rect 7072 11396 7096 11398
rect 7152 11396 7176 11398
rect 6936 11376 7232 11396
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6288 10130 6316 11222
rect 7392 11218 7420 11562
rect 7484 11354 7512 12718
rect 7576 12238 7604 12922
rect 7668 12782 7696 14282
rect 7760 14260 7788 17070
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7852 15978 7880 16390
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 7840 15972 7892 15978
rect 7840 15914 7892 15920
rect 7852 14890 7880 15914
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 7944 14890 7972 15438
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 7840 14884 7892 14890
rect 7840 14826 7892 14832
rect 7932 14884 7984 14890
rect 7932 14826 7984 14832
rect 7852 14362 7880 14826
rect 7944 14482 7972 14826
rect 8128 14482 8156 14894
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 7852 14334 7972 14362
rect 7760 14232 7880 14260
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7760 13394 7788 13874
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7852 13190 7880 14232
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7668 12374 7696 12718
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7668 11626 7696 12038
rect 7852 11898 7880 12718
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7944 11778 7972 14334
rect 8024 14340 8076 14346
rect 8024 14282 8076 14288
rect 8036 13870 8064 14282
rect 8220 14074 8248 16050
rect 8312 16046 8340 17002
rect 8588 16250 8616 19722
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 9926 19612 10222 19632
rect 9982 19610 10006 19612
rect 10062 19610 10086 19612
rect 10142 19610 10166 19612
rect 10004 19558 10006 19610
rect 10068 19558 10080 19610
rect 10142 19558 10144 19610
rect 9982 19556 10006 19558
rect 10062 19556 10086 19558
rect 10142 19556 10166 19558
rect 9926 19536 10222 19556
rect 9036 19236 9088 19242
rect 9036 19178 9088 19184
rect 9680 19236 9732 19242
rect 9680 19178 9732 19184
rect 9048 18426 9076 19178
rect 9692 18834 9720 19178
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9926 18524 10222 18544
rect 9982 18522 10006 18524
rect 10062 18522 10086 18524
rect 10142 18522 10166 18524
rect 10004 18470 10006 18522
rect 10068 18470 10080 18522
rect 10142 18470 10144 18522
rect 9982 18468 10006 18470
rect 10062 18468 10086 18470
rect 10142 18468 10166 18470
rect 9926 18448 10222 18468
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9692 17202 9720 17614
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9784 16658 9812 17478
rect 9926 17436 10222 17456
rect 9982 17434 10006 17436
rect 10062 17434 10086 17436
rect 10142 17434 10166 17436
rect 10004 17382 10006 17434
rect 10068 17382 10080 17434
rect 10142 17382 10144 17434
rect 9982 17380 10006 17382
rect 10062 17380 10086 17382
rect 10142 17380 10166 17382
rect 9926 17360 10222 17380
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9876 16538 9904 17138
rect 9784 16510 9904 16538
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 8588 16046 8616 16186
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 8036 12986 8064 13806
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 7852 11762 7972 11778
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7840 11756 7972 11762
rect 7892 11750 7972 11756
rect 7840 11698 7892 11704
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7208 11082 7236 11154
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 6936 10364 7232 10384
rect 6992 10362 7016 10364
rect 7072 10362 7096 10364
rect 7152 10362 7176 10364
rect 7014 10310 7016 10362
rect 7078 10310 7090 10362
rect 7152 10310 7154 10362
rect 6992 10308 7016 10310
rect 7072 10308 7096 10310
rect 7152 10308 7176 10310
rect 6936 10288 7232 10308
rect 7300 10146 7328 10950
rect 7392 10606 7420 11154
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7208 10130 7328 10146
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 7196 10124 7328 10130
rect 7248 10118 7328 10124
rect 7196 10066 7248 10072
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6656 9518 6684 9998
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6656 8974 6684 9454
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6552 8900 6604 8906
rect 6552 8842 6604 8848
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5736 3652 5764 5510
rect 5816 3664 5868 3670
rect 5736 3624 5816 3652
rect 5736 3126 5764 3624
rect 5816 3606 5868 3612
rect 5724 3120 5776 3126
rect 5724 3062 5776 3068
rect 5736 2990 5764 3062
rect 5920 2990 5948 7210
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 5920 2650 5948 2926
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 6564 2582 6592 8842
rect 6840 7206 6868 9862
rect 7300 9654 7328 10118
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7288 9512 7340 9518
rect 7392 9500 7420 10542
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7340 9472 7420 9500
rect 7288 9454 7340 9460
rect 6936 9276 7232 9296
rect 6992 9274 7016 9276
rect 7072 9274 7096 9276
rect 7152 9274 7176 9276
rect 7014 9222 7016 9274
rect 7078 9222 7090 9274
rect 7152 9222 7154 9274
rect 6992 9220 7016 9222
rect 7072 9220 7096 9222
rect 7152 9220 7176 9222
rect 6936 9200 7232 9220
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 6936 8188 7232 8208
rect 6992 8186 7016 8188
rect 7072 8186 7096 8188
rect 7152 8186 7176 8188
rect 7014 8134 7016 8186
rect 7078 8134 7090 8186
rect 7152 8134 7154 8186
rect 6992 8132 7016 8134
rect 7072 8132 7096 8134
rect 7152 8132 7176 8134
rect 6936 8112 7232 8132
rect 7300 7954 7328 8230
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6656 5914 6684 6190
rect 6840 5914 6868 7142
rect 6936 7100 7232 7120
rect 6992 7098 7016 7100
rect 7072 7098 7096 7100
rect 7152 7098 7176 7100
rect 7014 7046 7016 7098
rect 7078 7046 7090 7098
rect 7152 7046 7154 7098
rect 6992 7044 7016 7046
rect 7072 7044 7096 7046
rect 7152 7044 7176 7046
rect 6936 7024 7232 7044
rect 7392 6866 7420 7278
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 6936 6012 7232 6032
rect 6992 6010 7016 6012
rect 7072 6010 7096 6012
rect 7152 6010 7176 6012
rect 7014 5958 7016 6010
rect 7078 5958 7090 6010
rect 7152 5958 7154 6010
rect 6992 5956 7016 5958
rect 7072 5956 7096 5958
rect 7152 5956 7176 5958
rect 6936 5936 7232 5956
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6656 5166 6684 5850
rect 7392 5166 7420 6802
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 6936 4924 7232 4944
rect 6992 4922 7016 4924
rect 7072 4922 7096 4924
rect 7152 4922 7176 4924
rect 7014 4870 7016 4922
rect 7078 4870 7090 4922
rect 7152 4870 7154 4922
rect 6992 4868 7016 4870
rect 7072 4868 7096 4870
rect 7152 4868 7176 4870
rect 6936 4848 7232 4868
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 6936 3836 7232 3856
rect 6992 3834 7016 3836
rect 7072 3834 7096 3836
rect 7152 3834 7176 3836
rect 7014 3782 7016 3834
rect 7078 3782 7090 3834
rect 7152 3782 7154 3834
rect 6992 3780 7016 3782
rect 7072 3780 7096 3782
rect 7152 3780 7176 3782
rect 6936 3760 7232 3780
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6840 3058 6868 3674
rect 7300 3670 7328 4558
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7392 4146 7420 4422
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7484 4078 7512 9862
rect 7576 9722 7604 9998
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7576 9042 7604 9658
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7576 7342 7604 8434
rect 7760 8022 7788 11698
rect 7944 11082 7972 11750
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7944 10810 7972 11018
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 8036 10690 8064 12242
rect 8128 11014 8156 14010
rect 8220 13326 8248 14010
rect 8312 13938 8340 15982
rect 9416 15502 9444 15982
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9508 15366 9536 16050
rect 9600 16046 9628 16186
rect 9784 16096 9812 16510
rect 9926 16348 10222 16368
rect 9982 16346 10006 16348
rect 10062 16346 10086 16348
rect 10142 16346 10166 16348
rect 10004 16294 10006 16346
rect 10068 16294 10080 16346
rect 10142 16294 10144 16346
rect 9982 16292 10006 16294
rect 10062 16292 10086 16294
rect 10142 16292 10166 16294
rect 9926 16272 10222 16292
rect 9864 16108 9916 16114
rect 9784 16068 9864 16096
rect 9864 16050 9916 16056
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10244 15638 10272 15982
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9692 15162 9720 15506
rect 9926 15260 10222 15280
rect 9982 15258 10006 15260
rect 10062 15258 10086 15260
rect 10142 15258 10166 15260
rect 10004 15206 10006 15258
rect 10068 15206 10080 15258
rect 10142 15206 10144 15258
rect 9982 15204 10006 15206
rect 10062 15204 10086 15206
rect 10142 15204 10166 15206
rect 9926 15184 10222 15204
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 8220 12442 8248 13126
rect 8208 12436 8260 12442
rect 8404 12434 8432 14214
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9140 13530 9168 13806
rect 9232 13802 9260 14418
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9324 13870 9352 14214
rect 9926 14172 10222 14192
rect 9982 14170 10006 14172
rect 10062 14170 10086 14172
rect 10142 14170 10166 14172
rect 10004 14118 10006 14170
rect 10068 14118 10080 14170
rect 10142 14118 10144 14170
rect 9982 14116 10006 14118
rect 10062 14116 10086 14118
rect 10142 14116 10166 14118
rect 9926 14096 10222 14116
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9508 13394 9536 13806
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 10060 13462 10088 13670
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 8208 12378 8260 12384
rect 8312 12406 8432 12434
rect 9508 12434 9536 13330
rect 9926 13084 10222 13104
rect 9982 13082 10006 13084
rect 10062 13082 10086 13084
rect 10142 13082 10166 13084
rect 10004 13030 10006 13082
rect 10068 13030 10080 13082
rect 10142 13030 10144 13082
rect 9982 13028 10006 13030
rect 10062 13028 10086 13030
rect 10142 13028 10166 13030
rect 9926 13008 10222 13028
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9508 12406 9628 12434
rect 8220 12306 8248 12378
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8312 12102 8340 12406
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 7944 10662 8064 10690
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7576 7002 7604 7278
rect 7944 7206 7972 10662
rect 8128 10606 8156 10950
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8128 9024 8156 9998
rect 8220 9586 8248 11154
rect 8312 10130 8340 12038
rect 8496 11830 8524 12106
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8484 10600 8536 10606
rect 8404 10560 8484 10588
rect 8404 10130 8432 10560
rect 8484 10542 8536 10548
rect 8772 10470 8800 12242
rect 9416 12102 9444 12242
rect 9600 12170 9628 12406
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9416 11762 9444 12038
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9140 11286 9168 11630
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 9140 10606 9168 11222
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8404 9518 8432 10066
rect 8772 9738 8800 10406
rect 9048 10130 9076 10474
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 8772 9710 8984 9738
rect 8956 9518 8984 9710
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8208 9036 8260 9042
rect 8128 8996 8208 9024
rect 8208 8978 8260 8984
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7576 5710 7604 6938
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7576 4214 7604 5646
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7944 4826 7972 4966
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7668 4282 7696 4558
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 7564 4208 7616 4214
rect 7564 4150 7616 4156
rect 7668 4078 7696 4218
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7288 3664 7340 3670
rect 7288 3606 7340 3612
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6840 2854 6868 2994
rect 7944 2990 7972 3470
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 7944 2774 7972 2926
rect 6936 2748 7232 2768
rect 6992 2746 7016 2748
rect 7072 2746 7096 2748
rect 7152 2746 7176 2748
rect 7014 2694 7016 2746
rect 7078 2694 7090 2746
rect 7152 2694 7154 2746
rect 6992 2692 7016 2694
rect 7072 2692 7096 2694
rect 7152 2692 7176 2694
rect 6936 2672 7232 2692
rect 7852 2746 7972 2774
rect 7852 2650 7880 2746
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 2320 2576 2372 2582
rect 2320 2518 2372 2524
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 8036 2514 8064 8774
rect 8220 8362 8248 8978
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8128 6866 8156 8230
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 8128 5778 8156 6802
rect 8312 6798 8340 8366
rect 8496 8294 8524 9318
rect 8680 9110 8708 9454
rect 9324 9110 9352 11086
rect 9416 10674 9444 11698
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9508 10554 9536 11766
rect 9692 11150 9720 12106
rect 9784 11898 9812 12786
rect 9926 11996 10222 12016
rect 9982 11994 10006 11996
rect 10062 11994 10086 11996
rect 10142 11994 10166 11996
rect 10004 11942 10006 11994
rect 10068 11942 10080 11994
rect 10142 11942 10144 11994
rect 9982 11940 10006 11942
rect 10062 11940 10086 11942
rect 10142 11940 10166 11942
rect 9926 11920 10222 11940
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 10336 11778 10364 19654
rect 10600 19168 10652 19174
rect 10600 19110 10652 19116
rect 10612 18902 10640 19110
rect 10600 18896 10652 18902
rect 10600 18838 10652 18844
rect 10416 17536 10468 17542
rect 10416 17478 10468 17484
rect 10428 17202 10456 17478
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 10428 16726 10456 17138
rect 10416 16720 10468 16726
rect 10416 16662 10468 16668
rect 10508 16652 10560 16658
rect 10508 16594 10560 16600
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10428 15026 10456 16526
rect 10520 15706 10548 16594
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10428 12238 10456 13262
rect 10704 12646 10732 19722
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 16488 19712 16540 19718
rect 16488 19654 16540 19660
rect 10784 17128 10836 17134
rect 10782 17096 10784 17105
rect 10836 17096 10838 17105
rect 10782 17031 10838 17040
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10796 16658 10824 16934
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10888 14618 10916 14894
rect 10968 14884 11020 14890
rect 10968 14826 11020 14832
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10796 12102 10824 13806
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10336 11750 10456 11778
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9926 10908 10222 10928
rect 9982 10906 10006 10908
rect 10062 10906 10086 10908
rect 10142 10906 10166 10908
rect 10004 10854 10006 10906
rect 10068 10854 10080 10906
rect 10142 10854 10144 10906
rect 9982 10852 10006 10854
rect 10062 10852 10086 10854
rect 10142 10852 10166 10854
rect 9926 10832 10222 10852
rect 9416 10526 9536 10554
rect 10336 10538 10364 11630
rect 10324 10532 10376 10538
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 9312 9104 9364 9110
rect 9312 9046 9364 9052
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8772 7342 8800 8434
rect 9324 7954 9352 9046
rect 9416 8430 9444 10526
rect 10324 10474 10376 10480
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9508 10062 9536 10406
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9508 8974 9536 9318
rect 9600 9178 9628 10066
rect 9926 9820 10222 9840
rect 9982 9818 10006 9820
rect 10062 9818 10086 9820
rect 10142 9818 10166 9820
rect 10004 9766 10006 9818
rect 10068 9766 10080 9818
rect 10142 9766 10144 9818
rect 9982 9764 10006 9766
rect 10062 9764 10086 9766
rect 10142 9764 10166 9766
rect 9926 9744 10222 9764
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9508 7750 9536 8910
rect 9600 8906 9628 9114
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9600 8634 9628 8842
rect 9692 8838 9720 9386
rect 10336 8838 10364 10474
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9692 7954 9720 8774
rect 9926 8732 10222 8752
rect 9982 8730 10006 8732
rect 10062 8730 10086 8732
rect 10142 8730 10166 8732
rect 10004 8678 10006 8730
rect 10068 8678 10080 8730
rect 10142 8678 10144 8730
rect 9982 8676 10006 8678
rect 10062 8676 10086 8678
rect 10142 8676 10166 8678
rect 9926 8656 10222 8676
rect 10428 8362 10456 11750
rect 10796 11694 10824 12038
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10612 11354 10640 11630
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10704 9450 10732 10474
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 9128 7268 9180 7274
rect 9128 7210 9180 7216
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8588 6662 8616 7142
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8404 5302 8432 6190
rect 8588 5914 8616 6598
rect 8772 6322 8800 7142
rect 9140 6798 9168 7210
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 9140 6254 9168 6734
rect 9324 6254 9352 6802
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 9324 5778 9352 6190
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8128 2650 8156 3334
rect 8404 3194 8432 3674
rect 8680 3602 8708 4014
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8680 3126 8708 3538
rect 9508 3126 9536 6054
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 8668 3120 8720 3126
rect 8668 3062 8720 3068
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 9220 2916 9272 2922
rect 9220 2858 9272 2864
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 1872 800 1900 2314
rect 3252 800 3280 2450
rect 3946 2204 4242 2224
rect 4002 2202 4026 2204
rect 4082 2202 4106 2204
rect 4162 2202 4186 2204
rect 4024 2150 4026 2202
rect 4088 2150 4100 2202
rect 4162 2150 4164 2202
rect 4002 2148 4026 2150
rect 4082 2148 4106 2150
rect 4162 2148 4186 2150
rect 3946 2128 4242 2148
rect 4632 800 4660 2450
rect 6012 800 6040 2450
rect 7852 800 7880 2450
rect 9232 800 9260 2858
rect 9600 2446 9628 4150
rect 9692 2650 9720 7686
rect 9784 6866 9812 7754
rect 9926 7644 10222 7664
rect 9982 7642 10006 7644
rect 10062 7642 10086 7644
rect 10142 7642 10166 7644
rect 10004 7590 10006 7642
rect 10068 7590 10080 7642
rect 10142 7590 10144 7642
rect 9982 7588 10006 7590
rect 10062 7588 10086 7590
rect 10142 7588 10166 7590
rect 9926 7568 10222 7588
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9784 6254 9812 6802
rect 9926 6556 10222 6576
rect 9982 6554 10006 6556
rect 10062 6554 10086 6556
rect 10142 6554 10166 6556
rect 10004 6502 10006 6554
rect 10068 6502 10080 6554
rect 10142 6502 10144 6554
rect 9982 6500 10006 6502
rect 10062 6500 10086 6502
rect 10142 6500 10166 6502
rect 9926 6480 10222 6500
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 10704 5794 10732 8774
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10796 5914 10824 6190
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10508 5772 10560 5778
rect 10704 5766 10824 5794
rect 10508 5714 10560 5720
rect 9926 5468 10222 5488
rect 9982 5466 10006 5468
rect 10062 5466 10086 5468
rect 10142 5466 10166 5468
rect 10004 5414 10006 5466
rect 10068 5414 10080 5466
rect 10142 5414 10144 5466
rect 9982 5412 10006 5414
rect 10062 5412 10086 5414
rect 10142 5412 10166 5414
rect 9926 5392 10222 5412
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9784 4690 9812 5102
rect 10520 5030 10548 5714
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10520 4758 10548 4966
rect 10508 4752 10560 4758
rect 10508 4694 10560 4700
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9784 4282 9812 4626
rect 9926 4380 10222 4400
rect 9982 4378 10006 4380
rect 10062 4378 10086 4380
rect 10142 4378 10166 4380
rect 10004 4326 10006 4378
rect 10068 4326 10080 4378
rect 10142 4326 10144 4378
rect 9982 4324 10006 4326
rect 10062 4324 10086 4326
rect 10142 4324 10166 4326
rect 9926 4304 10222 4324
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 10324 4140 10376 4146
rect 10376 4100 10640 4128
rect 10324 4082 10376 4088
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 9926 3292 10222 3312
rect 9982 3290 10006 3292
rect 10062 3290 10086 3292
rect 10142 3290 10166 3292
rect 10004 3238 10006 3290
rect 10068 3238 10080 3290
rect 10142 3238 10144 3290
rect 9982 3236 10006 3238
rect 10062 3236 10086 3238
rect 10142 3236 10166 3238
rect 9926 3216 10222 3236
rect 10336 2990 10364 3470
rect 10520 3194 10548 3606
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 10324 2984 10376 2990
rect 10324 2926 10376 2932
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9784 2514 9812 2926
rect 10336 2650 10364 2926
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9926 2204 10222 2224
rect 9982 2202 10006 2204
rect 10062 2202 10086 2204
rect 10142 2202 10166 2204
rect 10004 2150 10006 2202
rect 10068 2150 10080 2202
rect 10142 2150 10144 2202
rect 9982 2148 10006 2150
rect 10062 2148 10086 2150
rect 10142 2148 10166 2150
rect 9926 2128 10222 2148
rect 10612 800 10640 4100
rect 10704 3602 10732 5034
rect 10796 3942 10824 5766
rect 10888 5166 10916 6802
rect 10876 5160 10928 5166
rect 10876 5102 10928 5108
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10980 2774 11008 14826
rect 11072 14482 11100 15302
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 11164 14074 11192 15982
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11072 12170 11100 13126
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 11164 11694 11192 12242
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 11072 10810 11100 11222
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11164 10674 11192 11494
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11164 10198 11192 10610
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11256 9178 11284 19654
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12176 18630 12204 18770
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 11704 18352 11756 18358
rect 11704 18294 11756 18300
rect 11716 17678 11744 18294
rect 12176 18290 12204 18566
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12164 18148 12216 18154
rect 12164 18090 12216 18096
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11808 17746 11836 18022
rect 12176 17746 12204 18090
rect 11796 17740 11848 17746
rect 12164 17740 12216 17746
rect 11796 17682 11848 17688
rect 12084 17700 12164 17728
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11992 15706 12020 15846
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 11992 15366 12020 15642
rect 12084 15434 12112 17700
rect 12164 17682 12216 17688
rect 12360 17134 12388 18702
rect 12452 18426 12480 18770
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12360 16810 12388 17070
rect 12452 16946 12480 18362
rect 12544 17524 12572 18702
rect 12624 18080 12676 18086
rect 12624 18022 12676 18028
rect 12636 17882 12664 18022
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12728 17678 12756 19654
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12820 18766 12848 19246
rect 13820 19236 13872 19242
rect 13820 19178 13872 19184
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 12916 19068 13212 19088
rect 12972 19066 12996 19068
rect 13052 19066 13076 19068
rect 13132 19066 13156 19068
rect 12994 19014 12996 19066
rect 13058 19014 13070 19066
rect 13132 19014 13134 19066
rect 12972 19012 12996 19014
rect 13052 19012 13076 19014
rect 13132 19012 13156 19014
rect 12916 18992 13212 19012
rect 13176 18828 13228 18834
rect 13176 18770 13228 18776
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 13188 18426 13216 18770
rect 13280 18698 13308 19110
rect 13464 18970 13492 19110
rect 13832 18970 13860 19178
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13268 18692 13320 18698
rect 13268 18634 13320 18640
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13464 18154 13492 18906
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13556 18154 13584 18838
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 13452 18148 13504 18154
rect 13452 18090 13504 18096
rect 13544 18148 13596 18154
rect 13544 18090 13596 18096
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12820 17814 12848 18022
rect 12916 17980 13212 18000
rect 12972 17978 12996 17980
rect 13052 17978 13076 17980
rect 13132 17978 13156 17980
rect 12994 17926 12996 17978
rect 13058 17926 13070 17978
rect 13132 17926 13134 17978
rect 12972 17924 12996 17926
rect 13052 17924 13076 17926
rect 13132 17924 13156 17926
rect 12916 17904 13212 17924
rect 12808 17808 12860 17814
rect 12808 17750 12860 17756
rect 13464 17746 13492 18090
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12544 17496 12848 17524
rect 12820 17202 12848 17496
rect 13464 17270 13492 17682
rect 13556 17610 13584 18090
rect 14200 17678 14228 18158
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 13544 17604 13596 17610
rect 13544 17546 13596 17552
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12452 16918 12572 16946
rect 12360 16782 12480 16810
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12176 16046 12204 16526
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 12164 16040 12216 16046
rect 12164 15982 12216 15988
rect 12176 15570 12204 15982
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 12268 15502 12296 16390
rect 12360 15978 12388 16594
rect 12452 16046 12480 16782
rect 12544 16114 12572 16918
rect 12728 16726 12756 17070
rect 12820 16794 12848 17138
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13544 17128 13596 17134
rect 13544 17070 13596 17076
rect 12916 16892 13212 16912
rect 12972 16890 12996 16892
rect 13052 16890 13076 16892
rect 13132 16890 13156 16892
rect 12994 16838 12996 16890
rect 13058 16838 13070 16890
rect 13132 16838 13134 16890
rect 12972 16836 12996 16838
rect 13052 16836 13076 16838
rect 13132 16836 13156 16838
rect 12916 16816 13212 16836
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 13372 16658 13400 17070
rect 13556 16794 13584 17070
rect 14200 16794 14228 17614
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 14200 16522 14228 16730
rect 14188 16516 14240 16522
rect 14188 16458 14240 16464
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 12348 15972 12400 15978
rect 12348 15914 12400 15920
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 12916 15804 13212 15824
rect 12972 15802 12996 15804
rect 13052 15802 13076 15804
rect 13132 15802 13156 15804
rect 12994 15750 12996 15802
rect 13058 15750 13070 15802
rect 13132 15750 13134 15802
rect 12972 15748 12996 15750
rect 13052 15748 13076 15750
rect 13132 15748 13156 15750
rect 12916 15728 13212 15748
rect 13464 15638 13492 15846
rect 13452 15632 13504 15638
rect 13452 15574 13504 15580
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11992 15026 12020 15302
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 12268 14958 12296 15438
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11532 14618 11560 14758
rect 12916 14716 13212 14736
rect 12972 14714 12996 14716
rect 13052 14714 13076 14716
rect 13132 14714 13156 14716
rect 12994 14662 12996 14714
rect 13058 14662 13070 14714
rect 13132 14662 13134 14714
rect 12972 14660 12996 14662
rect 13052 14660 13076 14662
rect 13132 14660 13156 14662
rect 12916 14640 13212 14660
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11532 14482 11560 14554
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11716 13530 11744 14350
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 12916 13628 13212 13648
rect 12972 13626 12996 13628
rect 13052 13626 13076 13628
rect 13132 13626 13156 13628
rect 12994 13574 12996 13626
rect 13058 13574 13070 13626
rect 13132 13574 13134 13626
rect 12972 13572 12996 13574
rect 13052 13572 13076 13574
rect 13132 13572 13156 13574
rect 12916 13552 13212 13572
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11428 13456 11480 13462
rect 11428 13398 11480 13404
rect 11440 12442 11468 13398
rect 13280 13394 13308 14214
rect 13372 13938 13400 14418
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13556 12918 13584 15982
rect 14004 15972 14056 15978
rect 14004 15914 14056 15920
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 13740 13530 13768 13738
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13740 13326 13768 13466
rect 13832 13394 13860 13670
rect 13924 13462 13952 13806
rect 14016 13734 14044 15914
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 13912 13456 13964 13462
rect 13912 13398 13964 13404
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13544 12912 13596 12918
rect 13544 12854 13596 12860
rect 13556 12782 13584 12854
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13832 12714 13860 13330
rect 13924 12850 13952 13398
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 13820 12708 13872 12714
rect 13820 12650 13872 12656
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11336 11620 11388 11626
rect 11336 11562 11388 11568
rect 11348 11354 11376 11562
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11532 11218 11560 12650
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12452 12374 12480 12582
rect 12916 12540 13212 12560
rect 12972 12538 12996 12540
rect 13052 12538 13076 12540
rect 13132 12538 13156 12540
rect 12994 12486 12996 12538
rect 13058 12486 13070 12538
rect 13132 12486 13134 12538
rect 12972 12484 12996 12486
rect 13052 12484 13076 12486
rect 13132 12484 13156 12486
rect 12916 12464 13212 12484
rect 13924 12442 13952 12786
rect 14016 12646 14044 13670
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 12440 12368 12492 12374
rect 12440 12310 12492 12316
rect 13360 12368 13412 12374
rect 14108 12322 14136 15642
rect 14200 15502 14228 16458
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 13360 12310 13412 12316
rect 13372 11898 13400 12310
rect 14016 12306 14136 12322
rect 14004 12300 14136 12306
rect 14056 12294 14136 12300
rect 14004 12242 14056 12248
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 14016 11694 14044 12242
rect 14200 12238 14228 15438
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 14200 11694 14228 12174
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 12916 11452 13212 11472
rect 12972 11450 12996 11452
rect 13052 11450 13076 11452
rect 13132 11450 13156 11452
rect 12994 11398 12996 11450
rect 13058 11398 13070 11450
rect 13132 11398 13134 11450
rect 12972 11396 12996 11398
rect 13052 11396 13076 11398
rect 13132 11396 13156 11398
rect 12916 11376 13212 11396
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 11440 10810 11468 11154
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11532 10674 11560 10950
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11716 10062 11744 11086
rect 12268 10130 12296 11154
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11716 8974 11744 9998
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11716 7324 11744 8910
rect 11808 8430 11836 8978
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 11808 7954 11836 8366
rect 12084 8090 12112 8366
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12268 8022 12296 10066
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11808 7478 11836 7890
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 11796 7472 11848 7478
rect 11796 7414 11848 7420
rect 11716 7296 11836 7324
rect 11808 6798 11836 7296
rect 12084 7002 12112 7686
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11532 4690 11560 5102
rect 11808 4690 11836 6734
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12360 6254 12388 6598
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12360 5778 12388 6190
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11532 3738 11560 4626
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11624 4214 11652 4558
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 12452 4078 12480 8502
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 12544 3670 12572 9998
rect 12636 7954 12664 11290
rect 14200 11150 14228 11630
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12820 10606 12848 10950
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 12916 10364 13212 10384
rect 12972 10362 12996 10364
rect 13052 10362 13076 10364
rect 13132 10362 13156 10364
rect 12994 10310 12996 10362
rect 13058 10310 13070 10362
rect 13132 10310 13134 10362
rect 12972 10308 12996 10310
rect 13052 10308 13076 10310
rect 13132 10308 13156 10310
rect 12916 10288 13212 10308
rect 13280 9586 13308 10406
rect 13464 10198 13492 10406
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 13556 10130 13584 10610
rect 14384 10606 14412 19654
rect 14924 19304 14976 19310
rect 14924 19246 14976 19252
rect 14936 18902 14964 19246
rect 15304 18902 15332 19654
rect 15906 19612 16202 19632
rect 15962 19610 15986 19612
rect 16042 19610 16066 19612
rect 16122 19610 16146 19612
rect 15984 19558 15986 19610
rect 16048 19558 16060 19610
rect 16122 19558 16124 19610
rect 15962 19556 15986 19558
rect 16042 19556 16066 19558
rect 16122 19556 16146 19558
rect 15906 19536 16202 19556
rect 15752 19236 15804 19242
rect 15752 19178 15804 19184
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15488 18902 15516 19110
rect 14924 18896 14976 18902
rect 14924 18838 14976 18844
rect 15292 18896 15344 18902
rect 15292 18838 15344 18844
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14660 18222 14688 18702
rect 14648 18216 14700 18222
rect 14648 18158 14700 18164
rect 14936 17746 14964 18838
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14476 16590 14504 17138
rect 14648 16652 14700 16658
rect 14648 16594 14700 16600
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 14476 16046 14504 16526
rect 14464 16040 14516 16046
rect 14464 15982 14516 15988
rect 14476 15094 14504 15982
rect 14660 15978 14688 16594
rect 14752 16028 14780 17682
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14844 17066 14872 17478
rect 14832 17060 14884 17066
rect 14832 17002 14884 17008
rect 14936 16046 14964 17682
rect 15382 17096 15438 17105
rect 15382 17031 15438 17040
rect 15396 16794 15424 17031
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 15764 16658 15792 19178
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 15906 18524 16202 18544
rect 15962 18522 15986 18524
rect 16042 18522 16066 18524
rect 16122 18522 16146 18524
rect 15984 18470 15986 18522
rect 16048 18470 16060 18522
rect 16122 18470 16124 18522
rect 15962 18468 15986 18470
rect 16042 18468 16066 18470
rect 16122 18468 16146 18470
rect 15906 18448 16202 18468
rect 16316 17814 16344 18566
rect 16304 17808 16356 17814
rect 16304 17750 16356 17756
rect 15906 17436 16202 17456
rect 15962 17434 15986 17436
rect 16042 17434 16066 17436
rect 16122 17434 16146 17436
rect 15984 17382 15986 17434
rect 16048 17382 16060 17434
rect 16122 17382 16124 17434
rect 15962 17380 15986 17382
rect 16042 17380 16066 17382
rect 16122 17380 16146 17382
rect 15906 17360 16202 17380
rect 16120 17264 16172 17270
rect 16120 17206 16172 17212
rect 16132 16658 16160 17206
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16408 16794 16436 17070
rect 16396 16788 16448 16794
rect 16396 16730 16448 16736
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 15906 16348 16202 16368
rect 15962 16346 15986 16348
rect 16042 16346 16066 16348
rect 16122 16346 16146 16348
rect 15984 16294 15986 16346
rect 16048 16294 16060 16346
rect 16122 16294 16124 16346
rect 15962 16292 15986 16294
rect 16042 16292 16066 16294
rect 16122 16292 16146 16294
rect 15906 16272 16202 16292
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 14832 16040 14884 16046
rect 14752 16000 14832 16028
rect 14832 15982 14884 15988
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 14648 15972 14700 15978
rect 14648 15914 14700 15920
rect 14464 15088 14516 15094
rect 14464 15030 14516 15036
rect 14476 14890 14504 15030
rect 14660 14958 14688 15914
rect 14844 15026 14872 15982
rect 14936 15706 14964 15982
rect 15016 15904 15068 15910
rect 15016 15846 15068 15852
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 15028 15638 15056 15846
rect 15580 15638 15608 15846
rect 15016 15632 15068 15638
rect 15016 15574 15068 15580
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14464 14884 14516 14890
rect 14464 14826 14516 14832
rect 14660 14618 14688 14894
rect 15108 14884 15160 14890
rect 15108 14826 15160 14832
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14476 11762 14504 13874
rect 15028 13870 15056 14418
rect 15120 13938 15148 14826
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14936 12986 14964 13806
rect 15028 13530 15056 13806
rect 15120 13734 15148 13874
rect 15212 13870 15240 14758
rect 15764 14618 15792 16118
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16224 15745 16252 15982
rect 16210 15736 16266 15745
rect 16210 15671 16266 15680
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 15906 15260 16202 15280
rect 15962 15258 15986 15260
rect 16042 15258 16066 15260
rect 16122 15258 16146 15260
rect 15984 15206 15986 15258
rect 16048 15206 16060 15258
rect 16122 15206 16124 15258
rect 15962 15204 15986 15206
rect 16042 15204 16066 15206
rect 16122 15204 16146 15206
rect 15906 15184 16202 15204
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16224 14618 16252 14894
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15108 13728 15160 13734
rect 15108 13670 15160 13676
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 15764 13410 15792 14554
rect 16316 14482 16344 15302
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 15906 14172 16202 14192
rect 15962 14170 15986 14172
rect 16042 14170 16066 14172
rect 16122 14170 16146 14172
rect 15984 14118 15986 14170
rect 16048 14118 16060 14170
rect 16122 14118 16124 14170
rect 15962 14116 15986 14118
rect 16042 14116 16066 14118
rect 16122 14116 16146 14118
rect 15906 14096 16202 14116
rect 15936 13796 15988 13802
rect 15936 13738 15988 13744
rect 15948 13530 15976 13738
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 15764 13394 15884 13410
rect 15108 13388 15160 13394
rect 15764 13388 15896 13394
rect 15764 13382 15844 13388
rect 15108 13330 15160 13336
rect 15844 13330 15896 13336
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 15028 12782 15056 13262
rect 15120 12918 15148 13330
rect 16316 13258 16344 14418
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 15752 13252 15804 13258
rect 15752 13194 15804 13200
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15304 12986 15332 13126
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15108 12912 15160 12918
rect 15108 12854 15160 12860
rect 15764 12782 15792 13194
rect 15906 13084 16202 13104
rect 15962 13082 15986 13084
rect 16042 13082 16066 13084
rect 16122 13082 16146 13084
rect 15984 13030 15986 13082
rect 16048 13030 16060 13082
rect 16122 13030 16124 13082
rect 15962 13028 15986 13030
rect 16042 13028 16066 13030
rect 16122 13028 16146 13030
rect 15906 13008 16202 13028
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 14924 12368 14976 12374
rect 14924 12310 14976 12316
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14936 11150 14964 12310
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15212 11626 15240 12038
rect 15764 11762 15792 12718
rect 15906 11996 16202 12016
rect 15962 11994 15986 11996
rect 16042 11994 16066 11996
rect 16122 11994 16146 11996
rect 15984 11942 15986 11994
rect 16048 11942 16060 11994
rect 16122 11942 16124 11994
rect 15962 11940 15986 11942
rect 16042 11940 16066 11942
rect 16122 11940 16146 11942
rect 15906 11920 16202 11940
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15200 11620 15252 11626
rect 15200 11562 15252 11568
rect 16408 11286 16436 13806
rect 16396 11280 16448 11286
rect 16396 11222 16448 11228
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12728 9110 12756 9318
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 12820 8634 12848 9454
rect 12916 9276 13212 9296
rect 12972 9274 12996 9276
rect 13052 9274 13076 9276
rect 13132 9274 13156 9276
rect 12994 9222 12996 9274
rect 13058 9222 13070 9274
rect 13132 9222 13134 9274
rect 12972 9220 12996 9222
rect 13052 9220 13076 9222
rect 13132 9220 13156 9222
rect 12916 9200 13212 9220
rect 13280 9042 13308 9522
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 14476 8430 14504 8774
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 12916 8188 13212 8208
rect 12972 8186 12996 8188
rect 13052 8186 13076 8188
rect 13132 8186 13156 8188
rect 12994 8134 12996 8186
rect 13058 8134 13070 8186
rect 13132 8134 13134 8186
rect 12972 8132 12996 8134
rect 13052 8132 13076 8134
rect 13132 8132 13156 8134
rect 12916 8112 13212 8132
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12636 7342 12664 7890
rect 13372 7546 13400 8026
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12916 7100 13212 7120
rect 12972 7098 12996 7100
rect 13052 7098 13076 7100
rect 13132 7098 13156 7100
rect 12994 7046 12996 7098
rect 13058 7046 13070 7098
rect 13132 7046 13134 7098
rect 12972 7044 12996 7046
rect 13052 7044 13076 7046
rect 13132 7044 13156 7046
rect 12916 7024 13212 7044
rect 13372 7002 13400 7482
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13464 6866 13492 7278
rect 13648 7002 13676 7754
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12728 6390 12756 6598
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12728 5846 12756 6054
rect 12916 6012 13212 6032
rect 12972 6010 12996 6012
rect 13052 6010 13076 6012
rect 13132 6010 13156 6012
rect 12994 5958 12996 6010
rect 13058 5958 13070 6010
rect 13132 5958 13134 6010
rect 12972 5956 12996 5958
rect 13052 5956 13076 5958
rect 13132 5956 13156 5958
rect 12916 5936 13212 5956
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12728 5166 12756 5782
rect 13464 5778 13492 6802
rect 14568 6798 14596 7278
rect 14936 6866 14964 11086
rect 15906 10908 16202 10928
rect 15962 10906 15986 10908
rect 16042 10906 16066 10908
rect 16122 10906 16146 10908
rect 15984 10854 15986 10906
rect 16048 10854 16060 10906
rect 16122 10854 16124 10906
rect 15962 10852 15986 10854
rect 16042 10852 16066 10854
rect 16122 10852 16146 10854
rect 15906 10832 16202 10852
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15016 10532 15068 10538
rect 15016 10474 15068 10480
rect 15028 10198 15056 10474
rect 15016 10192 15068 10198
rect 15016 10134 15068 10140
rect 15120 9994 15148 10542
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 15108 9988 15160 9994
rect 15108 9930 15160 9936
rect 15120 9586 15148 9930
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15304 9382 15332 10474
rect 15396 9518 15424 10542
rect 16500 10470 16528 19654
rect 17512 19394 17540 21540
rect 18892 19990 18920 21540
rect 18880 19984 18932 19990
rect 18880 19926 18932 19932
rect 18052 19780 18104 19786
rect 18052 19722 18104 19728
rect 17512 19366 17632 19394
rect 17604 19310 17632 19366
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17776 19236 17828 19242
rect 17776 19178 17828 19184
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16960 18290 16988 18702
rect 17144 18426 17172 18770
rect 17132 18420 17184 18426
rect 17132 18362 17184 18368
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16960 17882 16988 18226
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 17328 17814 17356 19110
rect 17316 17808 17368 17814
rect 17316 17750 17368 17756
rect 16856 17264 16908 17270
rect 16856 17206 16908 17212
rect 16868 14618 16896 17206
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16960 15706 16988 16526
rect 17236 16250 17264 17138
rect 17788 17134 17816 19178
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 17972 17882 18000 18090
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17684 17060 17736 17066
rect 17684 17002 17736 17008
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17500 16040 17552 16046
rect 17500 15982 17552 15988
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16868 12374 16896 12582
rect 16856 12368 16908 12374
rect 16856 12310 16908 12316
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 17052 10266 17080 15846
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 17144 13734 17172 15506
rect 17420 14958 17448 15846
rect 17512 15094 17540 15982
rect 17604 15366 17632 15982
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17500 15088 17552 15094
rect 17500 15030 17552 15036
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17328 13870 17356 14554
rect 17512 14482 17540 15030
rect 17604 14958 17632 15302
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17696 14618 17724 17002
rect 17776 16176 17828 16182
rect 17776 16118 17828 16124
rect 17788 15570 17816 16118
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 17684 14612 17736 14618
rect 17684 14554 17736 14560
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17512 13870 17540 14418
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 17500 13864 17552 13870
rect 17500 13806 17552 13812
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17144 13326 17172 13670
rect 17328 13530 17356 13806
rect 17592 13796 17644 13802
rect 17592 13738 17644 13744
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17604 13376 17632 13738
rect 17696 13530 17724 13806
rect 17684 13524 17736 13530
rect 17684 13466 17736 13472
rect 17684 13388 17736 13394
rect 17604 13348 17684 13376
rect 17684 13330 17736 13336
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17144 12782 17172 13262
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17696 12714 17724 13330
rect 17788 12782 17816 15506
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17880 13705 17908 14418
rect 17866 13696 17922 13705
rect 17866 13631 17922 13640
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17420 11286 17448 11494
rect 17696 11354 17724 12650
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17972 11898 18000 12242
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17408 11280 17460 11286
rect 17408 11222 17460 11228
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 15906 9820 16202 9840
rect 15962 9818 15986 9820
rect 16042 9818 16066 9820
rect 16122 9818 16146 9820
rect 15984 9766 15986 9818
rect 16048 9766 16060 9818
rect 16122 9766 16124 9818
rect 15962 9764 15986 9766
rect 16042 9764 16066 9766
rect 16122 9764 16146 9766
rect 15906 9744 16202 9764
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15304 9178 15332 9318
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15396 9110 15424 9454
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15396 8430 15424 9046
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15672 8566 15700 8774
rect 15906 8732 16202 8752
rect 15962 8730 15986 8732
rect 16042 8730 16066 8732
rect 16122 8730 16146 8732
rect 15984 8678 15986 8730
rect 16048 8678 16060 8730
rect 16122 8678 16124 8730
rect 15962 8676 15986 8678
rect 16042 8676 16066 8678
rect 16122 8676 16146 8678
rect 15906 8656 16202 8676
rect 15660 8560 15712 8566
rect 15660 8502 15712 8508
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 16500 8362 16528 8978
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16592 8362 16620 8774
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15764 7342 15792 7822
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 15906 7644 16202 7664
rect 15962 7642 15986 7644
rect 16042 7642 16066 7644
rect 16122 7642 16146 7644
rect 15984 7590 15986 7642
rect 16048 7590 16060 7642
rect 16122 7590 16124 7642
rect 15962 7588 15986 7590
rect 16042 7588 16066 7590
rect 16122 7588 16146 7590
rect 15906 7568 16202 7588
rect 16316 7546 16344 7686
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 16316 6934 16344 7482
rect 16592 7342 16620 8298
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14924 6860 14976 6866
rect 14924 6802 14976 6808
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14660 6322 14688 6734
rect 14844 6662 14872 6802
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14752 6458 14780 6598
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 15488 5914 15516 6870
rect 15906 6556 16202 6576
rect 15962 6554 15986 6556
rect 16042 6554 16066 6556
rect 16122 6554 16146 6556
rect 15984 6502 15986 6554
rect 16048 6502 16060 6554
rect 16122 6502 16124 6554
rect 15962 6500 15986 6502
rect 16042 6500 16066 6502
rect 16122 6500 16146 6502
rect 15906 6480 16202 6500
rect 16396 6384 16448 6390
rect 16396 6326 16448 6332
rect 15936 6248 15988 6254
rect 15936 6190 15988 6196
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15580 5778 15608 6054
rect 15856 5846 15884 6054
rect 15948 5846 15976 6190
rect 15844 5840 15896 5846
rect 15844 5782 15896 5788
rect 15936 5840 15988 5846
rect 15936 5782 15988 5788
rect 13452 5772 13504 5778
rect 13452 5714 13504 5720
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 15120 5370 15148 5714
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15672 5234 15700 5646
rect 15906 5468 16202 5488
rect 15962 5466 15986 5468
rect 16042 5466 16066 5468
rect 16122 5466 16146 5468
rect 15984 5414 15986 5466
rect 16048 5414 16060 5466
rect 16122 5414 16124 5466
rect 15962 5412 15986 5414
rect 16042 5412 16066 5414
rect 16122 5412 16146 5414
rect 15906 5392 16202 5412
rect 16316 5370 16344 5714
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 16408 5166 16436 6326
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16500 5166 16528 5714
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 16396 5160 16448 5166
rect 16396 5102 16448 5108
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12636 4146 12664 4966
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12728 4214 12756 4626
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12532 3664 12584 3670
rect 12584 3612 12664 3618
rect 12532 3606 12664 3612
rect 12544 3590 12664 3606
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 11072 3194 11100 3402
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 12084 3194 12112 3334
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12084 3074 12112 3130
rect 12084 3046 12204 3074
rect 12176 2922 12204 3046
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 10888 2746 11008 2774
rect 10888 2650 10916 2746
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 11992 800 12020 2790
rect 12452 2514 12480 2926
rect 12544 2650 12572 3470
rect 12636 2990 12664 3590
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12728 2446 12756 4150
rect 12820 2854 12848 5102
rect 16028 5092 16080 5098
rect 16028 5034 16080 5040
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 12916 4924 13212 4944
rect 12972 4922 12996 4924
rect 13052 4922 13076 4924
rect 13132 4922 13156 4924
rect 12994 4870 12996 4922
rect 13058 4870 13070 4922
rect 13132 4870 13134 4922
rect 12972 4868 12996 4870
rect 13052 4868 13076 4870
rect 13132 4868 13156 4870
rect 12916 4848 13212 4868
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13544 4752 13596 4758
rect 13544 4694 13596 4700
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 12912 4282 12940 4558
rect 13268 4548 13320 4554
rect 13268 4490 13320 4496
rect 12900 4276 12952 4282
rect 12900 4218 12952 4224
rect 12912 4078 12940 4218
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 12916 3836 13212 3856
rect 12972 3834 12996 3836
rect 13052 3834 13076 3836
rect 13132 3834 13156 3836
rect 12994 3782 12996 3834
rect 13058 3782 13070 3834
rect 13132 3782 13134 3834
rect 12972 3780 12996 3782
rect 13052 3780 13076 3782
rect 13132 3780 13156 3782
rect 12916 3760 13212 3780
rect 13280 3738 13308 4490
rect 13556 4078 13584 4694
rect 13648 4146 13676 4762
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 13372 3738 13400 3946
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 12916 2748 13212 2768
rect 12972 2746 12996 2748
rect 13052 2746 13076 2748
rect 13132 2746 13156 2748
rect 12994 2694 12996 2746
rect 13058 2694 13070 2746
rect 13132 2694 13134 2746
rect 12972 2692 12996 2694
rect 13052 2692 13076 2694
rect 13132 2692 13156 2694
rect 12916 2672 13212 2692
rect 13464 2514 13492 3946
rect 13556 3602 13584 4014
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13556 2990 13584 3538
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 15028 3482 15056 3878
rect 15120 3602 15148 3878
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 14752 2990 14780 3470
rect 15028 3454 15148 3482
rect 15488 3466 15516 4966
rect 16040 4826 16068 5034
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 15906 4380 16202 4400
rect 15962 4378 15986 4380
rect 16042 4378 16066 4380
rect 16122 4378 16146 4380
rect 15984 4326 15986 4378
rect 16048 4326 16060 4378
rect 16122 4326 16124 4378
rect 15962 4324 15986 4326
rect 16042 4324 16066 4326
rect 16122 4324 16146 4326
rect 15906 4304 16202 4324
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15120 3398 15148 3454
rect 15476 3460 15528 3466
rect 15476 3402 15528 3408
rect 15108 3392 15160 3398
rect 15108 3334 15160 3340
rect 15120 3194 15148 3334
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15580 3058 15608 3606
rect 15906 3292 16202 3312
rect 15962 3290 15986 3292
rect 16042 3290 16066 3292
rect 16122 3290 16146 3292
rect 15984 3238 15986 3290
rect 16048 3238 16060 3290
rect 16122 3238 16124 3290
rect 15962 3236 15986 3238
rect 16042 3236 16066 3238
rect 16122 3236 16146 3238
rect 15906 3216 16202 3236
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14752 2650 14780 2926
rect 15580 2922 15608 2994
rect 16408 2922 16436 4626
rect 15568 2916 15620 2922
rect 15568 2858 15620 2864
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 16408 2582 16436 2858
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 16396 2576 16448 2582
rect 16396 2518 16448 2524
rect 13452 2508 13504 2514
rect 13452 2450 13504 2456
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 13832 800 13860 2450
rect 15212 800 15240 2518
rect 16500 2446 16528 5102
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16684 4622 16712 4966
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 16592 3534 16620 4490
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16592 3126 16620 3470
rect 16960 3194 16988 10066
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17512 9042 17540 9862
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17512 8430 17540 8978
rect 17696 8498 17724 9114
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17500 8424 17552 8430
rect 17500 8366 17552 8372
rect 17696 8090 17724 8434
rect 17880 8430 17908 8978
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 18064 6390 18092 19722
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 18144 16720 18196 16726
rect 18144 16662 18196 16668
rect 18156 15162 18184 16662
rect 18248 15706 18276 18566
rect 18326 18456 18382 18465
rect 18326 18391 18382 18400
rect 18340 18358 18368 18391
rect 18328 18352 18380 18358
rect 18328 18294 18380 18300
rect 18420 18148 18472 18154
rect 18420 18090 18472 18096
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 18340 15570 18368 16390
rect 18328 15564 18380 15570
rect 18328 15506 18380 15512
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18340 13190 18368 13466
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18340 12646 18368 13126
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18340 12442 18368 12582
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18326 11656 18382 11665
rect 18326 11591 18382 11600
rect 18340 10606 18368 11591
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18144 10192 18196 10198
rect 18144 10134 18196 10140
rect 18156 9654 18184 10134
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18326 9616 18382 9625
rect 18326 9551 18382 9560
rect 18340 9518 18368 9551
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18326 6896 18382 6905
rect 18326 6831 18328 6840
rect 18380 6831 18382 6840
rect 18328 6802 18380 6808
rect 18052 6384 18104 6390
rect 18052 6326 18104 6332
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17144 5914 17172 6190
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 17144 5302 17172 5850
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 18156 4826 18184 5510
rect 18326 4856 18382 4865
rect 18144 4820 18196 4826
rect 18326 4791 18382 4800
rect 18144 4762 18196 4768
rect 18340 4690 18368 4791
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18432 4554 18460 18090
rect 18512 17740 18564 17746
rect 18512 17682 18564 17688
rect 18524 14958 18552 17682
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 18524 11694 18552 14894
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18420 4548 18472 4554
rect 18420 4490 18472 4496
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 15906 2204 16202 2224
rect 15962 2202 15986 2204
rect 16042 2202 16066 2204
rect 16122 2202 16146 2204
rect 15984 2150 15986 2202
rect 16048 2150 16060 2202
rect 16122 2150 16124 2202
rect 15962 2148 15986 2150
rect 16042 2148 16066 2150
rect 16122 2148 16146 2150
rect 15906 2128 16202 2148
rect 16592 800 16620 2926
rect 17328 2650 17356 3334
rect 18156 3194 18184 3674
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18340 2825 18368 3538
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 18326 2816 18382 2825
rect 18326 2751 18382 2760
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 17960 2372 18012 2378
rect 17960 2314 18012 2320
rect 17972 800 18000 2314
rect 478 0 534 800
rect 1858 0 1914 800
rect 3238 0 3294 800
rect 4618 0 4674 800
rect 5998 0 6054 800
rect 7838 0 7894 800
rect 9218 0 9274 800
rect 10598 0 10654 800
rect 11978 0 12034 800
rect 13818 0 13874 800
rect 15198 0 15254 800
rect 16578 0 16634 800
rect 17958 0 18014 800
rect 18432 785 18460 2926
rect 18418 776 18474 785
rect 18418 711 18474 720
<< via2 >>
rect 1490 20440 1546 20496
rect 6936 20154 6992 20156
rect 7016 20154 7072 20156
rect 7096 20154 7152 20156
rect 7176 20154 7232 20156
rect 6936 20102 6962 20154
rect 6962 20102 6992 20154
rect 7016 20102 7026 20154
rect 7026 20102 7072 20154
rect 7096 20102 7142 20154
rect 7142 20102 7152 20154
rect 7176 20102 7206 20154
rect 7206 20102 7232 20154
rect 6936 20100 6992 20102
rect 7016 20100 7072 20102
rect 7096 20100 7152 20102
rect 7176 20100 7232 20102
rect 1398 17740 1454 17776
rect 1398 17720 1400 17740
rect 1400 17720 1452 17740
rect 1452 17720 1454 17740
rect 1398 15680 1454 15736
rect 1398 13640 1454 13696
rect 1490 11600 1546 11656
rect 1398 8900 1454 8936
rect 1398 8880 1400 8900
rect 1400 8880 1452 8900
rect 1452 8880 1454 8900
rect 3946 19610 4002 19612
rect 4026 19610 4082 19612
rect 4106 19610 4162 19612
rect 4186 19610 4242 19612
rect 3946 19558 3972 19610
rect 3972 19558 4002 19610
rect 4026 19558 4036 19610
rect 4036 19558 4082 19610
rect 4106 19558 4152 19610
rect 4152 19558 4162 19610
rect 4186 19558 4216 19610
rect 4216 19558 4242 19610
rect 3946 19556 4002 19558
rect 4026 19556 4082 19558
rect 4106 19556 4162 19558
rect 4186 19556 4242 19558
rect 3946 18522 4002 18524
rect 4026 18522 4082 18524
rect 4106 18522 4162 18524
rect 4186 18522 4242 18524
rect 3946 18470 3972 18522
rect 3972 18470 4002 18522
rect 4026 18470 4036 18522
rect 4036 18470 4082 18522
rect 4106 18470 4152 18522
rect 4152 18470 4162 18522
rect 4186 18470 4216 18522
rect 4216 18470 4242 18522
rect 3946 18468 4002 18470
rect 4026 18468 4082 18470
rect 4106 18468 4162 18470
rect 4186 18468 4242 18470
rect 3946 17434 4002 17436
rect 4026 17434 4082 17436
rect 4106 17434 4162 17436
rect 4186 17434 4242 17436
rect 3946 17382 3972 17434
rect 3972 17382 4002 17434
rect 4026 17382 4036 17434
rect 4036 17382 4082 17434
rect 4106 17382 4152 17434
rect 4152 17382 4162 17434
rect 4186 17382 4216 17434
rect 4216 17382 4242 17434
rect 3946 17380 4002 17382
rect 4026 17380 4082 17382
rect 4106 17380 4162 17382
rect 4186 17380 4242 17382
rect 3946 16346 4002 16348
rect 4026 16346 4082 16348
rect 4106 16346 4162 16348
rect 4186 16346 4242 16348
rect 3946 16294 3972 16346
rect 3972 16294 4002 16346
rect 4026 16294 4036 16346
rect 4036 16294 4082 16346
rect 4106 16294 4152 16346
rect 4152 16294 4162 16346
rect 4186 16294 4216 16346
rect 4216 16294 4242 16346
rect 3946 16292 4002 16294
rect 4026 16292 4082 16294
rect 4106 16292 4162 16294
rect 4186 16292 4242 16294
rect 3946 15258 4002 15260
rect 4026 15258 4082 15260
rect 4106 15258 4162 15260
rect 4186 15258 4242 15260
rect 3946 15206 3972 15258
rect 3972 15206 4002 15258
rect 4026 15206 4036 15258
rect 4036 15206 4082 15258
rect 4106 15206 4152 15258
rect 4152 15206 4162 15258
rect 4186 15206 4216 15258
rect 4216 15206 4242 15258
rect 3946 15204 4002 15206
rect 4026 15204 4082 15206
rect 4106 15204 4162 15206
rect 4186 15204 4242 15206
rect 3946 14170 4002 14172
rect 4026 14170 4082 14172
rect 4106 14170 4162 14172
rect 4186 14170 4242 14172
rect 3946 14118 3972 14170
rect 3972 14118 4002 14170
rect 4026 14118 4036 14170
rect 4036 14118 4082 14170
rect 4106 14118 4152 14170
rect 4152 14118 4162 14170
rect 4186 14118 4216 14170
rect 4216 14118 4242 14170
rect 3946 14116 4002 14118
rect 4026 14116 4082 14118
rect 4106 14116 4162 14118
rect 4186 14116 4242 14118
rect 3946 13082 4002 13084
rect 4026 13082 4082 13084
rect 4106 13082 4162 13084
rect 4186 13082 4242 13084
rect 3946 13030 3972 13082
rect 3972 13030 4002 13082
rect 4026 13030 4036 13082
rect 4036 13030 4082 13082
rect 4106 13030 4152 13082
rect 4152 13030 4162 13082
rect 4186 13030 4216 13082
rect 4216 13030 4242 13082
rect 3946 13028 4002 13030
rect 4026 13028 4082 13030
rect 4106 13028 4162 13030
rect 4186 13028 4242 13030
rect 3946 11994 4002 11996
rect 4026 11994 4082 11996
rect 4106 11994 4162 11996
rect 4186 11994 4242 11996
rect 3946 11942 3972 11994
rect 3972 11942 4002 11994
rect 4026 11942 4036 11994
rect 4036 11942 4082 11994
rect 4106 11942 4152 11994
rect 4152 11942 4162 11994
rect 4186 11942 4216 11994
rect 4216 11942 4242 11994
rect 3946 11940 4002 11942
rect 4026 11940 4082 11942
rect 4106 11940 4162 11942
rect 4186 11940 4242 11942
rect 3946 10906 4002 10908
rect 4026 10906 4082 10908
rect 4106 10906 4162 10908
rect 4186 10906 4242 10908
rect 3946 10854 3972 10906
rect 3972 10854 4002 10906
rect 4026 10854 4036 10906
rect 4036 10854 4082 10906
rect 4106 10854 4152 10906
rect 4152 10854 4162 10906
rect 4186 10854 4216 10906
rect 4216 10854 4242 10906
rect 3946 10852 4002 10854
rect 4026 10852 4082 10854
rect 4106 10852 4162 10854
rect 4186 10852 4242 10854
rect 1398 6840 1454 6896
rect 3946 9818 4002 9820
rect 4026 9818 4082 9820
rect 4106 9818 4162 9820
rect 4186 9818 4242 9820
rect 3946 9766 3972 9818
rect 3972 9766 4002 9818
rect 4026 9766 4036 9818
rect 4036 9766 4082 9818
rect 4106 9766 4152 9818
rect 4152 9766 4162 9818
rect 4186 9766 4216 9818
rect 4216 9766 4242 9818
rect 3946 9764 4002 9766
rect 4026 9764 4082 9766
rect 4106 9764 4162 9766
rect 4186 9764 4242 9766
rect 3946 8730 4002 8732
rect 4026 8730 4082 8732
rect 4106 8730 4162 8732
rect 4186 8730 4242 8732
rect 3946 8678 3972 8730
rect 3972 8678 4002 8730
rect 4026 8678 4036 8730
rect 4036 8678 4082 8730
rect 4106 8678 4152 8730
rect 4152 8678 4162 8730
rect 4186 8678 4216 8730
rect 4216 8678 4242 8730
rect 3946 8676 4002 8678
rect 4026 8676 4082 8678
rect 4106 8676 4162 8678
rect 4186 8676 4242 8678
rect 1490 4820 1546 4856
rect 1490 4800 1492 4820
rect 1492 4800 1544 4820
rect 1544 4800 1546 4820
rect 1398 2760 1454 2816
rect 3946 7642 4002 7644
rect 4026 7642 4082 7644
rect 4106 7642 4162 7644
rect 4186 7642 4242 7644
rect 3946 7590 3972 7642
rect 3972 7590 4002 7642
rect 4026 7590 4036 7642
rect 4036 7590 4082 7642
rect 4106 7590 4152 7642
rect 4152 7590 4162 7642
rect 4186 7590 4216 7642
rect 4216 7590 4242 7642
rect 3946 7588 4002 7590
rect 4026 7588 4082 7590
rect 4106 7588 4162 7590
rect 4186 7588 4242 7590
rect 3946 6554 4002 6556
rect 4026 6554 4082 6556
rect 4106 6554 4162 6556
rect 4186 6554 4242 6556
rect 3946 6502 3972 6554
rect 3972 6502 4002 6554
rect 4026 6502 4036 6554
rect 4036 6502 4082 6554
rect 4106 6502 4152 6554
rect 4152 6502 4162 6554
rect 4186 6502 4216 6554
rect 4216 6502 4242 6554
rect 3946 6500 4002 6502
rect 4026 6500 4082 6502
rect 4106 6500 4162 6502
rect 4186 6500 4242 6502
rect 3946 5466 4002 5468
rect 4026 5466 4082 5468
rect 4106 5466 4162 5468
rect 4186 5466 4242 5468
rect 3946 5414 3972 5466
rect 3972 5414 4002 5466
rect 4026 5414 4036 5466
rect 4036 5414 4082 5466
rect 4106 5414 4152 5466
rect 4152 5414 4162 5466
rect 4186 5414 4216 5466
rect 4216 5414 4242 5466
rect 3946 5412 4002 5414
rect 4026 5412 4082 5414
rect 4106 5412 4162 5414
rect 4186 5412 4242 5414
rect 3946 4378 4002 4380
rect 4026 4378 4082 4380
rect 4106 4378 4162 4380
rect 4186 4378 4242 4380
rect 3946 4326 3972 4378
rect 3972 4326 4002 4378
rect 4026 4326 4036 4378
rect 4036 4326 4082 4378
rect 4106 4326 4152 4378
rect 4152 4326 4162 4378
rect 4186 4326 4216 4378
rect 4216 4326 4242 4378
rect 3946 4324 4002 4326
rect 4026 4324 4082 4326
rect 4106 4324 4162 4326
rect 4186 4324 4242 4326
rect 3946 3290 4002 3292
rect 4026 3290 4082 3292
rect 4106 3290 4162 3292
rect 4186 3290 4242 3292
rect 3946 3238 3972 3290
rect 3972 3238 4002 3290
rect 4026 3238 4036 3290
rect 4036 3238 4082 3290
rect 4106 3238 4152 3290
rect 4152 3238 4162 3290
rect 4186 3238 4216 3290
rect 4216 3238 4242 3290
rect 3946 3236 4002 3238
rect 4026 3236 4082 3238
rect 4106 3236 4162 3238
rect 4186 3236 4242 3238
rect 12916 20154 12972 20156
rect 12996 20154 13052 20156
rect 13076 20154 13132 20156
rect 13156 20154 13212 20156
rect 12916 20102 12942 20154
rect 12942 20102 12972 20154
rect 12996 20102 13006 20154
rect 13006 20102 13052 20154
rect 13076 20102 13122 20154
rect 13122 20102 13132 20154
rect 13156 20102 13186 20154
rect 13186 20102 13212 20154
rect 12916 20100 12972 20102
rect 12996 20100 13052 20102
rect 13076 20100 13132 20102
rect 13156 20100 13212 20102
rect 16486 20440 16542 20496
rect 6936 19066 6992 19068
rect 7016 19066 7072 19068
rect 7096 19066 7152 19068
rect 7176 19066 7232 19068
rect 6936 19014 6962 19066
rect 6962 19014 6992 19066
rect 7016 19014 7026 19066
rect 7026 19014 7072 19066
rect 7096 19014 7142 19066
rect 7142 19014 7152 19066
rect 7176 19014 7206 19066
rect 7206 19014 7232 19066
rect 6936 19012 6992 19014
rect 7016 19012 7072 19014
rect 7096 19012 7152 19014
rect 7176 19012 7232 19014
rect 6936 17978 6992 17980
rect 7016 17978 7072 17980
rect 7096 17978 7152 17980
rect 7176 17978 7232 17980
rect 6936 17926 6962 17978
rect 6962 17926 6992 17978
rect 7016 17926 7026 17978
rect 7026 17926 7072 17978
rect 7096 17926 7142 17978
rect 7142 17926 7152 17978
rect 7176 17926 7206 17978
rect 7206 17926 7232 17978
rect 6936 17924 6992 17926
rect 7016 17924 7072 17926
rect 7096 17924 7152 17926
rect 7176 17924 7232 17926
rect 6936 16890 6992 16892
rect 7016 16890 7072 16892
rect 7096 16890 7152 16892
rect 7176 16890 7232 16892
rect 6936 16838 6962 16890
rect 6962 16838 6992 16890
rect 7016 16838 7026 16890
rect 7026 16838 7072 16890
rect 7096 16838 7142 16890
rect 7142 16838 7152 16890
rect 7176 16838 7206 16890
rect 7206 16838 7232 16890
rect 6936 16836 6992 16838
rect 7016 16836 7072 16838
rect 7096 16836 7152 16838
rect 7176 16836 7232 16838
rect 6936 15802 6992 15804
rect 7016 15802 7072 15804
rect 7096 15802 7152 15804
rect 7176 15802 7232 15804
rect 6936 15750 6962 15802
rect 6962 15750 6992 15802
rect 7016 15750 7026 15802
rect 7026 15750 7072 15802
rect 7096 15750 7142 15802
rect 7142 15750 7152 15802
rect 7176 15750 7206 15802
rect 7206 15750 7232 15802
rect 6936 15748 6992 15750
rect 7016 15748 7072 15750
rect 7096 15748 7152 15750
rect 7176 15748 7232 15750
rect 6936 14714 6992 14716
rect 7016 14714 7072 14716
rect 7096 14714 7152 14716
rect 7176 14714 7232 14716
rect 6936 14662 6962 14714
rect 6962 14662 6992 14714
rect 7016 14662 7026 14714
rect 7026 14662 7072 14714
rect 7096 14662 7142 14714
rect 7142 14662 7152 14714
rect 7176 14662 7206 14714
rect 7206 14662 7232 14714
rect 6936 14660 6992 14662
rect 7016 14660 7072 14662
rect 7096 14660 7152 14662
rect 7176 14660 7232 14662
rect 6936 13626 6992 13628
rect 7016 13626 7072 13628
rect 7096 13626 7152 13628
rect 7176 13626 7232 13628
rect 6936 13574 6962 13626
rect 6962 13574 6992 13626
rect 7016 13574 7026 13626
rect 7026 13574 7072 13626
rect 7096 13574 7142 13626
rect 7142 13574 7152 13626
rect 7176 13574 7206 13626
rect 7206 13574 7232 13626
rect 6936 13572 6992 13574
rect 7016 13572 7072 13574
rect 7096 13572 7152 13574
rect 7176 13572 7232 13574
rect 6936 12538 6992 12540
rect 7016 12538 7072 12540
rect 7096 12538 7152 12540
rect 7176 12538 7232 12540
rect 6936 12486 6962 12538
rect 6962 12486 6992 12538
rect 7016 12486 7026 12538
rect 7026 12486 7072 12538
rect 7096 12486 7142 12538
rect 7142 12486 7152 12538
rect 7176 12486 7206 12538
rect 7206 12486 7232 12538
rect 6936 12484 6992 12486
rect 7016 12484 7072 12486
rect 7096 12484 7152 12486
rect 7176 12484 7232 12486
rect 6936 11450 6992 11452
rect 7016 11450 7072 11452
rect 7096 11450 7152 11452
rect 7176 11450 7232 11452
rect 6936 11398 6962 11450
rect 6962 11398 6992 11450
rect 7016 11398 7026 11450
rect 7026 11398 7072 11450
rect 7096 11398 7142 11450
rect 7142 11398 7152 11450
rect 7176 11398 7206 11450
rect 7206 11398 7232 11450
rect 6936 11396 6992 11398
rect 7016 11396 7072 11398
rect 7096 11396 7152 11398
rect 7176 11396 7232 11398
rect 9926 19610 9982 19612
rect 10006 19610 10062 19612
rect 10086 19610 10142 19612
rect 10166 19610 10222 19612
rect 9926 19558 9952 19610
rect 9952 19558 9982 19610
rect 10006 19558 10016 19610
rect 10016 19558 10062 19610
rect 10086 19558 10132 19610
rect 10132 19558 10142 19610
rect 10166 19558 10196 19610
rect 10196 19558 10222 19610
rect 9926 19556 9982 19558
rect 10006 19556 10062 19558
rect 10086 19556 10142 19558
rect 10166 19556 10222 19558
rect 9926 18522 9982 18524
rect 10006 18522 10062 18524
rect 10086 18522 10142 18524
rect 10166 18522 10222 18524
rect 9926 18470 9952 18522
rect 9952 18470 9982 18522
rect 10006 18470 10016 18522
rect 10016 18470 10062 18522
rect 10086 18470 10132 18522
rect 10132 18470 10142 18522
rect 10166 18470 10196 18522
rect 10196 18470 10222 18522
rect 9926 18468 9982 18470
rect 10006 18468 10062 18470
rect 10086 18468 10142 18470
rect 10166 18468 10222 18470
rect 9926 17434 9982 17436
rect 10006 17434 10062 17436
rect 10086 17434 10142 17436
rect 10166 17434 10222 17436
rect 9926 17382 9952 17434
rect 9952 17382 9982 17434
rect 10006 17382 10016 17434
rect 10016 17382 10062 17434
rect 10086 17382 10132 17434
rect 10132 17382 10142 17434
rect 10166 17382 10196 17434
rect 10196 17382 10222 17434
rect 9926 17380 9982 17382
rect 10006 17380 10062 17382
rect 10086 17380 10142 17382
rect 10166 17380 10222 17382
rect 6936 10362 6992 10364
rect 7016 10362 7072 10364
rect 7096 10362 7152 10364
rect 7176 10362 7232 10364
rect 6936 10310 6962 10362
rect 6962 10310 6992 10362
rect 7016 10310 7026 10362
rect 7026 10310 7072 10362
rect 7096 10310 7142 10362
rect 7142 10310 7152 10362
rect 7176 10310 7206 10362
rect 7206 10310 7232 10362
rect 6936 10308 6992 10310
rect 7016 10308 7072 10310
rect 7096 10308 7152 10310
rect 7176 10308 7232 10310
rect 6936 9274 6992 9276
rect 7016 9274 7072 9276
rect 7096 9274 7152 9276
rect 7176 9274 7232 9276
rect 6936 9222 6962 9274
rect 6962 9222 6992 9274
rect 7016 9222 7026 9274
rect 7026 9222 7072 9274
rect 7096 9222 7142 9274
rect 7142 9222 7152 9274
rect 7176 9222 7206 9274
rect 7206 9222 7232 9274
rect 6936 9220 6992 9222
rect 7016 9220 7072 9222
rect 7096 9220 7152 9222
rect 7176 9220 7232 9222
rect 6936 8186 6992 8188
rect 7016 8186 7072 8188
rect 7096 8186 7152 8188
rect 7176 8186 7232 8188
rect 6936 8134 6962 8186
rect 6962 8134 6992 8186
rect 7016 8134 7026 8186
rect 7026 8134 7072 8186
rect 7096 8134 7142 8186
rect 7142 8134 7152 8186
rect 7176 8134 7206 8186
rect 7206 8134 7232 8186
rect 6936 8132 6992 8134
rect 7016 8132 7072 8134
rect 7096 8132 7152 8134
rect 7176 8132 7232 8134
rect 6936 7098 6992 7100
rect 7016 7098 7072 7100
rect 7096 7098 7152 7100
rect 7176 7098 7232 7100
rect 6936 7046 6962 7098
rect 6962 7046 6992 7098
rect 7016 7046 7026 7098
rect 7026 7046 7072 7098
rect 7096 7046 7142 7098
rect 7142 7046 7152 7098
rect 7176 7046 7206 7098
rect 7206 7046 7232 7098
rect 6936 7044 6992 7046
rect 7016 7044 7072 7046
rect 7096 7044 7152 7046
rect 7176 7044 7232 7046
rect 6936 6010 6992 6012
rect 7016 6010 7072 6012
rect 7096 6010 7152 6012
rect 7176 6010 7232 6012
rect 6936 5958 6962 6010
rect 6962 5958 6992 6010
rect 7016 5958 7026 6010
rect 7026 5958 7072 6010
rect 7096 5958 7142 6010
rect 7142 5958 7152 6010
rect 7176 5958 7206 6010
rect 7206 5958 7232 6010
rect 6936 5956 6992 5958
rect 7016 5956 7072 5958
rect 7096 5956 7152 5958
rect 7176 5956 7232 5958
rect 6936 4922 6992 4924
rect 7016 4922 7072 4924
rect 7096 4922 7152 4924
rect 7176 4922 7232 4924
rect 6936 4870 6962 4922
rect 6962 4870 6992 4922
rect 7016 4870 7026 4922
rect 7026 4870 7072 4922
rect 7096 4870 7142 4922
rect 7142 4870 7152 4922
rect 7176 4870 7206 4922
rect 7206 4870 7232 4922
rect 6936 4868 6992 4870
rect 7016 4868 7072 4870
rect 7096 4868 7152 4870
rect 7176 4868 7232 4870
rect 6936 3834 6992 3836
rect 7016 3834 7072 3836
rect 7096 3834 7152 3836
rect 7176 3834 7232 3836
rect 6936 3782 6962 3834
rect 6962 3782 6992 3834
rect 7016 3782 7026 3834
rect 7026 3782 7072 3834
rect 7096 3782 7142 3834
rect 7142 3782 7152 3834
rect 7176 3782 7206 3834
rect 7206 3782 7232 3834
rect 6936 3780 6992 3782
rect 7016 3780 7072 3782
rect 7096 3780 7152 3782
rect 7176 3780 7232 3782
rect 9926 16346 9982 16348
rect 10006 16346 10062 16348
rect 10086 16346 10142 16348
rect 10166 16346 10222 16348
rect 9926 16294 9952 16346
rect 9952 16294 9982 16346
rect 10006 16294 10016 16346
rect 10016 16294 10062 16346
rect 10086 16294 10132 16346
rect 10132 16294 10142 16346
rect 10166 16294 10196 16346
rect 10196 16294 10222 16346
rect 9926 16292 9982 16294
rect 10006 16292 10062 16294
rect 10086 16292 10142 16294
rect 10166 16292 10222 16294
rect 9926 15258 9982 15260
rect 10006 15258 10062 15260
rect 10086 15258 10142 15260
rect 10166 15258 10222 15260
rect 9926 15206 9952 15258
rect 9952 15206 9982 15258
rect 10006 15206 10016 15258
rect 10016 15206 10062 15258
rect 10086 15206 10132 15258
rect 10132 15206 10142 15258
rect 10166 15206 10196 15258
rect 10196 15206 10222 15258
rect 9926 15204 9982 15206
rect 10006 15204 10062 15206
rect 10086 15204 10142 15206
rect 10166 15204 10222 15206
rect 9926 14170 9982 14172
rect 10006 14170 10062 14172
rect 10086 14170 10142 14172
rect 10166 14170 10222 14172
rect 9926 14118 9952 14170
rect 9952 14118 9982 14170
rect 10006 14118 10016 14170
rect 10016 14118 10062 14170
rect 10086 14118 10132 14170
rect 10132 14118 10142 14170
rect 10166 14118 10196 14170
rect 10196 14118 10222 14170
rect 9926 14116 9982 14118
rect 10006 14116 10062 14118
rect 10086 14116 10142 14118
rect 10166 14116 10222 14118
rect 9926 13082 9982 13084
rect 10006 13082 10062 13084
rect 10086 13082 10142 13084
rect 10166 13082 10222 13084
rect 9926 13030 9952 13082
rect 9952 13030 9982 13082
rect 10006 13030 10016 13082
rect 10016 13030 10062 13082
rect 10086 13030 10132 13082
rect 10132 13030 10142 13082
rect 10166 13030 10196 13082
rect 10196 13030 10222 13082
rect 9926 13028 9982 13030
rect 10006 13028 10062 13030
rect 10086 13028 10142 13030
rect 10166 13028 10222 13030
rect 6936 2746 6992 2748
rect 7016 2746 7072 2748
rect 7096 2746 7152 2748
rect 7176 2746 7232 2748
rect 6936 2694 6962 2746
rect 6962 2694 6992 2746
rect 7016 2694 7026 2746
rect 7026 2694 7072 2746
rect 7096 2694 7142 2746
rect 7142 2694 7152 2746
rect 7176 2694 7206 2746
rect 7206 2694 7232 2746
rect 6936 2692 6992 2694
rect 7016 2692 7072 2694
rect 7096 2692 7152 2694
rect 7176 2692 7232 2694
rect 9926 11994 9982 11996
rect 10006 11994 10062 11996
rect 10086 11994 10142 11996
rect 10166 11994 10222 11996
rect 9926 11942 9952 11994
rect 9952 11942 9982 11994
rect 10006 11942 10016 11994
rect 10016 11942 10062 11994
rect 10086 11942 10132 11994
rect 10132 11942 10142 11994
rect 10166 11942 10196 11994
rect 10196 11942 10222 11994
rect 9926 11940 9982 11942
rect 10006 11940 10062 11942
rect 10086 11940 10142 11942
rect 10166 11940 10222 11942
rect 10782 17076 10784 17096
rect 10784 17076 10836 17096
rect 10836 17076 10838 17096
rect 10782 17040 10838 17076
rect 9926 10906 9982 10908
rect 10006 10906 10062 10908
rect 10086 10906 10142 10908
rect 10166 10906 10222 10908
rect 9926 10854 9952 10906
rect 9952 10854 9982 10906
rect 10006 10854 10016 10906
rect 10016 10854 10062 10906
rect 10086 10854 10132 10906
rect 10132 10854 10142 10906
rect 10166 10854 10196 10906
rect 10196 10854 10222 10906
rect 9926 10852 9982 10854
rect 10006 10852 10062 10854
rect 10086 10852 10142 10854
rect 10166 10852 10222 10854
rect 9926 9818 9982 9820
rect 10006 9818 10062 9820
rect 10086 9818 10142 9820
rect 10166 9818 10222 9820
rect 9926 9766 9952 9818
rect 9952 9766 9982 9818
rect 10006 9766 10016 9818
rect 10016 9766 10062 9818
rect 10086 9766 10132 9818
rect 10132 9766 10142 9818
rect 10166 9766 10196 9818
rect 10196 9766 10222 9818
rect 9926 9764 9982 9766
rect 10006 9764 10062 9766
rect 10086 9764 10142 9766
rect 10166 9764 10222 9766
rect 9926 8730 9982 8732
rect 10006 8730 10062 8732
rect 10086 8730 10142 8732
rect 10166 8730 10222 8732
rect 9926 8678 9952 8730
rect 9952 8678 9982 8730
rect 10006 8678 10016 8730
rect 10016 8678 10062 8730
rect 10086 8678 10132 8730
rect 10132 8678 10142 8730
rect 10166 8678 10196 8730
rect 10196 8678 10222 8730
rect 9926 8676 9982 8678
rect 10006 8676 10062 8678
rect 10086 8676 10142 8678
rect 10166 8676 10222 8678
rect 3946 2202 4002 2204
rect 4026 2202 4082 2204
rect 4106 2202 4162 2204
rect 4186 2202 4242 2204
rect 3946 2150 3972 2202
rect 3972 2150 4002 2202
rect 4026 2150 4036 2202
rect 4036 2150 4082 2202
rect 4106 2150 4152 2202
rect 4152 2150 4162 2202
rect 4186 2150 4216 2202
rect 4216 2150 4242 2202
rect 3946 2148 4002 2150
rect 4026 2148 4082 2150
rect 4106 2148 4162 2150
rect 4186 2148 4242 2150
rect 9926 7642 9982 7644
rect 10006 7642 10062 7644
rect 10086 7642 10142 7644
rect 10166 7642 10222 7644
rect 9926 7590 9952 7642
rect 9952 7590 9982 7642
rect 10006 7590 10016 7642
rect 10016 7590 10062 7642
rect 10086 7590 10132 7642
rect 10132 7590 10142 7642
rect 10166 7590 10196 7642
rect 10196 7590 10222 7642
rect 9926 7588 9982 7590
rect 10006 7588 10062 7590
rect 10086 7588 10142 7590
rect 10166 7588 10222 7590
rect 9926 6554 9982 6556
rect 10006 6554 10062 6556
rect 10086 6554 10142 6556
rect 10166 6554 10222 6556
rect 9926 6502 9952 6554
rect 9952 6502 9982 6554
rect 10006 6502 10016 6554
rect 10016 6502 10062 6554
rect 10086 6502 10132 6554
rect 10132 6502 10142 6554
rect 10166 6502 10196 6554
rect 10196 6502 10222 6554
rect 9926 6500 9982 6502
rect 10006 6500 10062 6502
rect 10086 6500 10142 6502
rect 10166 6500 10222 6502
rect 9926 5466 9982 5468
rect 10006 5466 10062 5468
rect 10086 5466 10142 5468
rect 10166 5466 10222 5468
rect 9926 5414 9952 5466
rect 9952 5414 9982 5466
rect 10006 5414 10016 5466
rect 10016 5414 10062 5466
rect 10086 5414 10132 5466
rect 10132 5414 10142 5466
rect 10166 5414 10196 5466
rect 10196 5414 10222 5466
rect 9926 5412 9982 5414
rect 10006 5412 10062 5414
rect 10086 5412 10142 5414
rect 10166 5412 10222 5414
rect 9926 4378 9982 4380
rect 10006 4378 10062 4380
rect 10086 4378 10142 4380
rect 10166 4378 10222 4380
rect 9926 4326 9952 4378
rect 9952 4326 9982 4378
rect 10006 4326 10016 4378
rect 10016 4326 10062 4378
rect 10086 4326 10132 4378
rect 10132 4326 10142 4378
rect 10166 4326 10196 4378
rect 10196 4326 10222 4378
rect 9926 4324 9982 4326
rect 10006 4324 10062 4326
rect 10086 4324 10142 4326
rect 10166 4324 10222 4326
rect 9926 3290 9982 3292
rect 10006 3290 10062 3292
rect 10086 3290 10142 3292
rect 10166 3290 10222 3292
rect 9926 3238 9952 3290
rect 9952 3238 9982 3290
rect 10006 3238 10016 3290
rect 10016 3238 10062 3290
rect 10086 3238 10132 3290
rect 10132 3238 10142 3290
rect 10166 3238 10196 3290
rect 10196 3238 10222 3290
rect 9926 3236 9982 3238
rect 10006 3236 10062 3238
rect 10086 3236 10142 3238
rect 10166 3236 10222 3238
rect 9926 2202 9982 2204
rect 10006 2202 10062 2204
rect 10086 2202 10142 2204
rect 10166 2202 10222 2204
rect 9926 2150 9952 2202
rect 9952 2150 9982 2202
rect 10006 2150 10016 2202
rect 10016 2150 10062 2202
rect 10086 2150 10132 2202
rect 10132 2150 10142 2202
rect 10166 2150 10196 2202
rect 10196 2150 10222 2202
rect 9926 2148 9982 2150
rect 10006 2148 10062 2150
rect 10086 2148 10142 2150
rect 10166 2148 10222 2150
rect 12916 19066 12972 19068
rect 12996 19066 13052 19068
rect 13076 19066 13132 19068
rect 13156 19066 13212 19068
rect 12916 19014 12942 19066
rect 12942 19014 12972 19066
rect 12996 19014 13006 19066
rect 13006 19014 13052 19066
rect 13076 19014 13122 19066
rect 13122 19014 13132 19066
rect 13156 19014 13186 19066
rect 13186 19014 13212 19066
rect 12916 19012 12972 19014
rect 12996 19012 13052 19014
rect 13076 19012 13132 19014
rect 13156 19012 13212 19014
rect 12916 17978 12972 17980
rect 12996 17978 13052 17980
rect 13076 17978 13132 17980
rect 13156 17978 13212 17980
rect 12916 17926 12942 17978
rect 12942 17926 12972 17978
rect 12996 17926 13006 17978
rect 13006 17926 13052 17978
rect 13076 17926 13122 17978
rect 13122 17926 13132 17978
rect 13156 17926 13186 17978
rect 13186 17926 13212 17978
rect 12916 17924 12972 17926
rect 12996 17924 13052 17926
rect 13076 17924 13132 17926
rect 13156 17924 13212 17926
rect 12916 16890 12972 16892
rect 12996 16890 13052 16892
rect 13076 16890 13132 16892
rect 13156 16890 13212 16892
rect 12916 16838 12942 16890
rect 12942 16838 12972 16890
rect 12996 16838 13006 16890
rect 13006 16838 13052 16890
rect 13076 16838 13122 16890
rect 13122 16838 13132 16890
rect 13156 16838 13186 16890
rect 13186 16838 13212 16890
rect 12916 16836 12972 16838
rect 12996 16836 13052 16838
rect 13076 16836 13132 16838
rect 13156 16836 13212 16838
rect 12916 15802 12972 15804
rect 12996 15802 13052 15804
rect 13076 15802 13132 15804
rect 13156 15802 13212 15804
rect 12916 15750 12942 15802
rect 12942 15750 12972 15802
rect 12996 15750 13006 15802
rect 13006 15750 13052 15802
rect 13076 15750 13122 15802
rect 13122 15750 13132 15802
rect 13156 15750 13186 15802
rect 13186 15750 13212 15802
rect 12916 15748 12972 15750
rect 12996 15748 13052 15750
rect 13076 15748 13132 15750
rect 13156 15748 13212 15750
rect 12916 14714 12972 14716
rect 12996 14714 13052 14716
rect 13076 14714 13132 14716
rect 13156 14714 13212 14716
rect 12916 14662 12942 14714
rect 12942 14662 12972 14714
rect 12996 14662 13006 14714
rect 13006 14662 13052 14714
rect 13076 14662 13122 14714
rect 13122 14662 13132 14714
rect 13156 14662 13186 14714
rect 13186 14662 13212 14714
rect 12916 14660 12972 14662
rect 12996 14660 13052 14662
rect 13076 14660 13132 14662
rect 13156 14660 13212 14662
rect 12916 13626 12972 13628
rect 12996 13626 13052 13628
rect 13076 13626 13132 13628
rect 13156 13626 13212 13628
rect 12916 13574 12942 13626
rect 12942 13574 12972 13626
rect 12996 13574 13006 13626
rect 13006 13574 13052 13626
rect 13076 13574 13122 13626
rect 13122 13574 13132 13626
rect 13156 13574 13186 13626
rect 13186 13574 13212 13626
rect 12916 13572 12972 13574
rect 12996 13572 13052 13574
rect 13076 13572 13132 13574
rect 13156 13572 13212 13574
rect 12916 12538 12972 12540
rect 12996 12538 13052 12540
rect 13076 12538 13132 12540
rect 13156 12538 13212 12540
rect 12916 12486 12942 12538
rect 12942 12486 12972 12538
rect 12996 12486 13006 12538
rect 13006 12486 13052 12538
rect 13076 12486 13122 12538
rect 13122 12486 13132 12538
rect 13156 12486 13186 12538
rect 13186 12486 13212 12538
rect 12916 12484 12972 12486
rect 12996 12484 13052 12486
rect 13076 12484 13132 12486
rect 13156 12484 13212 12486
rect 12916 11450 12972 11452
rect 12996 11450 13052 11452
rect 13076 11450 13132 11452
rect 13156 11450 13212 11452
rect 12916 11398 12942 11450
rect 12942 11398 12972 11450
rect 12996 11398 13006 11450
rect 13006 11398 13052 11450
rect 13076 11398 13122 11450
rect 13122 11398 13132 11450
rect 13156 11398 13186 11450
rect 13186 11398 13212 11450
rect 12916 11396 12972 11398
rect 12996 11396 13052 11398
rect 13076 11396 13132 11398
rect 13156 11396 13212 11398
rect 12916 10362 12972 10364
rect 12996 10362 13052 10364
rect 13076 10362 13132 10364
rect 13156 10362 13212 10364
rect 12916 10310 12942 10362
rect 12942 10310 12972 10362
rect 12996 10310 13006 10362
rect 13006 10310 13052 10362
rect 13076 10310 13122 10362
rect 13122 10310 13132 10362
rect 13156 10310 13186 10362
rect 13186 10310 13212 10362
rect 12916 10308 12972 10310
rect 12996 10308 13052 10310
rect 13076 10308 13132 10310
rect 13156 10308 13212 10310
rect 15906 19610 15962 19612
rect 15986 19610 16042 19612
rect 16066 19610 16122 19612
rect 16146 19610 16202 19612
rect 15906 19558 15932 19610
rect 15932 19558 15962 19610
rect 15986 19558 15996 19610
rect 15996 19558 16042 19610
rect 16066 19558 16112 19610
rect 16112 19558 16122 19610
rect 16146 19558 16176 19610
rect 16176 19558 16202 19610
rect 15906 19556 15962 19558
rect 15986 19556 16042 19558
rect 16066 19556 16122 19558
rect 16146 19556 16202 19558
rect 15382 17040 15438 17096
rect 15906 18522 15962 18524
rect 15986 18522 16042 18524
rect 16066 18522 16122 18524
rect 16146 18522 16202 18524
rect 15906 18470 15932 18522
rect 15932 18470 15962 18522
rect 15986 18470 15996 18522
rect 15996 18470 16042 18522
rect 16066 18470 16112 18522
rect 16112 18470 16122 18522
rect 16146 18470 16176 18522
rect 16176 18470 16202 18522
rect 15906 18468 15962 18470
rect 15986 18468 16042 18470
rect 16066 18468 16122 18470
rect 16146 18468 16202 18470
rect 15906 17434 15962 17436
rect 15986 17434 16042 17436
rect 16066 17434 16122 17436
rect 16146 17434 16202 17436
rect 15906 17382 15932 17434
rect 15932 17382 15962 17434
rect 15986 17382 15996 17434
rect 15996 17382 16042 17434
rect 16066 17382 16112 17434
rect 16112 17382 16122 17434
rect 16146 17382 16176 17434
rect 16176 17382 16202 17434
rect 15906 17380 15962 17382
rect 15986 17380 16042 17382
rect 16066 17380 16122 17382
rect 16146 17380 16202 17382
rect 15906 16346 15962 16348
rect 15986 16346 16042 16348
rect 16066 16346 16122 16348
rect 16146 16346 16202 16348
rect 15906 16294 15932 16346
rect 15932 16294 15962 16346
rect 15986 16294 15996 16346
rect 15996 16294 16042 16346
rect 16066 16294 16112 16346
rect 16112 16294 16122 16346
rect 16146 16294 16176 16346
rect 16176 16294 16202 16346
rect 15906 16292 15962 16294
rect 15986 16292 16042 16294
rect 16066 16292 16122 16294
rect 16146 16292 16202 16294
rect 16210 15680 16266 15736
rect 15906 15258 15962 15260
rect 15986 15258 16042 15260
rect 16066 15258 16122 15260
rect 16146 15258 16202 15260
rect 15906 15206 15932 15258
rect 15932 15206 15962 15258
rect 15986 15206 15996 15258
rect 15996 15206 16042 15258
rect 16066 15206 16112 15258
rect 16112 15206 16122 15258
rect 16146 15206 16176 15258
rect 16176 15206 16202 15258
rect 15906 15204 15962 15206
rect 15986 15204 16042 15206
rect 16066 15204 16122 15206
rect 16146 15204 16202 15206
rect 15906 14170 15962 14172
rect 15986 14170 16042 14172
rect 16066 14170 16122 14172
rect 16146 14170 16202 14172
rect 15906 14118 15932 14170
rect 15932 14118 15962 14170
rect 15986 14118 15996 14170
rect 15996 14118 16042 14170
rect 16066 14118 16112 14170
rect 16112 14118 16122 14170
rect 16146 14118 16176 14170
rect 16176 14118 16202 14170
rect 15906 14116 15962 14118
rect 15986 14116 16042 14118
rect 16066 14116 16122 14118
rect 16146 14116 16202 14118
rect 15906 13082 15962 13084
rect 15986 13082 16042 13084
rect 16066 13082 16122 13084
rect 16146 13082 16202 13084
rect 15906 13030 15932 13082
rect 15932 13030 15962 13082
rect 15986 13030 15996 13082
rect 15996 13030 16042 13082
rect 16066 13030 16112 13082
rect 16112 13030 16122 13082
rect 16146 13030 16176 13082
rect 16176 13030 16202 13082
rect 15906 13028 15962 13030
rect 15986 13028 16042 13030
rect 16066 13028 16122 13030
rect 16146 13028 16202 13030
rect 15906 11994 15962 11996
rect 15986 11994 16042 11996
rect 16066 11994 16122 11996
rect 16146 11994 16202 11996
rect 15906 11942 15932 11994
rect 15932 11942 15962 11994
rect 15986 11942 15996 11994
rect 15996 11942 16042 11994
rect 16066 11942 16112 11994
rect 16112 11942 16122 11994
rect 16146 11942 16176 11994
rect 16176 11942 16202 11994
rect 15906 11940 15962 11942
rect 15986 11940 16042 11942
rect 16066 11940 16122 11942
rect 16146 11940 16202 11942
rect 12916 9274 12972 9276
rect 12996 9274 13052 9276
rect 13076 9274 13132 9276
rect 13156 9274 13212 9276
rect 12916 9222 12942 9274
rect 12942 9222 12972 9274
rect 12996 9222 13006 9274
rect 13006 9222 13052 9274
rect 13076 9222 13122 9274
rect 13122 9222 13132 9274
rect 13156 9222 13186 9274
rect 13186 9222 13212 9274
rect 12916 9220 12972 9222
rect 12996 9220 13052 9222
rect 13076 9220 13132 9222
rect 13156 9220 13212 9222
rect 12916 8186 12972 8188
rect 12996 8186 13052 8188
rect 13076 8186 13132 8188
rect 13156 8186 13212 8188
rect 12916 8134 12942 8186
rect 12942 8134 12972 8186
rect 12996 8134 13006 8186
rect 13006 8134 13052 8186
rect 13076 8134 13122 8186
rect 13122 8134 13132 8186
rect 13156 8134 13186 8186
rect 13186 8134 13212 8186
rect 12916 8132 12972 8134
rect 12996 8132 13052 8134
rect 13076 8132 13132 8134
rect 13156 8132 13212 8134
rect 12916 7098 12972 7100
rect 12996 7098 13052 7100
rect 13076 7098 13132 7100
rect 13156 7098 13212 7100
rect 12916 7046 12942 7098
rect 12942 7046 12972 7098
rect 12996 7046 13006 7098
rect 13006 7046 13052 7098
rect 13076 7046 13122 7098
rect 13122 7046 13132 7098
rect 13156 7046 13186 7098
rect 13186 7046 13212 7098
rect 12916 7044 12972 7046
rect 12996 7044 13052 7046
rect 13076 7044 13132 7046
rect 13156 7044 13212 7046
rect 12916 6010 12972 6012
rect 12996 6010 13052 6012
rect 13076 6010 13132 6012
rect 13156 6010 13212 6012
rect 12916 5958 12942 6010
rect 12942 5958 12972 6010
rect 12996 5958 13006 6010
rect 13006 5958 13052 6010
rect 13076 5958 13122 6010
rect 13122 5958 13132 6010
rect 13156 5958 13186 6010
rect 13186 5958 13212 6010
rect 12916 5956 12972 5958
rect 12996 5956 13052 5958
rect 13076 5956 13132 5958
rect 13156 5956 13212 5958
rect 15906 10906 15962 10908
rect 15986 10906 16042 10908
rect 16066 10906 16122 10908
rect 16146 10906 16202 10908
rect 15906 10854 15932 10906
rect 15932 10854 15962 10906
rect 15986 10854 15996 10906
rect 15996 10854 16042 10906
rect 16066 10854 16112 10906
rect 16112 10854 16122 10906
rect 16146 10854 16176 10906
rect 16176 10854 16202 10906
rect 15906 10852 15962 10854
rect 15986 10852 16042 10854
rect 16066 10852 16122 10854
rect 16146 10852 16202 10854
rect 17866 13640 17922 13696
rect 15906 9818 15962 9820
rect 15986 9818 16042 9820
rect 16066 9818 16122 9820
rect 16146 9818 16202 9820
rect 15906 9766 15932 9818
rect 15932 9766 15962 9818
rect 15986 9766 15996 9818
rect 15996 9766 16042 9818
rect 16066 9766 16112 9818
rect 16112 9766 16122 9818
rect 16146 9766 16176 9818
rect 16176 9766 16202 9818
rect 15906 9764 15962 9766
rect 15986 9764 16042 9766
rect 16066 9764 16122 9766
rect 16146 9764 16202 9766
rect 15906 8730 15962 8732
rect 15986 8730 16042 8732
rect 16066 8730 16122 8732
rect 16146 8730 16202 8732
rect 15906 8678 15932 8730
rect 15932 8678 15962 8730
rect 15986 8678 15996 8730
rect 15996 8678 16042 8730
rect 16066 8678 16112 8730
rect 16112 8678 16122 8730
rect 16146 8678 16176 8730
rect 16176 8678 16202 8730
rect 15906 8676 15962 8678
rect 15986 8676 16042 8678
rect 16066 8676 16122 8678
rect 16146 8676 16202 8678
rect 15906 7642 15962 7644
rect 15986 7642 16042 7644
rect 16066 7642 16122 7644
rect 16146 7642 16202 7644
rect 15906 7590 15932 7642
rect 15932 7590 15962 7642
rect 15986 7590 15996 7642
rect 15996 7590 16042 7642
rect 16066 7590 16112 7642
rect 16112 7590 16122 7642
rect 16146 7590 16176 7642
rect 16176 7590 16202 7642
rect 15906 7588 15962 7590
rect 15986 7588 16042 7590
rect 16066 7588 16122 7590
rect 16146 7588 16202 7590
rect 15906 6554 15962 6556
rect 15986 6554 16042 6556
rect 16066 6554 16122 6556
rect 16146 6554 16202 6556
rect 15906 6502 15932 6554
rect 15932 6502 15962 6554
rect 15986 6502 15996 6554
rect 15996 6502 16042 6554
rect 16066 6502 16112 6554
rect 16112 6502 16122 6554
rect 16146 6502 16176 6554
rect 16176 6502 16202 6554
rect 15906 6500 15962 6502
rect 15986 6500 16042 6502
rect 16066 6500 16122 6502
rect 16146 6500 16202 6502
rect 15906 5466 15962 5468
rect 15986 5466 16042 5468
rect 16066 5466 16122 5468
rect 16146 5466 16202 5468
rect 15906 5414 15932 5466
rect 15932 5414 15962 5466
rect 15986 5414 15996 5466
rect 15996 5414 16042 5466
rect 16066 5414 16112 5466
rect 16112 5414 16122 5466
rect 16146 5414 16176 5466
rect 16176 5414 16202 5466
rect 15906 5412 15962 5414
rect 15986 5412 16042 5414
rect 16066 5412 16122 5414
rect 16146 5412 16202 5414
rect 12916 4922 12972 4924
rect 12996 4922 13052 4924
rect 13076 4922 13132 4924
rect 13156 4922 13212 4924
rect 12916 4870 12942 4922
rect 12942 4870 12972 4922
rect 12996 4870 13006 4922
rect 13006 4870 13052 4922
rect 13076 4870 13122 4922
rect 13122 4870 13132 4922
rect 13156 4870 13186 4922
rect 13186 4870 13212 4922
rect 12916 4868 12972 4870
rect 12996 4868 13052 4870
rect 13076 4868 13132 4870
rect 13156 4868 13212 4870
rect 12916 3834 12972 3836
rect 12996 3834 13052 3836
rect 13076 3834 13132 3836
rect 13156 3834 13212 3836
rect 12916 3782 12942 3834
rect 12942 3782 12972 3834
rect 12996 3782 13006 3834
rect 13006 3782 13052 3834
rect 13076 3782 13122 3834
rect 13122 3782 13132 3834
rect 13156 3782 13186 3834
rect 13186 3782 13212 3834
rect 12916 3780 12972 3782
rect 12996 3780 13052 3782
rect 13076 3780 13132 3782
rect 13156 3780 13212 3782
rect 12916 2746 12972 2748
rect 12996 2746 13052 2748
rect 13076 2746 13132 2748
rect 13156 2746 13212 2748
rect 12916 2694 12942 2746
rect 12942 2694 12972 2746
rect 12996 2694 13006 2746
rect 13006 2694 13052 2746
rect 13076 2694 13122 2746
rect 13122 2694 13132 2746
rect 13156 2694 13186 2746
rect 13186 2694 13212 2746
rect 12916 2692 12972 2694
rect 12996 2692 13052 2694
rect 13076 2692 13132 2694
rect 13156 2692 13212 2694
rect 15906 4378 15962 4380
rect 15986 4378 16042 4380
rect 16066 4378 16122 4380
rect 16146 4378 16202 4380
rect 15906 4326 15932 4378
rect 15932 4326 15962 4378
rect 15986 4326 15996 4378
rect 15996 4326 16042 4378
rect 16066 4326 16112 4378
rect 16112 4326 16122 4378
rect 16146 4326 16176 4378
rect 16176 4326 16202 4378
rect 15906 4324 15962 4326
rect 15986 4324 16042 4326
rect 16066 4324 16122 4326
rect 16146 4324 16202 4326
rect 15906 3290 15962 3292
rect 15986 3290 16042 3292
rect 16066 3290 16122 3292
rect 16146 3290 16202 3292
rect 15906 3238 15932 3290
rect 15932 3238 15962 3290
rect 15986 3238 15996 3290
rect 15996 3238 16042 3290
rect 16066 3238 16112 3290
rect 16112 3238 16122 3290
rect 16146 3238 16176 3290
rect 16176 3238 16202 3290
rect 15906 3236 15962 3238
rect 15986 3236 16042 3238
rect 16066 3236 16122 3238
rect 16146 3236 16202 3238
rect 18326 18400 18382 18456
rect 18326 11600 18382 11656
rect 18326 9560 18382 9616
rect 18326 6860 18382 6896
rect 18326 6840 18328 6860
rect 18328 6840 18380 6860
rect 18380 6840 18382 6860
rect 18326 4800 18382 4856
rect 15906 2202 15962 2204
rect 15986 2202 16042 2204
rect 16066 2202 16122 2204
rect 16146 2202 16202 2204
rect 15906 2150 15932 2202
rect 15932 2150 15962 2202
rect 15986 2150 15996 2202
rect 15996 2150 16042 2202
rect 16066 2150 16112 2202
rect 16112 2150 16122 2202
rect 16146 2150 16176 2202
rect 16176 2150 16202 2202
rect 15906 2148 15962 2150
rect 15986 2148 16042 2150
rect 16066 2148 16122 2150
rect 16146 2148 16202 2150
rect 18326 2760 18382 2816
rect 18418 720 18474 776
<< metal3 >>
rect 0 20498 800 20528
rect 1485 20498 1551 20501
rect 0 20496 1551 20498
rect 0 20440 1490 20496
rect 1546 20440 1551 20496
rect 0 20438 1551 20440
rect 0 20408 800 20438
rect 1485 20435 1551 20438
rect 16481 20498 16547 20501
rect 19396 20498 20196 20528
rect 16481 20496 20196 20498
rect 16481 20440 16486 20496
rect 16542 20440 20196 20496
rect 16481 20438 20196 20440
rect 16481 20435 16547 20438
rect 19396 20408 20196 20438
rect 6924 20160 7244 20161
rect 6924 20096 6932 20160
rect 6996 20096 7012 20160
rect 7076 20096 7092 20160
rect 7156 20096 7172 20160
rect 7236 20096 7244 20160
rect 6924 20095 7244 20096
rect 12904 20160 13224 20161
rect 12904 20096 12912 20160
rect 12976 20096 12992 20160
rect 13056 20096 13072 20160
rect 13136 20096 13152 20160
rect 13216 20096 13224 20160
rect 12904 20095 13224 20096
rect 3934 19616 4254 19617
rect 3934 19552 3942 19616
rect 4006 19552 4022 19616
rect 4086 19552 4102 19616
rect 4166 19552 4182 19616
rect 4246 19552 4254 19616
rect 3934 19551 4254 19552
rect 9914 19616 10234 19617
rect 9914 19552 9922 19616
rect 9986 19552 10002 19616
rect 10066 19552 10082 19616
rect 10146 19552 10162 19616
rect 10226 19552 10234 19616
rect 9914 19551 10234 19552
rect 15894 19616 16214 19617
rect 15894 19552 15902 19616
rect 15966 19552 15982 19616
rect 16046 19552 16062 19616
rect 16126 19552 16142 19616
rect 16206 19552 16214 19616
rect 15894 19551 16214 19552
rect 6924 19072 7244 19073
rect 6924 19008 6932 19072
rect 6996 19008 7012 19072
rect 7076 19008 7092 19072
rect 7156 19008 7172 19072
rect 7236 19008 7244 19072
rect 6924 19007 7244 19008
rect 12904 19072 13224 19073
rect 12904 19008 12912 19072
rect 12976 19008 12992 19072
rect 13056 19008 13072 19072
rect 13136 19008 13152 19072
rect 13216 19008 13224 19072
rect 12904 19007 13224 19008
rect 3934 18528 4254 18529
rect 3934 18464 3942 18528
rect 4006 18464 4022 18528
rect 4086 18464 4102 18528
rect 4166 18464 4182 18528
rect 4246 18464 4254 18528
rect 3934 18463 4254 18464
rect 9914 18528 10234 18529
rect 9914 18464 9922 18528
rect 9986 18464 10002 18528
rect 10066 18464 10082 18528
rect 10146 18464 10162 18528
rect 10226 18464 10234 18528
rect 9914 18463 10234 18464
rect 15894 18528 16214 18529
rect 15894 18464 15902 18528
rect 15966 18464 15982 18528
rect 16046 18464 16062 18528
rect 16126 18464 16142 18528
rect 16206 18464 16214 18528
rect 15894 18463 16214 18464
rect 18321 18458 18387 18461
rect 19396 18458 20196 18488
rect 18321 18456 20196 18458
rect 18321 18400 18326 18456
rect 18382 18400 20196 18456
rect 18321 18398 20196 18400
rect 18321 18395 18387 18398
rect 19396 18368 20196 18398
rect 6924 17984 7244 17985
rect 6924 17920 6932 17984
rect 6996 17920 7012 17984
rect 7076 17920 7092 17984
rect 7156 17920 7172 17984
rect 7236 17920 7244 17984
rect 6924 17919 7244 17920
rect 12904 17984 13224 17985
rect 12904 17920 12912 17984
rect 12976 17920 12992 17984
rect 13056 17920 13072 17984
rect 13136 17920 13152 17984
rect 13216 17920 13224 17984
rect 12904 17919 13224 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 3934 17440 4254 17441
rect 3934 17376 3942 17440
rect 4006 17376 4022 17440
rect 4086 17376 4102 17440
rect 4166 17376 4182 17440
rect 4246 17376 4254 17440
rect 3934 17375 4254 17376
rect 9914 17440 10234 17441
rect 9914 17376 9922 17440
rect 9986 17376 10002 17440
rect 10066 17376 10082 17440
rect 10146 17376 10162 17440
rect 10226 17376 10234 17440
rect 9914 17375 10234 17376
rect 15894 17440 16214 17441
rect 15894 17376 15902 17440
rect 15966 17376 15982 17440
rect 16046 17376 16062 17440
rect 16126 17376 16142 17440
rect 16206 17376 16214 17440
rect 15894 17375 16214 17376
rect 10777 17098 10843 17101
rect 15377 17098 15443 17101
rect 10777 17096 15443 17098
rect 10777 17040 10782 17096
rect 10838 17040 15382 17096
rect 15438 17040 15443 17096
rect 10777 17038 15443 17040
rect 10777 17035 10843 17038
rect 15377 17035 15443 17038
rect 6924 16896 7244 16897
rect 6924 16832 6932 16896
rect 6996 16832 7012 16896
rect 7076 16832 7092 16896
rect 7156 16832 7172 16896
rect 7236 16832 7244 16896
rect 6924 16831 7244 16832
rect 12904 16896 13224 16897
rect 12904 16832 12912 16896
rect 12976 16832 12992 16896
rect 13056 16832 13072 16896
rect 13136 16832 13152 16896
rect 13216 16832 13224 16896
rect 12904 16831 13224 16832
rect 3934 16352 4254 16353
rect 3934 16288 3942 16352
rect 4006 16288 4022 16352
rect 4086 16288 4102 16352
rect 4166 16288 4182 16352
rect 4246 16288 4254 16352
rect 3934 16287 4254 16288
rect 9914 16352 10234 16353
rect 9914 16288 9922 16352
rect 9986 16288 10002 16352
rect 10066 16288 10082 16352
rect 10146 16288 10162 16352
rect 10226 16288 10234 16352
rect 9914 16287 10234 16288
rect 15894 16352 16214 16353
rect 15894 16288 15902 16352
rect 15966 16288 15982 16352
rect 16046 16288 16062 16352
rect 16126 16288 16142 16352
rect 16206 16288 16214 16352
rect 15894 16287 16214 16288
rect 6924 15808 7244 15809
rect 0 15738 800 15768
rect 6924 15744 6932 15808
rect 6996 15744 7012 15808
rect 7076 15744 7092 15808
rect 7156 15744 7172 15808
rect 7236 15744 7244 15808
rect 6924 15743 7244 15744
rect 12904 15808 13224 15809
rect 12904 15744 12912 15808
rect 12976 15744 12992 15808
rect 13056 15744 13072 15808
rect 13136 15744 13152 15808
rect 13216 15744 13224 15808
rect 12904 15743 13224 15744
rect 1393 15738 1459 15741
rect 0 15736 1459 15738
rect 0 15680 1398 15736
rect 1454 15680 1459 15736
rect 0 15678 1459 15680
rect 0 15648 800 15678
rect 1393 15675 1459 15678
rect 16205 15738 16271 15741
rect 19396 15738 20196 15768
rect 16205 15736 20196 15738
rect 16205 15680 16210 15736
rect 16266 15680 20196 15736
rect 16205 15678 20196 15680
rect 16205 15675 16271 15678
rect 19396 15648 20196 15678
rect 3934 15264 4254 15265
rect 3934 15200 3942 15264
rect 4006 15200 4022 15264
rect 4086 15200 4102 15264
rect 4166 15200 4182 15264
rect 4246 15200 4254 15264
rect 3934 15199 4254 15200
rect 9914 15264 10234 15265
rect 9914 15200 9922 15264
rect 9986 15200 10002 15264
rect 10066 15200 10082 15264
rect 10146 15200 10162 15264
rect 10226 15200 10234 15264
rect 9914 15199 10234 15200
rect 15894 15264 16214 15265
rect 15894 15200 15902 15264
rect 15966 15200 15982 15264
rect 16046 15200 16062 15264
rect 16126 15200 16142 15264
rect 16206 15200 16214 15264
rect 15894 15199 16214 15200
rect 6924 14720 7244 14721
rect 6924 14656 6932 14720
rect 6996 14656 7012 14720
rect 7076 14656 7092 14720
rect 7156 14656 7172 14720
rect 7236 14656 7244 14720
rect 6924 14655 7244 14656
rect 12904 14720 13224 14721
rect 12904 14656 12912 14720
rect 12976 14656 12992 14720
rect 13056 14656 13072 14720
rect 13136 14656 13152 14720
rect 13216 14656 13224 14720
rect 12904 14655 13224 14656
rect 3934 14176 4254 14177
rect 3934 14112 3942 14176
rect 4006 14112 4022 14176
rect 4086 14112 4102 14176
rect 4166 14112 4182 14176
rect 4246 14112 4254 14176
rect 3934 14111 4254 14112
rect 9914 14176 10234 14177
rect 9914 14112 9922 14176
rect 9986 14112 10002 14176
rect 10066 14112 10082 14176
rect 10146 14112 10162 14176
rect 10226 14112 10234 14176
rect 9914 14111 10234 14112
rect 15894 14176 16214 14177
rect 15894 14112 15902 14176
rect 15966 14112 15982 14176
rect 16046 14112 16062 14176
rect 16126 14112 16142 14176
rect 16206 14112 16214 14176
rect 15894 14111 16214 14112
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 17861 13698 17927 13701
rect 19396 13698 20196 13728
rect 17861 13696 20196 13698
rect 17861 13640 17866 13696
rect 17922 13640 20196 13696
rect 17861 13638 20196 13640
rect 17861 13635 17927 13638
rect 6924 13632 7244 13633
rect 6924 13568 6932 13632
rect 6996 13568 7012 13632
rect 7076 13568 7092 13632
rect 7156 13568 7172 13632
rect 7236 13568 7244 13632
rect 6924 13567 7244 13568
rect 12904 13632 13224 13633
rect 12904 13568 12912 13632
rect 12976 13568 12992 13632
rect 13056 13568 13072 13632
rect 13136 13568 13152 13632
rect 13216 13568 13224 13632
rect 19396 13608 20196 13638
rect 12904 13567 13224 13568
rect 3934 13088 4254 13089
rect 3934 13024 3942 13088
rect 4006 13024 4022 13088
rect 4086 13024 4102 13088
rect 4166 13024 4182 13088
rect 4246 13024 4254 13088
rect 3934 13023 4254 13024
rect 9914 13088 10234 13089
rect 9914 13024 9922 13088
rect 9986 13024 10002 13088
rect 10066 13024 10082 13088
rect 10146 13024 10162 13088
rect 10226 13024 10234 13088
rect 9914 13023 10234 13024
rect 15894 13088 16214 13089
rect 15894 13024 15902 13088
rect 15966 13024 15982 13088
rect 16046 13024 16062 13088
rect 16126 13024 16142 13088
rect 16206 13024 16214 13088
rect 15894 13023 16214 13024
rect 6924 12544 7244 12545
rect 6924 12480 6932 12544
rect 6996 12480 7012 12544
rect 7076 12480 7092 12544
rect 7156 12480 7172 12544
rect 7236 12480 7244 12544
rect 6924 12479 7244 12480
rect 12904 12544 13224 12545
rect 12904 12480 12912 12544
rect 12976 12480 12992 12544
rect 13056 12480 13072 12544
rect 13136 12480 13152 12544
rect 13216 12480 13224 12544
rect 12904 12479 13224 12480
rect 3934 12000 4254 12001
rect 3934 11936 3942 12000
rect 4006 11936 4022 12000
rect 4086 11936 4102 12000
rect 4166 11936 4182 12000
rect 4246 11936 4254 12000
rect 3934 11935 4254 11936
rect 9914 12000 10234 12001
rect 9914 11936 9922 12000
rect 9986 11936 10002 12000
rect 10066 11936 10082 12000
rect 10146 11936 10162 12000
rect 10226 11936 10234 12000
rect 9914 11935 10234 11936
rect 15894 12000 16214 12001
rect 15894 11936 15902 12000
rect 15966 11936 15982 12000
rect 16046 11936 16062 12000
rect 16126 11936 16142 12000
rect 16206 11936 16214 12000
rect 15894 11935 16214 11936
rect 0 11658 800 11688
rect 1485 11658 1551 11661
rect 0 11656 1551 11658
rect 0 11600 1490 11656
rect 1546 11600 1551 11656
rect 0 11598 1551 11600
rect 0 11568 800 11598
rect 1485 11595 1551 11598
rect 18321 11658 18387 11661
rect 19396 11658 20196 11688
rect 18321 11656 20196 11658
rect 18321 11600 18326 11656
rect 18382 11600 20196 11656
rect 18321 11598 20196 11600
rect 18321 11595 18387 11598
rect 19396 11568 20196 11598
rect 6924 11456 7244 11457
rect 6924 11392 6932 11456
rect 6996 11392 7012 11456
rect 7076 11392 7092 11456
rect 7156 11392 7172 11456
rect 7236 11392 7244 11456
rect 6924 11391 7244 11392
rect 12904 11456 13224 11457
rect 12904 11392 12912 11456
rect 12976 11392 12992 11456
rect 13056 11392 13072 11456
rect 13136 11392 13152 11456
rect 13216 11392 13224 11456
rect 12904 11391 13224 11392
rect 3934 10912 4254 10913
rect 3934 10848 3942 10912
rect 4006 10848 4022 10912
rect 4086 10848 4102 10912
rect 4166 10848 4182 10912
rect 4246 10848 4254 10912
rect 3934 10847 4254 10848
rect 9914 10912 10234 10913
rect 9914 10848 9922 10912
rect 9986 10848 10002 10912
rect 10066 10848 10082 10912
rect 10146 10848 10162 10912
rect 10226 10848 10234 10912
rect 9914 10847 10234 10848
rect 15894 10912 16214 10913
rect 15894 10848 15902 10912
rect 15966 10848 15982 10912
rect 16046 10848 16062 10912
rect 16126 10848 16142 10912
rect 16206 10848 16214 10912
rect 15894 10847 16214 10848
rect 6924 10368 7244 10369
rect 6924 10304 6932 10368
rect 6996 10304 7012 10368
rect 7076 10304 7092 10368
rect 7156 10304 7172 10368
rect 7236 10304 7244 10368
rect 6924 10303 7244 10304
rect 12904 10368 13224 10369
rect 12904 10304 12912 10368
rect 12976 10304 12992 10368
rect 13056 10304 13072 10368
rect 13136 10304 13152 10368
rect 13216 10304 13224 10368
rect 12904 10303 13224 10304
rect 3934 9824 4254 9825
rect 3934 9760 3942 9824
rect 4006 9760 4022 9824
rect 4086 9760 4102 9824
rect 4166 9760 4182 9824
rect 4246 9760 4254 9824
rect 3934 9759 4254 9760
rect 9914 9824 10234 9825
rect 9914 9760 9922 9824
rect 9986 9760 10002 9824
rect 10066 9760 10082 9824
rect 10146 9760 10162 9824
rect 10226 9760 10234 9824
rect 9914 9759 10234 9760
rect 15894 9824 16214 9825
rect 15894 9760 15902 9824
rect 15966 9760 15982 9824
rect 16046 9760 16062 9824
rect 16126 9760 16142 9824
rect 16206 9760 16214 9824
rect 15894 9759 16214 9760
rect 18321 9618 18387 9621
rect 19396 9618 20196 9648
rect 18321 9616 20196 9618
rect 18321 9560 18326 9616
rect 18382 9560 20196 9616
rect 18321 9558 20196 9560
rect 18321 9555 18387 9558
rect 19396 9528 20196 9558
rect 6924 9280 7244 9281
rect 6924 9216 6932 9280
rect 6996 9216 7012 9280
rect 7076 9216 7092 9280
rect 7156 9216 7172 9280
rect 7236 9216 7244 9280
rect 6924 9215 7244 9216
rect 12904 9280 13224 9281
rect 12904 9216 12912 9280
rect 12976 9216 12992 9280
rect 13056 9216 13072 9280
rect 13136 9216 13152 9280
rect 13216 9216 13224 9280
rect 12904 9215 13224 9216
rect 0 8938 800 8968
rect 1393 8938 1459 8941
rect 0 8936 1459 8938
rect 0 8880 1398 8936
rect 1454 8880 1459 8936
rect 0 8878 1459 8880
rect 0 8848 800 8878
rect 1393 8875 1459 8878
rect 3934 8736 4254 8737
rect 3934 8672 3942 8736
rect 4006 8672 4022 8736
rect 4086 8672 4102 8736
rect 4166 8672 4182 8736
rect 4246 8672 4254 8736
rect 3934 8671 4254 8672
rect 9914 8736 10234 8737
rect 9914 8672 9922 8736
rect 9986 8672 10002 8736
rect 10066 8672 10082 8736
rect 10146 8672 10162 8736
rect 10226 8672 10234 8736
rect 9914 8671 10234 8672
rect 15894 8736 16214 8737
rect 15894 8672 15902 8736
rect 15966 8672 15982 8736
rect 16046 8672 16062 8736
rect 16126 8672 16142 8736
rect 16206 8672 16214 8736
rect 15894 8671 16214 8672
rect 6924 8192 7244 8193
rect 6924 8128 6932 8192
rect 6996 8128 7012 8192
rect 7076 8128 7092 8192
rect 7156 8128 7172 8192
rect 7236 8128 7244 8192
rect 6924 8127 7244 8128
rect 12904 8192 13224 8193
rect 12904 8128 12912 8192
rect 12976 8128 12992 8192
rect 13056 8128 13072 8192
rect 13136 8128 13152 8192
rect 13216 8128 13224 8192
rect 12904 8127 13224 8128
rect 3934 7648 4254 7649
rect 3934 7584 3942 7648
rect 4006 7584 4022 7648
rect 4086 7584 4102 7648
rect 4166 7584 4182 7648
rect 4246 7584 4254 7648
rect 3934 7583 4254 7584
rect 9914 7648 10234 7649
rect 9914 7584 9922 7648
rect 9986 7584 10002 7648
rect 10066 7584 10082 7648
rect 10146 7584 10162 7648
rect 10226 7584 10234 7648
rect 9914 7583 10234 7584
rect 15894 7648 16214 7649
rect 15894 7584 15902 7648
rect 15966 7584 15982 7648
rect 16046 7584 16062 7648
rect 16126 7584 16142 7648
rect 16206 7584 16214 7648
rect 15894 7583 16214 7584
rect 6924 7104 7244 7105
rect 6924 7040 6932 7104
rect 6996 7040 7012 7104
rect 7076 7040 7092 7104
rect 7156 7040 7172 7104
rect 7236 7040 7244 7104
rect 6924 7039 7244 7040
rect 12904 7104 13224 7105
rect 12904 7040 12912 7104
rect 12976 7040 12992 7104
rect 13056 7040 13072 7104
rect 13136 7040 13152 7104
rect 13216 7040 13224 7104
rect 12904 7039 13224 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 18321 6898 18387 6901
rect 19396 6898 20196 6928
rect 18321 6896 20196 6898
rect 18321 6840 18326 6896
rect 18382 6840 20196 6896
rect 18321 6838 20196 6840
rect 18321 6835 18387 6838
rect 19396 6808 20196 6838
rect 3934 6560 4254 6561
rect 3934 6496 3942 6560
rect 4006 6496 4022 6560
rect 4086 6496 4102 6560
rect 4166 6496 4182 6560
rect 4246 6496 4254 6560
rect 3934 6495 4254 6496
rect 9914 6560 10234 6561
rect 9914 6496 9922 6560
rect 9986 6496 10002 6560
rect 10066 6496 10082 6560
rect 10146 6496 10162 6560
rect 10226 6496 10234 6560
rect 9914 6495 10234 6496
rect 15894 6560 16214 6561
rect 15894 6496 15902 6560
rect 15966 6496 15982 6560
rect 16046 6496 16062 6560
rect 16126 6496 16142 6560
rect 16206 6496 16214 6560
rect 15894 6495 16214 6496
rect 6924 6016 7244 6017
rect 6924 5952 6932 6016
rect 6996 5952 7012 6016
rect 7076 5952 7092 6016
rect 7156 5952 7172 6016
rect 7236 5952 7244 6016
rect 6924 5951 7244 5952
rect 12904 6016 13224 6017
rect 12904 5952 12912 6016
rect 12976 5952 12992 6016
rect 13056 5952 13072 6016
rect 13136 5952 13152 6016
rect 13216 5952 13224 6016
rect 12904 5951 13224 5952
rect 3934 5472 4254 5473
rect 3934 5408 3942 5472
rect 4006 5408 4022 5472
rect 4086 5408 4102 5472
rect 4166 5408 4182 5472
rect 4246 5408 4254 5472
rect 3934 5407 4254 5408
rect 9914 5472 10234 5473
rect 9914 5408 9922 5472
rect 9986 5408 10002 5472
rect 10066 5408 10082 5472
rect 10146 5408 10162 5472
rect 10226 5408 10234 5472
rect 9914 5407 10234 5408
rect 15894 5472 16214 5473
rect 15894 5408 15902 5472
rect 15966 5408 15982 5472
rect 16046 5408 16062 5472
rect 16126 5408 16142 5472
rect 16206 5408 16214 5472
rect 15894 5407 16214 5408
rect 6924 4928 7244 4929
rect 0 4858 800 4888
rect 6924 4864 6932 4928
rect 6996 4864 7012 4928
rect 7076 4864 7092 4928
rect 7156 4864 7172 4928
rect 7236 4864 7244 4928
rect 6924 4863 7244 4864
rect 12904 4928 13224 4929
rect 12904 4864 12912 4928
rect 12976 4864 12992 4928
rect 13056 4864 13072 4928
rect 13136 4864 13152 4928
rect 13216 4864 13224 4928
rect 12904 4863 13224 4864
rect 1485 4858 1551 4861
rect 0 4856 1551 4858
rect 0 4800 1490 4856
rect 1546 4800 1551 4856
rect 0 4798 1551 4800
rect 0 4768 800 4798
rect 1485 4795 1551 4798
rect 18321 4858 18387 4861
rect 19396 4858 20196 4888
rect 18321 4856 20196 4858
rect 18321 4800 18326 4856
rect 18382 4800 20196 4856
rect 18321 4798 20196 4800
rect 18321 4795 18387 4798
rect 19396 4768 20196 4798
rect 3934 4384 4254 4385
rect 3934 4320 3942 4384
rect 4006 4320 4022 4384
rect 4086 4320 4102 4384
rect 4166 4320 4182 4384
rect 4246 4320 4254 4384
rect 3934 4319 4254 4320
rect 9914 4384 10234 4385
rect 9914 4320 9922 4384
rect 9986 4320 10002 4384
rect 10066 4320 10082 4384
rect 10146 4320 10162 4384
rect 10226 4320 10234 4384
rect 9914 4319 10234 4320
rect 15894 4384 16214 4385
rect 15894 4320 15902 4384
rect 15966 4320 15982 4384
rect 16046 4320 16062 4384
rect 16126 4320 16142 4384
rect 16206 4320 16214 4384
rect 15894 4319 16214 4320
rect 6924 3840 7244 3841
rect 6924 3776 6932 3840
rect 6996 3776 7012 3840
rect 7076 3776 7092 3840
rect 7156 3776 7172 3840
rect 7236 3776 7244 3840
rect 6924 3775 7244 3776
rect 12904 3840 13224 3841
rect 12904 3776 12912 3840
rect 12976 3776 12992 3840
rect 13056 3776 13072 3840
rect 13136 3776 13152 3840
rect 13216 3776 13224 3840
rect 12904 3775 13224 3776
rect 3934 3296 4254 3297
rect 3934 3232 3942 3296
rect 4006 3232 4022 3296
rect 4086 3232 4102 3296
rect 4166 3232 4182 3296
rect 4246 3232 4254 3296
rect 3934 3231 4254 3232
rect 9914 3296 10234 3297
rect 9914 3232 9922 3296
rect 9986 3232 10002 3296
rect 10066 3232 10082 3296
rect 10146 3232 10162 3296
rect 10226 3232 10234 3296
rect 9914 3231 10234 3232
rect 15894 3296 16214 3297
rect 15894 3232 15902 3296
rect 15966 3232 15982 3296
rect 16046 3232 16062 3296
rect 16126 3232 16142 3296
rect 16206 3232 16214 3296
rect 15894 3231 16214 3232
rect 0 2818 800 2848
rect 1393 2818 1459 2821
rect 0 2816 1459 2818
rect 0 2760 1398 2816
rect 1454 2760 1459 2816
rect 0 2758 1459 2760
rect 0 2728 800 2758
rect 1393 2755 1459 2758
rect 18321 2818 18387 2821
rect 19396 2818 20196 2848
rect 18321 2816 20196 2818
rect 18321 2760 18326 2816
rect 18382 2760 20196 2816
rect 18321 2758 20196 2760
rect 18321 2755 18387 2758
rect 6924 2752 7244 2753
rect 6924 2688 6932 2752
rect 6996 2688 7012 2752
rect 7076 2688 7092 2752
rect 7156 2688 7172 2752
rect 7236 2688 7244 2752
rect 6924 2687 7244 2688
rect 12904 2752 13224 2753
rect 12904 2688 12912 2752
rect 12976 2688 12992 2752
rect 13056 2688 13072 2752
rect 13136 2688 13152 2752
rect 13216 2688 13224 2752
rect 19396 2728 20196 2758
rect 12904 2687 13224 2688
rect 3934 2208 4254 2209
rect 3934 2144 3942 2208
rect 4006 2144 4022 2208
rect 4086 2144 4102 2208
rect 4166 2144 4182 2208
rect 4246 2144 4254 2208
rect 3934 2143 4254 2144
rect 9914 2208 10234 2209
rect 9914 2144 9922 2208
rect 9986 2144 10002 2208
rect 10066 2144 10082 2208
rect 10146 2144 10162 2208
rect 10226 2144 10234 2208
rect 9914 2143 10234 2144
rect 15894 2208 16214 2209
rect 15894 2144 15902 2208
rect 15966 2144 15982 2208
rect 16046 2144 16062 2208
rect 16126 2144 16142 2208
rect 16206 2144 16214 2208
rect 15894 2143 16214 2144
rect 18413 778 18479 781
rect 19396 778 20196 808
rect 18413 776 20196 778
rect 18413 720 18418 776
rect 18474 720 20196 776
rect 18413 718 20196 720
rect 18413 715 18479 718
rect 19396 688 20196 718
<< via3 >>
rect 6932 20156 6996 20160
rect 6932 20100 6936 20156
rect 6936 20100 6992 20156
rect 6992 20100 6996 20156
rect 6932 20096 6996 20100
rect 7012 20156 7076 20160
rect 7012 20100 7016 20156
rect 7016 20100 7072 20156
rect 7072 20100 7076 20156
rect 7012 20096 7076 20100
rect 7092 20156 7156 20160
rect 7092 20100 7096 20156
rect 7096 20100 7152 20156
rect 7152 20100 7156 20156
rect 7092 20096 7156 20100
rect 7172 20156 7236 20160
rect 7172 20100 7176 20156
rect 7176 20100 7232 20156
rect 7232 20100 7236 20156
rect 7172 20096 7236 20100
rect 12912 20156 12976 20160
rect 12912 20100 12916 20156
rect 12916 20100 12972 20156
rect 12972 20100 12976 20156
rect 12912 20096 12976 20100
rect 12992 20156 13056 20160
rect 12992 20100 12996 20156
rect 12996 20100 13052 20156
rect 13052 20100 13056 20156
rect 12992 20096 13056 20100
rect 13072 20156 13136 20160
rect 13072 20100 13076 20156
rect 13076 20100 13132 20156
rect 13132 20100 13136 20156
rect 13072 20096 13136 20100
rect 13152 20156 13216 20160
rect 13152 20100 13156 20156
rect 13156 20100 13212 20156
rect 13212 20100 13216 20156
rect 13152 20096 13216 20100
rect 3942 19612 4006 19616
rect 3942 19556 3946 19612
rect 3946 19556 4002 19612
rect 4002 19556 4006 19612
rect 3942 19552 4006 19556
rect 4022 19612 4086 19616
rect 4022 19556 4026 19612
rect 4026 19556 4082 19612
rect 4082 19556 4086 19612
rect 4022 19552 4086 19556
rect 4102 19612 4166 19616
rect 4102 19556 4106 19612
rect 4106 19556 4162 19612
rect 4162 19556 4166 19612
rect 4102 19552 4166 19556
rect 4182 19612 4246 19616
rect 4182 19556 4186 19612
rect 4186 19556 4242 19612
rect 4242 19556 4246 19612
rect 4182 19552 4246 19556
rect 9922 19612 9986 19616
rect 9922 19556 9926 19612
rect 9926 19556 9982 19612
rect 9982 19556 9986 19612
rect 9922 19552 9986 19556
rect 10002 19612 10066 19616
rect 10002 19556 10006 19612
rect 10006 19556 10062 19612
rect 10062 19556 10066 19612
rect 10002 19552 10066 19556
rect 10082 19612 10146 19616
rect 10082 19556 10086 19612
rect 10086 19556 10142 19612
rect 10142 19556 10146 19612
rect 10082 19552 10146 19556
rect 10162 19612 10226 19616
rect 10162 19556 10166 19612
rect 10166 19556 10222 19612
rect 10222 19556 10226 19612
rect 10162 19552 10226 19556
rect 15902 19612 15966 19616
rect 15902 19556 15906 19612
rect 15906 19556 15962 19612
rect 15962 19556 15966 19612
rect 15902 19552 15966 19556
rect 15982 19612 16046 19616
rect 15982 19556 15986 19612
rect 15986 19556 16042 19612
rect 16042 19556 16046 19612
rect 15982 19552 16046 19556
rect 16062 19612 16126 19616
rect 16062 19556 16066 19612
rect 16066 19556 16122 19612
rect 16122 19556 16126 19612
rect 16062 19552 16126 19556
rect 16142 19612 16206 19616
rect 16142 19556 16146 19612
rect 16146 19556 16202 19612
rect 16202 19556 16206 19612
rect 16142 19552 16206 19556
rect 6932 19068 6996 19072
rect 6932 19012 6936 19068
rect 6936 19012 6992 19068
rect 6992 19012 6996 19068
rect 6932 19008 6996 19012
rect 7012 19068 7076 19072
rect 7012 19012 7016 19068
rect 7016 19012 7072 19068
rect 7072 19012 7076 19068
rect 7012 19008 7076 19012
rect 7092 19068 7156 19072
rect 7092 19012 7096 19068
rect 7096 19012 7152 19068
rect 7152 19012 7156 19068
rect 7092 19008 7156 19012
rect 7172 19068 7236 19072
rect 7172 19012 7176 19068
rect 7176 19012 7232 19068
rect 7232 19012 7236 19068
rect 7172 19008 7236 19012
rect 12912 19068 12976 19072
rect 12912 19012 12916 19068
rect 12916 19012 12972 19068
rect 12972 19012 12976 19068
rect 12912 19008 12976 19012
rect 12992 19068 13056 19072
rect 12992 19012 12996 19068
rect 12996 19012 13052 19068
rect 13052 19012 13056 19068
rect 12992 19008 13056 19012
rect 13072 19068 13136 19072
rect 13072 19012 13076 19068
rect 13076 19012 13132 19068
rect 13132 19012 13136 19068
rect 13072 19008 13136 19012
rect 13152 19068 13216 19072
rect 13152 19012 13156 19068
rect 13156 19012 13212 19068
rect 13212 19012 13216 19068
rect 13152 19008 13216 19012
rect 3942 18524 4006 18528
rect 3942 18468 3946 18524
rect 3946 18468 4002 18524
rect 4002 18468 4006 18524
rect 3942 18464 4006 18468
rect 4022 18524 4086 18528
rect 4022 18468 4026 18524
rect 4026 18468 4082 18524
rect 4082 18468 4086 18524
rect 4022 18464 4086 18468
rect 4102 18524 4166 18528
rect 4102 18468 4106 18524
rect 4106 18468 4162 18524
rect 4162 18468 4166 18524
rect 4102 18464 4166 18468
rect 4182 18524 4246 18528
rect 4182 18468 4186 18524
rect 4186 18468 4242 18524
rect 4242 18468 4246 18524
rect 4182 18464 4246 18468
rect 9922 18524 9986 18528
rect 9922 18468 9926 18524
rect 9926 18468 9982 18524
rect 9982 18468 9986 18524
rect 9922 18464 9986 18468
rect 10002 18524 10066 18528
rect 10002 18468 10006 18524
rect 10006 18468 10062 18524
rect 10062 18468 10066 18524
rect 10002 18464 10066 18468
rect 10082 18524 10146 18528
rect 10082 18468 10086 18524
rect 10086 18468 10142 18524
rect 10142 18468 10146 18524
rect 10082 18464 10146 18468
rect 10162 18524 10226 18528
rect 10162 18468 10166 18524
rect 10166 18468 10222 18524
rect 10222 18468 10226 18524
rect 10162 18464 10226 18468
rect 15902 18524 15966 18528
rect 15902 18468 15906 18524
rect 15906 18468 15962 18524
rect 15962 18468 15966 18524
rect 15902 18464 15966 18468
rect 15982 18524 16046 18528
rect 15982 18468 15986 18524
rect 15986 18468 16042 18524
rect 16042 18468 16046 18524
rect 15982 18464 16046 18468
rect 16062 18524 16126 18528
rect 16062 18468 16066 18524
rect 16066 18468 16122 18524
rect 16122 18468 16126 18524
rect 16062 18464 16126 18468
rect 16142 18524 16206 18528
rect 16142 18468 16146 18524
rect 16146 18468 16202 18524
rect 16202 18468 16206 18524
rect 16142 18464 16206 18468
rect 6932 17980 6996 17984
rect 6932 17924 6936 17980
rect 6936 17924 6992 17980
rect 6992 17924 6996 17980
rect 6932 17920 6996 17924
rect 7012 17980 7076 17984
rect 7012 17924 7016 17980
rect 7016 17924 7072 17980
rect 7072 17924 7076 17980
rect 7012 17920 7076 17924
rect 7092 17980 7156 17984
rect 7092 17924 7096 17980
rect 7096 17924 7152 17980
rect 7152 17924 7156 17980
rect 7092 17920 7156 17924
rect 7172 17980 7236 17984
rect 7172 17924 7176 17980
rect 7176 17924 7232 17980
rect 7232 17924 7236 17980
rect 7172 17920 7236 17924
rect 12912 17980 12976 17984
rect 12912 17924 12916 17980
rect 12916 17924 12972 17980
rect 12972 17924 12976 17980
rect 12912 17920 12976 17924
rect 12992 17980 13056 17984
rect 12992 17924 12996 17980
rect 12996 17924 13052 17980
rect 13052 17924 13056 17980
rect 12992 17920 13056 17924
rect 13072 17980 13136 17984
rect 13072 17924 13076 17980
rect 13076 17924 13132 17980
rect 13132 17924 13136 17980
rect 13072 17920 13136 17924
rect 13152 17980 13216 17984
rect 13152 17924 13156 17980
rect 13156 17924 13212 17980
rect 13212 17924 13216 17980
rect 13152 17920 13216 17924
rect 3942 17436 4006 17440
rect 3942 17380 3946 17436
rect 3946 17380 4002 17436
rect 4002 17380 4006 17436
rect 3942 17376 4006 17380
rect 4022 17436 4086 17440
rect 4022 17380 4026 17436
rect 4026 17380 4082 17436
rect 4082 17380 4086 17436
rect 4022 17376 4086 17380
rect 4102 17436 4166 17440
rect 4102 17380 4106 17436
rect 4106 17380 4162 17436
rect 4162 17380 4166 17436
rect 4102 17376 4166 17380
rect 4182 17436 4246 17440
rect 4182 17380 4186 17436
rect 4186 17380 4242 17436
rect 4242 17380 4246 17436
rect 4182 17376 4246 17380
rect 9922 17436 9986 17440
rect 9922 17380 9926 17436
rect 9926 17380 9982 17436
rect 9982 17380 9986 17436
rect 9922 17376 9986 17380
rect 10002 17436 10066 17440
rect 10002 17380 10006 17436
rect 10006 17380 10062 17436
rect 10062 17380 10066 17436
rect 10002 17376 10066 17380
rect 10082 17436 10146 17440
rect 10082 17380 10086 17436
rect 10086 17380 10142 17436
rect 10142 17380 10146 17436
rect 10082 17376 10146 17380
rect 10162 17436 10226 17440
rect 10162 17380 10166 17436
rect 10166 17380 10222 17436
rect 10222 17380 10226 17436
rect 10162 17376 10226 17380
rect 15902 17436 15966 17440
rect 15902 17380 15906 17436
rect 15906 17380 15962 17436
rect 15962 17380 15966 17436
rect 15902 17376 15966 17380
rect 15982 17436 16046 17440
rect 15982 17380 15986 17436
rect 15986 17380 16042 17436
rect 16042 17380 16046 17436
rect 15982 17376 16046 17380
rect 16062 17436 16126 17440
rect 16062 17380 16066 17436
rect 16066 17380 16122 17436
rect 16122 17380 16126 17436
rect 16062 17376 16126 17380
rect 16142 17436 16206 17440
rect 16142 17380 16146 17436
rect 16146 17380 16202 17436
rect 16202 17380 16206 17436
rect 16142 17376 16206 17380
rect 6932 16892 6996 16896
rect 6932 16836 6936 16892
rect 6936 16836 6992 16892
rect 6992 16836 6996 16892
rect 6932 16832 6996 16836
rect 7012 16892 7076 16896
rect 7012 16836 7016 16892
rect 7016 16836 7072 16892
rect 7072 16836 7076 16892
rect 7012 16832 7076 16836
rect 7092 16892 7156 16896
rect 7092 16836 7096 16892
rect 7096 16836 7152 16892
rect 7152 16836 7156 16892
rect 7092 16832 7156 16836
rect 7172 16892 7236 16896
rect 7172 16836 7176 16892
rect 7176 16836 7232 16892
rect 7232 16836 7236 16892
rect 7172 16832 7236 16836
rect 12912 16892 12976 16896
rect 12912 16836 12916 16892
rect 12916 16836 12972 16892
rect 12972 16836 12976 16892
rect 12912 16832 12976 16836
rect 12992 16892 13056 16896
rect 12992 16836 12996 16892
rect 12996 16836 13052 16892
rect 13052 16836 13056 16892
rect 12992 16832 13056 16836
rect 13072 16892 13136 16896
rect 13072 16836 13076 16892
rect 13076 16836 13132 16892
rect 13132 16836 13136 16892
rect 13072 16832 13136 16836
rect 13152 16892 13216 16896
rect 13152 16836 13156 16892
rect 13156 16836 13212 16892
rect 13212 16836 13216 16892
rect 13152 16832 13216 16836
rect 3942 16348 4006 16352
rect 3942 16292 3946 16348
rect 3946 16292 4002 16348
rect 4002 16292 4006 16348
rect 3942 16288 4006 16292
rect 4022 16348 4086 16352
rect 4022 16292 4026 16348
rect 4026 16292 4082 16348
rect 4082 16292 4086 16348
rect 4022 16288 4086 16292
rect 4102 16348 4166 16352
rect 4102 16292 4106 16348
rect 4106 16292 4162 16348
rect 4162 16292 4166 16348
rect 4102 16288 4166 16292
rect 4182 16348 4246 16352
rect 4182 16292 4186 16348
rect 4186 16292 4242 16348
rect 4242 16292 4246 16348
rect 4182 16288 4246 16292
rect 9922 16348 9986 16352
rect 9922 16292 9926 16348
rect 9926 16292 9982 16348
rect 9982 16292 9986 16348
rect 9922 16288 9986 16292
rect 10002 16348 10066 16352
rect 10002 16292 10006 16348
rect 10006 16292 10062 16348
rect 10062 16292 10066 16348
rect 10002 16288 10066 16292
rect 10082 16348 10146 16352
rect 10082 16292 10086 16348
rect 10086 16292 10142 16348
rect 10142 16292 10146 16348
rect 10082 16288 10146 16292
rect 10162 16348 10226 16352
rect 10162 16292 10166 16348
rect 10166 16292 10222 16348
rect 10222 16292 10226 16348
rect 10162 16288 10226 16292
rect 15902 16348 15966 16352
rect 15902 16292 15906 16348
rect 15906 16292 15962 16348
rect 15962 16292 15966 16348
rect 15902 16288 15966 16292
rect 15982 16348 16046 16352
rect 15982 16292 15986 16348
rect 15986 16292 16042 16348
rect 16042 16292 16046 16348
rect 15982 16288 16046 16292
rect 16062 16348 16126 16352
rect 16062 16292 16066 16348
rect 16066 16292 16122 16348
rect 16122 16292 16126 16348
rect 16062 16288 16126 16292
rect 16142 16348 16206 16352
rect 16142 16292 16146 16348
rect 16146 16292 16202 16348
rect 16202 16292 16206 16348
rect 16142 16288 16206 16292
rect 6932 15804 6996 15808
rect 6932 15748 6936 15804
rect 6936 15748 6992 15804
rect 6992 15748 6996 15804
rect 6932 15744 6996 15748
rect 7012 15804 7076 15808
rect 7012 15748 7016 15804
rect 7016 15748 7072 15804
rect 7072 15748 7076 15804
rect 7012 15744 7076 15748
rect 7092 15804 7156 15808
rect 7092 15748 7096 15804
rect 7096 15748 7152 15804
rect 7152 15748 7156 15804
rect 7092 15744 7156 15748
rect 7172 15804 7236 15808
rect 7172 15748 7176 15804
rect 7176 15748 7232 15804
rect 7232 15748 7236 15804
rect 7172 15744 7236 15748
rect 12912 15804 12976 15808
rect 12912 15748 12916 15804
rect 12916 15748 12972 15804
rect 12972 15748 12976 15804
rect 12912 15744 12976 15748
rect 12992 15804 13056 15808
rect 12992 15748 12996 15804
rect 12996 15748 13052 15804
rect 13052 15748 13056 15804
rect 12992 15744 13056 15748
rect 13072 15804 13136 15808
rect 13072 15748 13076 15804
rect 13076 15748 13132 15804
rect 13132 15748 13136 15804
rect 13072 15744 13136 15748
rect 13152 15804 13216 15808
rect 13152 15748 13156 15804
rect 13156 15748 13212 15804
rect 13212 15748 13216 15804
rect 13152 15744 13216 15748
rect 3942 15260 4006 15264
rect 3942 15204 3946 15260
rect 3946 15204 4002 15260
rect 4002 15204 4006 15260
rect 3942 15200 4006 15204
rect 4022 15260 4086 15264
rect 4022 15204 4026 15260
rect 4026 15204 4082 15260
rect 4082 15204 4086 15260
rect 4022 15200 4086 15204
rect 4102 15260 4166 15264
rect 4102 15204 4106 15260
rect 4106 15204 4162 15260
rect 4162 15204 4166 15260
rect 4102 15200 4166 15204
rect 4182 15260 4246 15264
rect 4182 15204 4186 15260
rect 4186 15204 4242 15260
rect 4242 15204 4246 15260
rect 4182 15200 4246 15204
rect 9922 15260 9986 15264
rect 9922 15204 9926 15260
rect 9926 15204 9982 15260
rect 9982 15204 9986 15260
rect 9922 15200 9986 15204
rect 10002 15260 10066 15264
rect 10002 15204 10006 15260
rect 10006 15204 10062 15260
rect 10062 15204 10066 15260
rect 10002 15200 10066 15204
rect 10082 15260 10146 15264
rect 10082 15204 10086 15260
rect 10086 15204 10142 15260
rect 10142 15204 10146 15260
rect 10082 15200 10146 15204
rect 10162 15260 10226 15264
rect 10162 15204 10166 15260
rect 10166 15204 10222 15260
rect 10222 15204 10226 15260
rect 10162 15200 10226 15204
rect 15902 15260 15966 15264
rect 15902 15204 15906 15260
rect 15906 15204 15962 15260
rect 15962 15204 15966 15260
rect 15902 15200 15966 15204
rect 15982 15260 16046 15264
rect 15982 15204 15986 15260
rect 15986 15204 16042 15260
rect 16042 15204 16046 15260
rect 15982 15200 16046 15204
rect 16062 15260 16126 15264
rect 16062 15204 16066 15260
rect 16066 15204 16122 15260
rect 16122 15204 16126 15260
rect 16062 15200 16126 15204
rect 16142 15260 16206 15264
rect 16142 15204 16146 15260
rect 16146 15204 16202 15260
rect 16202 15204 16206 15260
rect 16142 15200 16206 15204
rect 6932 14716 6996 14720
rect 6932 14660 6936 14716
rect 6936 14660 6992 14716
rect 6992 14660 6996 14716
rect 6932 14656 6996 14660
rect 7012 14716 7076 14720
rect 7012 14660 7016 14716
rect 7016 14660 7072 14716
rect 7072 14660 7076 14716
rect 7012 14656 7076 14660
rect 7092 14716 7156 14720
rect 7092 14660 7096 14716
rect 7096 14660 7152 14716
rect 7152 14660 7156 14716
rect 7092 14656 7156 14660
rect 7172 14716 7236 14720
rect 7172 14660 7176 14716
rect 7176 14660 7232 14716
rect 7232 14660 7236 14716
rect 7172 14656 7236 14660
rect 12912 14716 12976 14720
rect 12912 14660 12916 14716
rect 12916 14660 12972 14716
rect 12972 14660 12976 14716
rect 12912 14656 12976 14660
rect 12992 14716 13056 14720
rect 12992 14660 12996 14716
rect 12996 14660 13052 14716
rect 13052 14660 13056 14716
rect 12992 14656 13056 14660
rect 13072 14716 13136 14720
rect 13072 14660 13076 14716
rect 13076 14660 13132 14716
rect 13132 14660 13136 14716
rect 13072 14656 13136 14660
rect 13152 14716 13216 14720
rect 13152 14660 13156 14716
rect 13156 14660 13212 14716
rect 13212 14660 13216 14716
rect 13152 14656 13216 14660
rect 3942 14172 4006 14176
rect 3942 14116 3946 14172
rect 3946 14116 4002 14172
rect 4002 14116 4006 14172
rect 3942 14112 4006 14116
rect 4022 14172 4086 14176
rect 4022 14116 4026 14172
rect 4026 14116 4082 14172
rect 4082 14116 4086 14172
rect 4022 14112 4086 14116
rect 4102 14172 4166 14176
rect 4102 14116 4106 14172
rect 4106 14116 4162 14172
rect 4162 14116 4166 14172
rect 4102 14112 4166 14116
rect 4182 14172 4246 14176
rect 4182 14116 4186 14172
rect 4186 14116 4242 14172
rect 4242 14116 4246 14172
rect 4182 14112 4246 14116
rect 9922 14172 9986 14176
rect 9922 14116 9926 14172
rect 9926 14116 9982 14172
rect 9982 14116 9986 14172
rect 9922 14112 9986 14116
rect 10002 14172 10066 14176
rect 10002 14116 10006 14172
rect 10006 14116 10062 14172
rect 10062 14116 10066 14172
rect 10002 14112 10066 14116
rect 10082 14172 10146 14176
rect 10082 14116 10086 14172
rect 10086 14116 10142 14172
rect 10142 14116 10146 14172
rect 10082 14112 10146 14116
rect 10162 14172 10226 14176
rect 10162 14116 10166 14172
rect 10166 14116 10222 14172
rect 10222 14116 10226 14172
rect 10162 14112 10226 14116
rect 15902 14172 15966 14176
rect 15902 14116 15906 14172
rect 15906 14116 15962 14172
rect 15962 14116 15966 14172
rect 15902 14112 15966 14116
rect 15982 14172 16046 14176
rect 15982 14116 15986 14172
rect 15986 14116 16042 14172
rect 16042 14116 16046 14172
rect 15982 14112 16046 14116
rect 16062 14172 16126 14176
rect 16062 14116 16066 14172
rect 16066 14116 16122 14172
rect 16122 14116 16126 14172
rect 16062 14112 16126 14116
rect 16142 14172 16206 14176
rect 16142 14116 16146 14172
rect 16146 14116 16202 14172
rect 16202 14116 16206 14172
rect 16142 14112 16206 14116
rect 6932 13628 6996 13632
rect 6932 13572 6936 13628
rect 6936 13572 6992 13628
rect 6992 13572 6996 13628
rect 6932 13568 6996 13572
rect 7012 13628 7076 13632
rect 7012 13572 7016 13628
rect 7016 13572 7072 13628
rect 7072 13572 7076 13628
rect 7012 13568 7076 13572
rect 7092 13628 7156 13632
rect 7092 13572 7096 13628
rect 7096 13572 7152 13628
rect 7152 13572 7156 13628
rect 7092 13568 7156 13572
rect 7172 13628 7236 13632
rect 7172 13572 7176 13628
rect 7176 13572 7232 13628
rect 7232 13572 7236 13628
rect 7172 13568 7236 13572
rect 12912 13628 12976 13632
rect 12912 13572 12916 13628
rect 12916 13572 12972 13628
rect 12972 13572 12976 13628
rect 12912 13568 12976 13572
rect 12992 13628 13056 13632
rect 12992 13572 12996 13628
rect 12996 13572 13052 13628
rect 13052 13572 13056 13628
rect 12992 13568 13056 13572
rect 13072 13628 13136 13632
rect 13072 13572 13076 13628
rect 13076 13572 13132 13628
rect 13132 13572 13136 13628
rect 13072 13568 13136 13572
rect 13152 13628 13216 13632
rect 13152 13572 13156 13628
rect 13156 13572 13212 13628
rect 13212 13572 13216 13628
rect 13152 13568 13216 13572
rect 3942 13084 4006 13088
rect 3942 13028 3946 13084
rect 3946 13028 4002 13084
rect 4002 13028 4006 13084
rect 3942 13024 4006 13028
rect 4022 13084 4086 13088
rect 4022 13028 4026 13084
rect 4026 13028 4082 13084
rect 4082 13028 4086 13084
rect 4022 13024 4086 13028
rect 4102 13084 4166 13088
rect 4102 13028 4106 13084
rect 4106 13028 4162 13084
rect 4162 13028 4166 13084
rect 4102 13024 4166 13028
rect 4182 13084 4246 13088
rect 4182 13028 4186 13084
rect 4186 13028 4242 13084
rect 4242 13028 4246 13084
rect 4182 13024 4246 13028
rect 9922 13084 9986 13088
rect 9922 13028 9926 13084
rect 9926 13028 9982 13084
rect 9982 13028 9986 13084
rect 9922 13024 9986 13028
rect 10002 13084 10066 13088
rect 10002 13028 10006 13084
rect 10006 13028 10062 13084
rect 10062 13028 10066 13084
rect 10002 13024 10066 13028
rect 10082 13084 10146 13088
rect 10082 13028 10086 13084
rect 10086 13028 10142 13084
rect 10142 13028 10146 13084
rect 10082 13024 10146 13028
rect 10162 13084 10226 13088
rect 10162 13028 10166 13084
rect 10166 13028 10222 13084
rect 10222 13028 10226 13084
rect 10162 13024 10226 13028
rect 15902 13084 15966 13088
rect 15902 13028 15906 13084
rect 15906 13028 15962 13084
rect 15962 13028 15966 13084
rect 15902 13024 15966 13028
rect 15982 13084 16046 13088
rect 15982 13028 15986 13084
rect 15986 13028 16042 13084
rect 16042 13028 16046 13084
rect 15982 13024 16046 13028
rect 16062 13084 16126 13088
rect 16062 13028 16066 13084
rect 16066 13028 16122 13084
rect 16122 13028 16126 13084
rect 16062 13024 16126 13028
rect 16142 13084 16206 13088
rect 16142 13028 16146 13084
rect 16146 13028 16202 13084
rect 16202 13028 16206 13084
rect 16142 13024 16206 13028
rect 6932 12540 6996 12544
rect 6932 12484 6936 12540
rect 6936 12484 6992 12540
rect 6992 12484 6996 12540
rect 6932 12480 6996 12484
rect 7012 12540 7076 12544
rect 7012 12484 7016 12540
rect 7016 12484 7072 12540
rect 7072 12484 7076 12540
rect 7012 12480 7076 12484
rect 7092 12540 7156 12544
rect 7092 12484 7096 12540
rect 7096 12484 7152 12540
rect 7152 12484 7156 12540
rect 7092 12480 7156 12484
rect 7172 12540 7236 12544
rect 7172 12484 7176 12540
rect 7176 12484 7232 12540
rect 7232 12484 7236 12540
rect 7172 12480 7236 12484
rect 12912 12540 12976 12544
rect 12912 12484 12916 12540
rect 12916 12484 12972 12540
rect 12972 12484 12976 12540
rect 12912 12480 12976 12484
rect 12992 12540 13056 12544
rect 12992 12484 12996 12540
rect 12996 12484 13052 12540
rect 13052 12484 13056 12540
rect 12992 12480 13056 12484
rect 13072 12540 13136 12544
rect 13072 12484 13076 12540
rect 13076 12484 13132 12540
rect 13132 12484 13136 12540
rect 13072 12480 13136 12484
rect 13152 12540 13216 12544
rect 13152 12484 13156 12540
rect 13156 12484 13212 12540
rect 13212 12484 13216 12540
rect 13152 12480 13216 12484
rect 3942 11996 4006 12000
rect 3942 11940 3946 11996
rect 3946 11940 4002 11996
rect 4002 11940 4006 11996
rect 3942 11936 4006 11940
rect 4022 11996 4086 12000
rect 4022 11940 4026 11996
rect 4026 11940 4082 11996
rect 4082 11940 4086 11996
rect 4022 11936 4086 11940
rect 4102 11996 4166 12000
rect 4102 11940 4106 11996
rect 4106 11940 4162 11996
rect 4162 11940 4166 11996
rect 4102 11936 4166 11940
rect 4182 11996 4246 12000
rect 4182 11940 4186 11996
rect 4186 11940 4242 11996
rect 4242 11940 4246 11996
rect 4182 11936 4246 11940
rect 9922 11996 9986 12000
rect 9922 11940 9926 11996
rect 9926 11940 9982 11996
rect 9982 11940 9986 11996
rect 9922 11936 9986 11940
rect 10002 11996 10066 12000
rect 10002 11940 10006 11996
rect 10006 11940 10062 11996
rect 10062 11940 10066 11996
rect 10002 11936 10066 11940
rect 10082 11996 10146 12000
rect 10082 11940 10086 11996
rect 10086 11940 10142 11996
rect 10142 11940 10146 11996
rect 10082 11936 10146 11940
rect 10162 11996 10226 12000
rect 10162 11940 10166 11996
rect 10166 11940 10222 11996
rect 10222 11940 10226 11996
rect 10162 11936 10226 11940
rect 15902 11996 15966 12000
rect 15902 11940 15906 11996
rect 15906 11940 15962 11996
rect 15962 11940 15966 11996
rect 15902 11936 15966 11940
rect 15982 11996 16046 12000
rect 15982 11940 15986 11996
rect 15986 11940 16042 11996
rect 16042 11940 16046 11996
rect 15982 11936 16046 11940
rect 16062 11996 16126 12000
rect 16062 11940 16066 11996
rect 16066 11940 16122 11996
rect 16122 11940 16126 11996
rect 16062 11936 16126 11940
rect 16142 11996 16206 12000
rect 16142 11940 16146 11996
rect 16146 11940 16202 11996
rect 16202 11940 16206 11996
rect 16142 11936 16206 11940
rect 6932 11452 6996 11456
rect 6932 11396 6936 11452
rect 6936 11396 6992 11452
rect 6992 11396 6996 11452
rect 6932 11392 6996 11396
rect 7012 11452 7076 11456
rect 7012 11396 7016 11452
rect 7016 11396 7072 11452
rect 7072 11396 7076 11452
rect 7012 11392 7076 11396
rect 7092 11452 7156 11456
rect 7092 11396 7096 11452
rect 7096 11396 7152 11452
rect 7152 11396 7156 11452
rect 7092 11392 7156 11396
rect 7172 11452 7236 11456
rect 7172 11396 7176 11452
rect 7176 11396 7232 11452
rect 7232 11396 7236 11452
rect 7172 11392 7236 11396
rect 12912 11452 12976 11456
rect 12912 11396 12916 11452
rect 12916 11396 12972 11452
rect 12972 11396 12976 11452
rect 12912 11392 12976 11396
rect 12992 11452 13056 11456
rect 12992 11396 12996 11452
rect 12996 11396 13052 11452
rect 13052 11396 13056 11452
rect 12992 11392 13056 11396
rect 13072 11452 13136 11456
rect 13072 11396 13076 11452
rect 13076 11396 13132 11452
rect 13132 11396 13136 11452
rect 13072 11392 13136 11396
rect 13152 11452 13216 11456
rect 13152 11396 13156 11452
rect 13156 11396 13212 11452
rect 13212 11396 13216 11452
rect 13152 11392 13216 11396
rect 3942 10908 4006 10912
rect 3942 10852 3946 10908
rect 3946 10852 4002 10908
rect 4002 10852 4006 10908
rect 3942 10848 4006 10852
rect 4022 10908 4086 10912
rect 4022 10852 4026 10908
rect 4026 10852 4082 10908
rect 4082 10852 4086 10908
rect 4022 10848 4086 10852
rect 4102 10908 4166 10912
rect 4102 10852 4106 10908
rect 4106 10852 4162 10908
rect 4162 10852 4166 10908
rect 4102 10848 4166 10852
rect 4182 10908 4246 10912
rect 4182 10852 4186 10908
rect 4186 10852 4242 10908
rect 4242 10852 4246 10908
rect 4182 10848 4246 10852
rect 9922 10908 9986 10912
rect 9922 10852 9926 10908
rect 9926 10852 9982 10908
rect 9982 10852 9986 10908
rect 9922 10848 9986 10852
rect 10002 10908 10066 10912
rect 10002 10852 10006 10908
rect 10006 10852 10062 10908
rect 10062 10852 10066 10908
rect 10002 10848 10066 10852
rect 10082 10908 10146 10912
rect 10082 10852 10086 10908
rect 10086 10852 10142 10908
rect 10142 10852 10146 10908
rect 10082 10848 10146 10852
rect 10162 10908 10226 10912
rect 10162 10852 10166 10908
rect 10166 10852 10222 10908
rect 10222 10852 10226 10908
rect 10162 10848 10226 10852
rect 15902 10908 15966 10912
rect 15902 10852 15906 10908
rect 15906 10852 15962 10908
rect 15962 10852 15966 10908
rect 15902 10848 15966 10852
rect 15982 10908 16046 10912
rect 15982 10852 15986 10908
rect 15986 10852 16042 10908
rect 16042 10852 16046 10908
rect 15982 10848 16046 10852
rect 16062 10908 16126 10912
rect 16062 10852 16066 10908
rect 16066 10852 16122 10908
rect 16122 10852 16126 10908
rect 16062 10848 16126 10852
rect 16142 10908 16206 10912
rect 16142 10852 16146 10908
rect 16146 10852 16202 10908
rect 16202 10852 16206 10908
rect 16142 10848 16206 10852
rect 6932 10364 6996 10368
rect 6932 10308 6936 10364
rect 6936 10308 6992 10364
rect 6992 10308 6996 10364
rect 6932 10304 6996 10308
rect 7012 10364 7076 10368
rect 7012 10308 7016 10364
rect 7016 10308 7072 10364
rect 7072 10308 7076 10364
rect 7012 10304 7076 10308
rect 7092 10364 7156 10368
rect 7092 10308 7096 10364
rect 7096 10308 7152 10364
rect 7152 10308 7156 10364
rect 7092 10304 7156 10308
rect 7172 10364 7236 10368
rect 7172 10308 7176 10364
rect 7176 10308 7232 10364
rect 7232 10308 7236 10364
rect 7172 10304 7236 10308
rect 12912 10364 12976 10368
rect 12912 10308 12916 10364
rect 12916 10308 12972 10364
rect 12972 10308 12976 10364
rect 12912 10304 12976 10308
rect 12992 10364 13056 10368
rect 12992 10308 12996 10364
rect 12996 10308 13052 10364
rect 13052 10308 13056 10364
rect 12992 10304 13056 10308
rect 13072 10364 13136 10368
rect 13072 10308 13076 10364
rect 13076 10308 13132 10364
rect 13132 10308 13136 10364
rect 13072 10304 13136 10308
rect 13152 10364 13216 10368
rect 13152 10308 13156 10364
rect 13156 10308 13212 10364
rect 13212 10308 13216 10364
rect 13152 10304 13216 10308
rect 3942 9820 4006 9824
rect 3942 9764 3946 9820
rect 3946 9764 4002 9820
rect 4002 9764 4006 9820
rect 3942 9760 4006 9764
rect 4022 9820 4086 9824
rect 4022 9764 4026 9820
rect 4026 9764 4082 9820
rect 4082 9764 4086 9820
rect 4022 9760 4086 9764
rect 4102 9820 4166 9824
rect 4102 9764 4106 9820
rect 4106 9764 4162 9820
rect 4162 9764 4166 9820
rect 4102 9760 4166 9764
rect 4182 9820 4246 9824
rect 4182 9764 4186 9820
rect 4186 9764 4242 9820
rect 4242 9764 4246 9820
rect 4182 9760 4246 9764
rect 9922 9820 9986 9824
rect 9922 9764 9926 9820
rect 9926 9764 9982 9820
rect 9982 9764 9986 9820
rect 9922 9760 9986 9764
rect 10002 9820 10066 9824
rect 10002 9764 10006 9820
rect 10006 9764 10062 9820
rect 10062 9764 10066 9820
rect 10002 9760 10066 9764
rect 10082 9820 10146 9824
rect 10082 9764 10086 9820
rect 10086 9764 10142 9820
rect 10142 9764 10146 9820
rect 10082 9760 10146 9764
rect 10162 9820 10226 9824
rect 10162 9764 10166 9820
rect 10166 9764 10222 9820
rect 10222 9764 10226 9820
rect 10162 9760 10226 9764
rect 15902 9820 15966 9824
rect 15902 9764 15906 9820
rect 15906 9764 15962 9820
rect 15962 9764 15966 9820
rect 15902 9760 15966 9764
rect 15982 9820 16046 9824
rect 15982 9764 15986 9820
rect 15986 9764 16042 9820
rect 16042 9764 16046 9820
rect 15982 9760 16046 9764
rect 16062 9820 16126 9824
rect 16062 9764 16066 9820
rect 16066 9764 16122 9820
rect 16122 9764 16126 9820
rect 16062 9760 16126 9764
rect 16142 9820 16206 9824
rect 16142 9764 16146 9820
rect 16146 9764 16202 9820
rect 16202 9764 16206 9820
rect 16142 9760 16206 9764
rect 6932 9276 6996 9280
rect 6932 9220 6936 9276
rect 6936 9220 6992 9276
rect 6992 9220 6996 9276
rect 6932 9216 6996 9220
rect 7012 9276 7076 9280
rect 7012 9220 7016 9276
rect 7016 9220 7072 9276
rect 7072 9220 7076 9276
rect 7012 9216 7076 9220
rect 7092 9276 7156 9280
rect 7092 9220 7096 9276
rect 7096 9220 7152 9276
rect 7152 9220 7156 9276
rect 7092 9216 7156 9220
rect 7172 9276 7236 9280
rect 7172 9220 7176 9276
rect 7176 9220 7232 9276
rect 7232 9220 7236 9276
rect 7172 9216 7236 9220
rect 12912 9276 12976 9280
rect 12912 9220 12916 9276
rect 12916 9220 12972 9276
rect 12972 9220 12976 9276
rect 12912 9216 12976 9220
rect 12992 9276 13056 9280
rect 12992 9220 12996 9276
rect 12996 9220 13052 9276
rect 13052 9220 13056 9276
rect 12992 9216 13056 9220
rect 13072 9276 13136 9280
rect 13072 9220 13076 9276
rect 13076 9220 13132 9276
rect 13132 9220 13136 9276
rect 13072 9216 13136 9220
rect 13152 9276 13216 9280
rect 13152 9220 13156 9276
rect 13156 9220 13212 9276
rect 13212 9220 13216 9276
rect 13152 9216 13216 9220
rect 3942 8732 4006 8736
rect 3942 8676 3946 8732
rect 3946 8676 4002 8732
rect 4002 8676 4006 8732
rect 3942 8672 4006 8676
rect 4022 8732 4086 8736
rect 4022 8676 4026 8732
rect 4026 8676 4082 8732
rect 4082 8676 4086 8732
rect 4022 8672 4086 8676
rect 4102 8732 4166 8736
rect 4102 8676 4106 8732
rect 4106 8676 4162 8732
rect 4162 8676 4166 8732
rect 4102 8672 4166 8676
rect 4182 8732 4246 8736
rect 4182 8676 4186 8732
rect 4186 8676 4242 8732
rect 4242 8676 4246 8732
rect 4182 8672 4246 8676
rect 9922 8732 9986 8736
rect 9922 8676 9926 8732
rect 9926 8676 9982 8732
rect 9982 8676 9986 8732
rect 9922 8672 9986 8676
rect 10002 8732 10066 8736
rect 10002 8676 10006 8732
rect 10006 8676 10062 8732
rect 10062 8676 10066 8732
rect 10002 8672 10066 8676
rect 10082 8732 10146 8736
rect 10082 8676 10086 8732
rect 10086 8676 10142 8732
rect 10142 8676 10146 8732
rect 10082 8672 10146 8676
rect 10162 8732 10226 8736
rect 10162 8676 10166 8732
rect 10166 8676 10222 8732
rect 10222 8676 10226 8732
rect 10162 8672 10226 8676
rect 15902 8732 15966 8736
rect 15902 8676 15906 8732
rect 15906 8676 15962 8732
rect 15962 8676 15966 8732
rect 15902 8672 15966 8676
rect 15982 8732 16046 8736
rect 15982 8676 15986 8732
rect 15986 8676 16042 8732
rect 16042 8676 16046 8732
rect 15982 8672 16046 8676
rect 16062 8732 16126 8736
rect 16062 8676 16066 8732
rect 16066 8676 16122 8732
rect 16122 8676 16126 8732
rect 16062 8672 16126 8676
rect 16142 8732 16206 8736
rect 16142 8676 16146 8732
rect 16146 8676 16202 8732
rect 16202 8676 16206 8732
rect 16142 8672 16206 8676
rect 6932 8188 6996 8192
rect 6932 8132 6936 8188
rect 6936 8132 6992 8188
rect 6992 8132 6996 8188
rect 6932 8128 6996 8132
rect 7012 8188 7076 8192
rect 7012 8132 7016 8188
rect 7016 8132 7072 8188
rect 7072 8132 7076 8188
rect 7012 8128 7076 8132
rect 7092 8188 7156 8192
rect 7092 8132 7096 8188
rect 7096 8132 7152 8188
rect 7152 8132 7156 8188
rect 7092 8128 7156 8132
rect 7172 8188 7236 8192
rect 7172 8132 7176 8188
rect 7176 8132 7232 8188
rect 7232 8132 7236 8188
rect 7172 8128 7236 8132
rect 12912 8188 12976 8192
rect 12912 8132 12916 8188
rect 12916 8132 12972 8188
rect 12972 8132 12976 8188
rect 12912 8128 12976 8132
rect 12992 8188 13056 8192
rect 12992 8132 12996 8188
rect 12996 8132 13052 8188
rect 13052 8132 13056 8188
rect 12992 8128 13056 8132
rect 13072 8188 13136 8192
rect 13072 8132 13076 8188
rect 13076 8132 13132 8188
rect 13132 8132 13136 8188
rect 13072 8128 13136 8132
rect 13152 8188 13216 8192
rect 13152 8132 13156 8188
rect 13156 8132 13212 8188
rect 13212 8132 13216 8188
rect 13152 8128 13216 8132
rect 3942 7644 4006 7648
rect 3942 7588 3946 7644
rect 3946 7588 4002 7644
rect 4002 7588 4006 7644
rect 3942 7584 4006 7588
rect 4022 7644 4086 7648
rect 4022 7588 4026 7644
rect 4026 7588 4082 7644
rect 4082 7588 4086 7644
rect 4022 7584 4086 7588
rect 4102 7644 4166 7648
rect 4102 7588 4106 7644
rect 4106 7588 4162 7644
rect 4162 7588 4166 7644
rect 4102 7584 4166 7588
rect 4182 7644 4246 7648
rect 4182 7588 4186 7644
rect 4186 7588 4242 7644
rect 4242 7588 4246 7644
rect 4182 7584 4246 7588
rect 9922 7644 9986 7648
rect 9922 7588 9926 7644
rect 9926 7588 9982 7644
rect 9982 7588 9986 7644
rect 9922 7584 9986 7588
rect 10002 7644 10066 7648
rect 10002 7588 10006 7644
rect 10006 7588 10062 7644
rect 10062 7588 10066 7644
rect 10002 7584 10066 7588
rect 10082 7644 10146 7648
rect 10082 7588 10086 7644
rect 10086 7588 10142 7644
rect 10142 7588 10146 7644
rect 10082 7584 10146 7588
rect 10162 7644 10226 7648
rect 10162 7588 10166 7644
rect 10166 7588 10222 7644
rect 10222 7588 10226 7644
rect 10162 7584 10226 7588
rect 15902 7644 15966 7648
rect 15902 7588 15906 7644
rect 15906 7588 15962 7644
rect 15962 7588 15966 7644
rect 15902 7584 15966 7588
rect 15982 7644 16046 7648
rect 15982 7588 15986 7644
rect 15986 7588 16042 7644
rect 16042 7588 16046 7644
rect 15982 7584 16046 7588
rect 16062 7644 16126 7648
rect 16062 7588 16066 7644
rect 16066 7588 16122 7644
rect 16122 7588 16126 7644
rect 16062 7584 16126 7588
rect 16142 7644 16206 7648
rect 16142 7588 16146 7644
rect 16146 7588 16202 7644
rect 16202 7588 16206 7644
rect 16142 7584 16206 7588
rect 6932 7100 6996 7104
rect 6932 7044 6936 7100
rect 6936 7044 6992 7100
rect 6992 7044 6996 7100
rect 6932 7040 6996 7044
rect 7012 7100 7076 7104
rect 7012 7044 7016 7100
rect 7016 7044 7072 7100
rect 7072 7044 7076 7100
rect 7012 7040 7076 7044
rect 7092 7100 7156 7104
rect 7092 7044 7096 7100
rect 7096 7044 7152 7100
rect 7152 7044 7156 7100
rect 7092 7040 7156 7044
rect 7172 7100 7236 7104
rect 7172 7044 7176 7100
rect 7176 7044 7232 7100
rect 7232 7044 7236 7100
rect 7172 7040 7236 7044
rect 12912 7100 12976 7104
rect 12912 7044 12916 7100
rect 12916 7044 12972 7100
rect 12972 7044 12976 7100
rect 12912 7040 12976 7044
rect 12992 7100 13056 7104
rect 12992 7044 12996 7100
rect 12996 7044 13052 7100
rect 13052 7044 13056 7100
rect 12992 7040 13056 7044
rect 13072 7100 13136 7104
rect 13072 7044 13076 7100
rect 13076 7044 13132 7100
rect 13132 7044 13136 7100
rect 13072 7040 13136 7044
rect 13152 7100 13216 7104
rect 13152 7044 13156 7100
rect 13156 7044 13212 7100
rect 13212 7044 13216 7100
rect 13152 7040 13216 7044
rect 3942 6556 4006 6560
rect 3942 6500 3946 6556
rect 3946 6500 4002 6556
rect 4002 6500 4006 6556
rect 3942 6496 4006 6500
rect 4022 6556 4086 6560
rect 4022 6500 4026 6556
rect 4026 6500 4082 6556
rect 4082 6500 4086 6556
rect 4022 6496 4086 6500
rect 4102 6556 4166 6560
rect 4102 6500 4106 6556
rect 4106 6500 4162 6556
rect 4162 6500 4166 6556
rect 4102 6496 4166 6500
rect 4182 6556 4246 6560
rect 4182 6500 4186 6556
rect 4186 6500 4242 6556
rect 4242 6500 4246 6556
rect 4182 6496 4246 6500
rect 9922 6556 9986 6560
rect 9922 6500 9926 6556
rect 9926 6500 9982 6556
rect 9982 6500 9986 6556
rect 9922 6496 9986 6500
rect 10002 6556 10066 6560
rect 10002 6500 10006 6556
rect 10006 6500 10062 6556
rect 10062 6500 10066 6556
rect 10002 6496 10066 6500
rect 10082 6556 10146 6560
rect 10082 6500 10086 6556
rect 10086 6500 10142 6556
rect 10142 6500 10146 6556
rect 10082 6496 10146 6500
rect 10162 6556 10226 6560
rect 10162 6500 10166 6556
rect 10166 6500 10222 6556
rect 10222 6500 10226 6556
rect 10162 6496 10226 6500
rect 15902 6556 15966 6560
rect 15902 6500 15906 6556
rect 15906 6500 15962 6556
rect 15962 6500 15966 6556
rect 15902 6496 15966 6500
rect 15982 6556 16046 6560
rect 15982 6500 15986 6556
rect 15986 6500 16042 6556
rect 16042 6500 16046 6556
rect 15982 6496 16046 6500
rect 16062 6556 16126 6560
rect 16062 6500 16066 6556
rect 16066 6500 16122 6556
rect 16122 6500 16126 6556
rect 16062 6496 16126 6500
rect 16142 6556 16206 6560
rect 16142 6500 16146 6556
rect 16146 6500 16202 6556
rect 16202 6500 16206 6556
rect 16142 6496 16206 6500
rect 6932 6012 6996 6016
rect 6932 5956 6936 6012
rect 6936 5956 6992 6012
rect 6992 5956 6996 6012
rect 6932 5952 6996 5956
rect 7012 6012 7076 6016
rect 7012 5956 7016 6012
rect 7016 5956 7072 6012
rect 7072 5956 7076 6012
rect 7012 5952 7076 5956
rect 7092 6012 7156 6016
rect 7092 5956 7096 6012
rect 7096 5956 7152 6012
rect 7152 5956 7156 6012
rect 7092 5952 7156 5956
rect 7172 6012 7236 6016
rect 7172 5956 7176 6012
rect 7176 5956 7232 6012
rect 7232 5956 7236 6012
rect 7172 5952 7236 5956
rect 12912 6012 12976 6016
rect 12912 5956 12916 6012
rect 12916 5956 12972 6012
rect 12972 5956 12976 6012
rect 12912 5952 12976 5956
rect 12992 6012 13056 6016
rect 12992 5956 12996 6012
rect 12996 5956 13052 6012
rect 13052 5956 13056 6012
rect 12992 5952 13056 5956
rect 13072 6012 13136 6016
rect 13072 5956 13076 6012
rect 13076 5956 13132 6012
rect 13132 5956 13136 6012
rect 13072 5952 13136 5956
rect 13152 6012 13216 6016
rect 13152 5956 13156 6012
rect 13156 5956 13212 6012
rect 13212 5956 13216 6012
rect 13152 5952 13216 5956
rect 3942 5468 4006 5472
rect 3942 5412 3946 5468
rect 3946 5412 4002 5468
rect 4002 5412 4006 5468
rect 3942 5408 4006 5412
rect 4022 5468 4086 5472
rect 4022 5412 4026 5468
rect 4026 5412 4082 5468
rect 4082 5412 4086 5468
rect 4022 5408 4086 5412
rect 4102 5468 4166 5472
rect 4102 5412 4106 5468
rect 4106 5412 4162 5468
rect 4162 5412 4166 5468
rect 4102 5408 4166 5412
rect 4182 5468 4246 5472
rect 4182 5412 4186 5468
rect 4186 5412 4242 5468
rect 4242 5412 4246 5468
rect 4182 5408 4246 5412
rect 9922 5468 9986 5472
rect 9922 5412 9926 5468
rect 9926 5412 9982 5468
rect 9982 5412 9986 5468
rect 9922 5408 9986 5412
rect 10002 5468 10066 5472
rect 10002 5412 10006 5468
rect 10006 5412 10062 5468
rect 10062 5412 10066 5468
rect 10002 5408 10066 5412
rect 10082 5468 10146 5472
rect 10082 5412 10086 5468
rect 10086 5412 10142 5468
rect 10142 5412 10146 5468
rect 10082 5408 10146 5412
rect 10162 5468 10226 5472
rect 10162 5412 10166 5468
rect 10166 5412 10222 5468
rect 10222 5412 10226 5468
rect 10162 5408 10226 5412
rect 15902 5468 15966 5472
rect 15902 5412 15906 5468
rect 15906 5412 15962 5468
rect 15962 5412 15966 5468
rect 15902 5408 15966 5412
rect 15982 5468 16046 5472
rect 15982 5412 15986 5468
rect 15986 5412 16042 5468
rect 16042 5412 16046 5468
rect 15982 5408 16046 5412
rect 16062 5468 16126 5472
rect 16062 5412 16066 5468
rect 16066 5412 16122 5468
rect 16122 5412 16126 5468
rect 16062 5408 16126 5412
rect 16142 5468 16206 5472
rect 16142 5412 16146 5468
rect 16146 5412 16202 5468
rect 16202 5412 16206 5468
rect 16142 5408 16206 5412
rect 6932 4924 6996 4928
rect 6932 4868 6936 4924
rect 6936 4868 6992 4924
rect 6992 4868 6996 4924
rect 6932 4864 6996 4868
rect 7012 4924 7076 4928
rect 7012 4868 7016 4924
rect 7016 4868 7072 4924
rect 7072 4868 7076 4924
rect 7012 4864 7076 4868
rect 7092 4924 7156 4928
rect 7092 4868 7096 4924
rect 7096 4868 7152 4924
rect 7152 4868 7156 4924
rect 7092 4864 7156 4868
rect 7172 4924 7236 4928
rect 7172 4868 7176 4924
rect 7176 4868 7232 4924
rect 7232 4868 7236 4924
rect 7172 4864 7236 4868
rect 12912 4924 12976 4928
rect 12912 4868 12916 4924
rect 12916 4868 12972 4924
rect 12972 4868 12976 4924
rect 12912 4864 12976 4868
rect 12992 4924 13056 4928
rect 12992 4868 12996 4924
rect 12996 4868 13052 4924
rect 13052 4868 13056 4924
rect 12992 4864 13056 4868
rect 13072 4924 13136 4928
rect 13072 4868 13076 4924
rect 13076 4868 13132 4924
rect 13132 4868 13136 4924
rect 13072 4864 13136 4868
rect 13152 4924 13216 4928
rect 13152 4868 13156 4924
rect 13156 4868 13212 4924
rect 13212 4868 13216 4924
rect 13152 4864 13216 4868
rect 3942 4380 4006 4384
rect 3942 4324 3946 4380
rect 3946 4324 4002 4380
rect 4002 4324 4006 4380
rect 3942 4320 4006 4324
rect 4022 4380 4086 4384
rect 4022 4324 4026 4380
rect 4026 4324 4082 4380
rect 4082 4324 4086 4380
rect 4022 4320 4086 4324
rect 4102 4380 4166 4384
rect 4102 4324 4106 4380
rect 4106 4324 4162 4380
rect 4162 4324 4166 4380
rect 4102 4320 4166 4324
rect 4182 4380 4246 4384
rect 4182 4324 4186 4380
rect 4186 4324 4242 4380
rect 4242 4324 4246 4380
rect 4182 4320 4246 4324
rect 9922 4380 9986 4384
rect 9922 4324 9926 4380
rect 9926 4324 9982 4380
rect 9982 4324 9986 4380
rect 9922 4320 9986 4324
rect 10002 4380 10066 4384
rect 10002 4324 10006 4380
rect 10006 4324 10062 4380
rect 10062 4324 10066 4380
rect 10002 4320 10066 4324
rect 10082 4380 10146 4384
rect 10082 4324 10086 4380
rect 10086 4324 10142 4380
rect 10142 4324 10146 4380
rect 10082 4320 10146 4324
rect 10162 4380 10226 4384
rect 10162 4324 10166 4380
rect 10166 4324 10222 4380
rect 10222 4324 10226 4380
rect 10162 4320 10226 4324
rect 15902 4380 15966 4384
rect 15902 4324 15906 4380
rect 15906 4324 15962 4380
rect 15962 4324 15966 4380
rect 15902 4320 15966 4324
rect 15982 4380 16046 4384
rect 15982 4324 15986 4380
rect 15986 4324 16042 4380
rect 16042 4324 16046 4380
rect 15982 4320 16046 4324
rect 16062 4380 16126 4384
rect 16062 4324 16066 4380
rect 16066 4324 16122 4380
rect 16122 4324 16126 4380
rect 16062 4320 16126 4324
rect 16142 4380 16206 4384
rect 16142 4324 16146 4380
rect 16146 4324 16202 4380
rect 16202 4324 16206 4380
rect 16142 4320 16206 4324
rect 6932 3836 6996 3840
rect 6932 3780 6936 3836
rect 6936 3780 6992 3836
rect 6992 3780 6996 3836
rect 6932 3776 6996 3780
rect 7012 3836 7076 3840
rect 7012 3780 7016 3836
rect 7016 3780 7072 3836
rect 7072 3780 7076 3836
rect 7012 3776 7076 3780
rect 7092 3836 7156 3840
rect 7092 3780 7096 3836
rect 7096 3780 7152 3836
rect 7152 3780 7156 3836
rect 7092 3776 7156 3780
rect 7172 3836 7236 3840
rect 7172 3780 7176 3836
rect 7176 3780 7232 3836
rect 7232 3780 7236 3836
rect 7172 3776 7236 3780
rect 12912 3836 12976 3840
rect 12912 3780 12916 3836
rect 12916 3780 12972 3836
rect 12972 3780 12976 3836
rect 12912 3776 12976 3780
rect 12992 3836 13056 3840
rect 12992 3780 12996 3836
rect 12996 3780 13052 3836
rect 13052 3780 13056 3836
rect 12992 3776 13056 3780
rect 13072 3836 13136 3840
rect 13072 3780 13076 3836
rect 13076 3780 13132 3836
rect 13132 3780 13136 3836
rect 13072 3776 13136 3780
rect 13152 3836 13216 3840
rect 13152 3780 13156 3836
rect 13156 3780 13212 3836
rect 13212 3780 13216 3836
rect 13152 3776 13216 3780
rect 3942 3292 4006 3296
rect 3942 3236 3946 3292
rect 3946 3236 4002 3292
rect 4002 3236 4006 3292
rect 3942 3232 4006 3236
rect 4022 3292 4086 3296
rect 4022 3236 4026 3292
rect 4026 3236 4082 3292
rect 4082 3236 4086 3292
rect 4022 3232 4086 3236
rect 4102 3292 4166 3296
rect 4102 3236 4106 3292
rect 4106 3236 4162 3292
rect 4162 3236 4166 3292
rect 4102 3232 4166 3236
rect 4182 3292 4246 3296
rect 4182 3236 4186 3292
rect 4186 3236 4242 3292
rect 4242 3236 4246 3292
rect 4182 3232 4246 3236
rect 9922 3292 9986 3296
rect 9922 3236 9926 3292
rect 9926 3236 9982 3292
rect 9982 3236 9986 3292
rect 9922 3232 9986 3236
rect 10002 3292 10066 3296
rect 10002 3236 10006 3292
rect 10006 3236 10062 3292
rect 10062 3236 10066 3292
rect 10002 3232 10066 3236
rect 10082 3292 10146 3296
rect 10082 3236 10086 3292
rect 10086 3236 10142 3292
rect 10142 3236 10146 3292
rect 10082 3232 10146 3236
rect 10162 3292 10226 3296
rect 10162 3236 10166 3292
rect 10166 3236 10222 3292
rect 10222 3236 10226 3292
rect 10162 3232 10226 3236
rect 15902 3292 15966 3296
rect 15902 3236 15906 3292
rect 15906 3236 15962 3292
rect 15962 3236 15966 3292
rect 15902 3232 15966 3236
rect 15982 3292 16046 3296
rect 15982 3236 15986 3292
rect 15986 3236 16042 3292
rect 16042 3236 16046 3292
rect 15982 3232 16046 3236
rect 16062 3292 16126 3296
rect 16062 3236 16066 3292
rect 16066 3236 16122 3292
rect 16122 3236 16126 3292
rect 16062 3232 16126 3236
rect 16142 3292 16206 3296
rect 16142 3236 16146 3292
rect 16146 3236 16202 3292
rect 16202 3236 16206 3292
rect 16142 3232 16206 3236
rect 6932 2748 6996 2752
rect 6932 2692 6936 2748
rect 6936 2692 6992 2748
rect 6992 2692 6996 2748
rect 6932 2688 6996 2692
rect 7012 2748 7076 2752
rect 7012 2692 7016 2748
rect 7016 2692 7072 2748
rect 7072 2692 7076 2748
rect 7012 2688 7076 2692
rect 7092 2748 7156 2752
rect 7092 2692 7096 2748
rect 7096 2692 7152 2748
rect 7152 2692 7156 2748
rect 7092 2688 7156 2692
rect 7172 2748 7236 2752
rect 7172 2692 7176 2748
rect 7176 2692 7232 2748
rect 7232 2692 7236 2748
rect 7172 2688 7236 2692
rect 12912 2748 12976 2752
rect 12912 2692 12916 2748
rect 12916 2692 12972 2748
rect 12972 2692 12976 2748
rect 12912 2688 12976 2692
rect 12992 2748 13056 2752
rect 12992 2692 12996 2748
rect 12996 2692 13052 2748
rect 13052 2692 13056 2748
rect 12992 2688 13056 2692
rect 13072 2748 13136 2752
rect 13072 2692 13076 2748
rect 13076 2692 13132 2748
rect 13132 2692 13136 2748
rect 13072 2688 13136 2692
rect 13152 2748 13216 2752
rect 13152 2692 13156 2748
rect 13156 2692 13212 2748
rect 13212 2692 13216 2748
rect 13152 2688 13216 2692
rect 3942 2204 4006 2208
rect 3942 2148 3946 2204
rect 3946 2148 4002 2204
rect 4002 2148 4006 2204
rect 3942 2144 4006 2148
rect 4022 2204 4086 2208
rect 4022 2148 4026 2204
rect 4026 2148 4082 2204
rect 4082 2148 4086 2204
rect 4022 2144 4086 2148
rect 4102 2204 4166 2208
rect 4102 2148 4106 2204
rect 4106 2148 4162 2204
rect 4162 2148 4166 2204
rect 4102 2144 4166 2148
rect 4182 2204 4246 2208
rect 4182 2148 4186 2204
rect 4186 2148 4242 2204
rect 4242 2148 4246 2204
rect 4182 2144 4246 2148
rect 9922 2204 9986 2208
rect 9922 2148 9926 2204
rect 9926 2148 9982 2204
rect 9982 2148 9986 2204
rect 9922 2144 9986 2148
rect 10002 2204 10066 2208
rect 10002 2148 10006 2204
rect 10006 2148 10062 2204
rect 10062 2148 10066 2204
rect 10002 2144 10066 2148
rect 10082 2204 10146 2208
rect 10082 2148 10086 2204
rect 10086 2148 10142 2204
rect 10142 2148 10146 2204
rect 10082 2144 10146 2148
rect 10162 2204 10226 2208
rect 10162 2148 10166 2204
rect 10166 2148 10222 2204
rect 10222 2148 10226 2204
rect 10162 2144 10226 2148
rect 15902 2204 15966 2208
rect 15902 2148 15906 2204
rect 15906 2148 15962 2204
rect 15962 2148 15966 2204
rect 15902 2144 15966 2148
rect 15982 2204 16046 2208
rect 15982 2148 15986 2204
rect 15986 2148 16042 2204
rect 16042 2148 16046 2204
rect 15982 2144 16046 2148
rect 16062 2204 16126 2208
rect 16062 2148 16066 2204
rect 16066 2148 16122 2204
rect 16122 2148 16126 2204
rect 16062 2144 16126 2148
rect 16142 2204 16206 2208
rect 16142 2148 16146 2204
rect 16146 2148 16202 2204
rect 16202 2148 16206 2204
rect 16142 2144 16206 2148
<< metal4 >>
rect -916 22106 -596 22148
rect -916 21870 -874 22106
rect -638 21870 -596 22106
rect -916 14214 -596 21870
rect -916 13978 -874 14214
rect -638 13978 -596 14214
rect -916 8230 -596 13978
rect -916 7994 -874 8230
rect -638 7994 -596 8230
rect -916 434 -596 7994
rect -256 21446 64 21488
rect -256 21210 -214 21446
rect 22 21210 64 21446
rect -256 17206 64 21210
rect -256 16970 -214 17206
rect 22 16970 64 17206
rect -256 11222 64 16970
rect -256 10986 -214 11222
rect 22 10986 64 11222
rect -256 5238 64 10986
rect -256 5002 -214 5238
rect 22 5002 64 5238
rect -256 1094 64 5002
rect -256 858 -214 1094
rect 22 858 64 1094
rect -256 816 64 858
rect 3934 21446 4254 22148
rect 3934 21210 3976 21446
rect 4212 21210 4254 21446
rect 3934 19616 4254 21210
rect 3934 19552 3942 19616
rect 4006 19552 4022 19616
rect 4086 19552 4102 19616
rect 4166 19552 4182 19616
rect 4246 19552 4254 19616
rect 3934 18528 4254 19552
rect 3934 18464 3942 18528
rect 4006 18464 4022 18528
rect 4086 18464 4102 18528
rect 4166 18464 4182 18528
rect 4246 18464 4254 18528
rect 3934 17440 4254 18464
rect 3934 17376 3942 17440
rect 4006 17376 4022 17440
rect 4086 17376 4102 17440
rect 4166 17376 4182 17440
rect 4246 17376 4254 17440
rect 3934 17206 4254 17376
rect 3934 16970 3976 17206
rect 4212 16970 4254 17206
rect 3934 16352 4254 16970
rect 3934 16288 3942 16352
rect 4006 16288 4022 16352
rect 4086 16288 4102 16352
rect 4166 16288 4182 16352
rect 4246 16288 4254 16352
rect 3934 15264 4254 16288
rect 3934 15200 3942 15264
rect 4006 15200 4022 15264
rect 4086 15200 4102 15264
rect 4166 15200 4182 15264
rect 4246 15200 4254 15264
rect 3934 14176 4254 15200
rect 3934 14112 3942 14176
rect 4006 14112 4022 14176
rect 4086 14112 4102 14176
rect 4166 14112 4182 14176
rect 4246 14112 4254 14176
rect 3934 13088 4254 14112
rect 3934 13024 3942 13088
rect 4006 13024 4022 13088
rect 4086 13024 4102 13088
rect 4166 13024 4182 13088
rect 4246 13024 4254 13088
rect 3934 12000 4254 13024
rect 3934 11936 3942 12000
rect 4006 11936 4022 12000
rect 4086 11936 4102 12000
rect 4166 11936 4182 12000
rect 4246 11936 4254 12000
rect 3934 11222 4254 11936
rect 3934 10986 3976 11222
rect 4212 10986 4254 11222
rect 3934 10912 4254 10986
rect 3934 10848 3942 10912
rect 4006 10848 4022 10912
rect 4086 10848 4102 10912
rect 4166 10848 4182 10912
rect 4246 10848 4254 10912
rect 3934 9824 4254 10848
rect 3934 9760 3942 9824
rect 4006 9760 4022 9824
rect 4086 9760 4102 9824
rect 4166 9760 4182 9824
rect 4246 9760 4254 9824
rect 3934 8736 4254 9760
rect 3934 8672 3942 8736
rect 4006 8672 4022 8736
rect 4086 8672 4102 8736
rect 4166 8672 4182 8736
rect 4246 8672 4254 8736
rect 3934 7648 4254 8672
rect 3934 7584 3942 7648
rect 4006 7584 4022 7648
rect 4086 7584 4102 7648
rect 4166 7584 4182 7648
rect 4246 7584 4254 7648
rect 3934 6560 4254 7584
rect 3934 6496 3942 6560
rect 4006 6496 4022 6560
rect 4086 6496 4102 6560
rect 4166 6496 4182 6560
rect 4246 6496 4254 6560
rect 3934 5472 4254 6496
rect 3934 5408 3942 5472
rect 4006 5408 4022 5472
rect 4086 5408 4102 5472
rect 4166 5408 4182 5472
rect 4246 5408 4254 5472
rect 3934 5238 4254 5408
rect 3934 5002 3976 5238
rect 4212 5002 4254 5238
rect 3934 4384 4254 5002
rect 3934 4320 3942 4384
rect 4006 4320 4022 4384
rect 4086 4320 4102 4384
rect 4166 4320 4182 4384
rect 4246 4320 4254 4384
rect 3934 3296 4254 4320
rect 3934 3232 3942 3296
rect 4006 3232 4022 3296
rect 4086 3232 4102 3296
rect 4166 3232 4182 3296
rect 4246 3232 4254 3296
rect 3934 2208 4254 3232
rect 3934 2144 3942 2208
rect 4006 2144 4022 2208
rect 4086 2144 4102 2208
rect 4166 2144 4182 2208
rect 4246 2144 4254 2208
rect 3934 1094 4254 2144
rect 3934 858 3976 1094
rect 4212 858 4254 1094
rect -916 198 -874 434
rect -638 198 -596 434
rect -916 156 -596 198
rect 3934 156 4254 858
rect 6924 22106 7244 22148
rect 6924 21870 6966 22106
rect 7202 21870 7244 22106
rect 6924 20160 7244 21870
rect 6924 20096 6932 20160
rect 6996 20096 7012 20160
rect 7076 20096 7092 20160
rect 7156 20096 7172 20160
rect 7236 20096 7244 20160
rect 6924 19072 7244 20096
rect 6924 19008 6932 19072
rect 6996 19008 7012 19072
rect 7076 19008 7092 19072
rect 7156 19008 7172 19072
rect 7236 19008 7244 19072
rect 6924 17984 7244 19008
rect 6924 17920 6932 17984
rect 6996 17920 7012 17984
rect 7076 17920 7092 17984
rect 7156 17920 7172 17984
rect 7236 17920 7244 17984
rect 6924 16896 7244 17920
rect 6924 16832 6932 16896
rect 6996 16832 7012 16896
rect 7076 16832 7092 16896
rect 7156 16832 7172 16896
rect 7236 16832 7244 16896
rect 6924 15808 7244 16832
rect 6924 15744 6932 15808
rect 6996 15744 7012 15808
rect 7076 15744 7092 15808
rect 7156 15744 7172 15808
rect 7236 15744 7244 15808
rect 6924 14720 7244 15744
rect 6924 14656 6932 14720
rect 6996 14656 7012 14720
rect 7076 14656 7092 14720
rect 7156 14656 7172 14720
rect 7236 14656 7244 14720
rect 6924 14214 7244 14656
rect 6924 13978 6966 14214
rect 7202 13978 7244 14214
rect 6924 13632 7244 13978
rect 6924 13568 6932 13632
rect 6996 13568 7012 13632
rect 7076 13568 7092 13632
rect 7156 13568 7172 13632
rect 7236 13568 7244 13632
rect 6924 12544 7244 13568
rect 6924 12480 6932 12544
rect 6996 12480 7012 12544
rect 7076 12480 7092 12544
rect 7156 12480 7172 12544
rect 7236 12480 7244 12544
rect 6924 11456 7244 12480
rect 6924 11392 6932 11456
rect 6996 11392 7012 11456
rect 7076 11392 7092 11456
rect 7156 11392 7172 11456
rect 7236 11392 7244 11456
rect 6924 10368 7244 11392
rect 6924 10304 6932 10368
rect 6996 10304 7012 10368
rect 7076 10304 7092 10368
rect 7156 10304 7172 10368
rect 7236 10304 7244 10368
rect 6924 9280 7244 10304
rect 6924 9216 6932 9280
rect 6996 9216 7012 9280
rect 7076 9216 7092 9280
rect 7156 9216 7172 9280
rect 7236 9216 7244 9280
rect 6924 8230 7244 9216
rect 6924 8192 6966 8230
rect 7202 8192 7244 8230
rect 6924 8128 6932 8192
rect 7236 8128 7244 8192
rect 6924 7994 6966 8128
rect 7202 7994 7244 8128
rect 6924 7104 7244 7994
rect 6924 7040 6932 7104
rect 6996 7040 7012 7104
rect 7076 7040 7092 7104
rect 7156 7040 7172 7104
rect 7236 7040 7244 7104
rect 6924 6016 7244 7040
rect 6924 5952 6932 6016
rect 6996 5952 7012 6016
rect 7076 5952 7092 6016
rect 7156 5952 7172 6016
rect 7236 5952 7244 6016
rect 6924 4928 7244 5952
rect 6924 4864 6932 4928
rect 6996 4864 7012 4928
rect 7076 4864 7092 4928
rect 7156 4864 7172 4928
rect 7236 4864 7244 4928
rect 6924 3840 7244 4864
rect 6924 3776 6932 3840
rect 6996 3776 7012 3840
rect 7076 3776 7092 3840
rect 7156 3776 7172 3840
rect 7236 3776 7244 3840
rect 6924 2752 7244 3776
rect 6924 2688 6932 2752
rect 6996 2688 7012 2752
rect 7076 2688 7092 2752
rect 7156 2688 7172 2752
rect 7236 2688 7244 2752
rect 6924 434 7244 2688
rect 6924 198 6966 434
rect 7202 198 7244 434
rect 6924 156 7244 198
rect 9914 21446 10234 22148
rect 9914 21210 9956 21446
rect 10192 21210 10234 21446
rect 9914 19616 10234 21210
rect 9914 19552 9922 19616
rect 9986 19552 10002 19616
rect 10066 19552 10082 19616
rect 10146 19552 10162 19616
rect 10226 19552 10234 19616
rect 9914 18528 10234 19552
rect 9914 18464 9922 18528
rect 9986 18464 10002 18528
rect 10066 18464 10082 18528
rect 10146 18464 10162 18528
rect 10226 18464 10234 18528
rect 9914 17440 10234 18464
rect 9914 17376 9922 17440
rect 9986 17376 10002 17440
rect 10066 17376 10082 17440
rect 10146 17376 10162 17440
rect 10226 17376 10234 17440
rect 9914 17206 10234 17376
rect 9914 16970 9956 17206
rect 10192 16970 10234 17206
rect 9914 16352 10234 16970
rect 9914 16288 9922 16352
rect 9986 16288 10002 16352
rect 10066 16288 10082 16352
rect 10146 16288 10162 16352
rect 10226 16288 10234 16352
rect 9914 15264 10234 16288
rect 9914 15200 9922 15264
rect 9986 15200 10002 15264
rect 10066 15200 10082 15264
rect 10146 15200 10162 15264
rect 10226 15200 10234 15264
rect 9914 14176 10234 15200
rect 9914 14112 9922 14176
rect 9986 14112 10002 14176
rect 10066 14112 10082 14176
rect 10146 14112 10162 14176
rect 10226 14112 10234 14176
rect 9914 13088 10234 14112
rect 9914 13024 9922 13088
rect 9986 13024 10002 13088
rect 10066 13024 10082 13088
rect 10146 13024 10162 13088
rect 10226 13024 10234 13088
rect 9914 12000 10234 13024
rect 9914 11936 9922 12000
rect 9986 11936 10002 12000
rect 10066 11936 10082 12000
rect 10146 11936 10162 12000
rect 10226 11936 10234 12000
rect 9914 11222 10234 11936
rect 9914 10986 9956 11222
rect 10192 10986 10234 11222
rect 9914 10912 10234 10986
rect 9914 10848 9922 10912
rect 9986 10848 10002 10912
rect 10066 10848 10082 10912
rect 10146 10848 10162 10912
rect 10226 10848 10234 10912
rect 9914 9824 10234 10848
rect 9914 9760 9922 9824
rect 9986 9760 10002 9824
rect 10066 9760 10082 9824
rect 10146 9760 10162 9824
rect 10226 9760 10234 9824
rect 9914 8736 10234 9760
rect 9914 8672 9922 8736
rect 9986 8672 10002 8736
rect 10066 8672 10082 8736
rect 10146 8672 10162 8736
rect 10226 8672 10234 8736
rect 9914 7648 10234 8672
rect 9914 7584 9922 7648
rect 9986 7584 10002 7648
rect 10066 7584 10082 7648
rect 10146 7584 10162 7648
rect 10226 7584 10234 7648
rect 9914 6560 10234 7584
rect 9914 6496 9922 6560
rect 9986 6496 10002 6560
rect 10066 6496 10082 6560
rect 10146 6496 10162 6560
rect 10226 6496 10234 6560
rect 9914 5472 10234 6496
rect 9914 5408 9922 5472
rect 9986 5408 10002 5472
rect 10066 5408 10082 5472
rect 10146 5408 10162 5472
rect 10226 5408 10234 5472
rect 9914 5238 10234 5408
rect 9914 5002 9956 5238
rect 10192 5002 10234 5238
rect 9914 4384 10234 5002
rect 9914 4320 9922 4384
rect 9986 4320 10002 4384
rect 10066 4320 10082 4384
rect 10146 4320 10162 4384
rect 10226 4320 10234 4384
rect 9914 3296 10234 4320
rect 9914 3232 9922 3296
rect 9986 3232 10002 3296
rect 10066 3232 10082 3296
rect 10146 3232 10162 3296
rect 10226 3232 10234 3296
rect 9914 2208 10234 3232
rect 9914 2144 9922 2208
rect 9986 2144 10002 2208
rect 10066 2144 10082 2208
rect 10146 2144 10162 2208
rect 10226 2144 10234 2208
rect 9914 1094 10234 2144
rect 9914 858 9956 1094
rect 10192 858 10234 1094
rect 9914 156 10234 858
rect 12904 22106 13224 22148
rect 12904 21870 12946 22106
rect 13182 21870 13224 22106
rect 12904 20160 13224 21870
rect 12904 20096 12912 20160
rect 12976 20096 12992 20160
rect 13056 20096 13072 20160
rect 13136 20096 13152 20160
rect 13216 20096 13224 20160
rect 12904 19072 13224 20096
rect 12904 19008 12912 19072
rect 12976 19008 12992 19072
rect 13056 19008 13072 19072
rect 13136 19008 13152 19072
rect 13216 19008 13224 19072
rect 12904 17984 13224 19008
rect 12904 17920 12912 17984
rect 12976 17920 12992 17984
rect 13056 17920 13072 17984
rect 13136 17920 13152 17984
rect 13216 17920 13224 17984
rect 12904 16896 13224 17920
rect 12904 16832 12912 16896
rect 12976 16832 12992 16896
rect 13056 16832 13072 16896
rect 13136 16832 13152 16896
rect 13216 16832 13224 16896
rect 12904 15808 13224 16832
rect 12904 15744 12912 15808
rect 12976 15744 12992 15808
rect 13056 15744 13072 15808
rect 13136 15744 13152 15808
rect 13216 15744 13224 15808
rect 12904 14720 13224 15744
rect 12904 14656 12912 14720
rect 12976 14656 12992 14720
rect 13056 14656 13072 14720
rect 13136 14656 13152 14720
rect 13216 14656 13224 14720
rect 12904 14214 13224 14656
rect 12904 13978 12946 14214
rect 13182 13978 13224 14214
rect 12904 13632 13224 13978
rect 12904 13568 12912 13632
rect 12976 13568 12992 13632
rect 13056 13568 13072 13632
rect 13136 13568 13152 13632
rect 13216 13568 13224 13632
rect 12904 12544 13224 13568
rect 12904 12480 12912 12544
rect 12976 12480 12992 12544
rect 13056 12480 13072 12544
rect 13136 12480 13152 12544
rect 13216 12480 13224 12544
rect 12904 11456 13224 12480
rect 12904 11392 12912 11456
rect 12976 11392 12992 11456
rect 13056 11392 13072 11456
rect 13136 11392 13152 11456
rect 13216 11392 13224 11456
rect 12904 10368 13224 11392
rect 12904 10304 12912 10368
rect 12976 10304 12992 10368
rect 13056 10304 13072 10368
rect 13136 10304 13152 10368
rect 13216 10304 13224 10368
rect 12904 9280 13224 10304
rect 12904 9216 12912 9280
rect 12976 9216 12992 9280
rect 13056 9216 13072 9280
rect 13136 9216 13152 9280
rect 13216 9216 13224 9280
rect 12904 8230 13224 9216
rect 12904 8192 12946 8230
rect 13182 8192 13224 8230
rect 12904 8128 12912 8192
rect 13216 8128 13224 8192
rect 12904 7994 12946 8128
rect 13182 7994 13224 8128
rect 12904 7104 13224 7994
rect 12904 7040 12912 7104
rect 12976 7040 12992 7104
rect 13056 7040 13072 7104
rect 13136 7040 13152 7104
rect 13216 7040 13224 7104
rect 12904 6016 13224 7040
rect 12904 5952 12912 6016
rect 12976 5952 12992 6016
rect 13056 5952 13072 6016
rect 13136 5952 13152 6016
rect 13216 5952 13224 6016
rect 12904 4928 13224 5952
rect 12904 4864 12912 4928
rect 12976 4864 12992 4928
rect 13056 4864 13072 4928
rect 13136 4864 13152 4928
rect 13216 4864 13224 4928
rect 12904 3840 13224 4864
rect 12904 3776 12912 3840
rect 12976 3776 12992 3840
rect 13056 3776 13072 3840
rect 13136 3776 13152 3840
rect 13216 3776 13224 3840
rect 12904 2752 13224 3776
rect 12904 2688 12912 2752
rect 12976 2688 12992 2752
rect 13056 2688 13072 2752
rect 13136 2688 13152 2752
rect 13216 2688 13224 2752
rect 12904 434 13224 2688
rect 12904 198 12946 434
rect 13182 198 13224 434
rect 12904 156 13224 198
rect 15894 21446 16214 22148
rect 20744 22106 21064 22148
rect 20744 21870 20786 22106
rect 21022 21870 21064 22106
rect 15894 21210 15936 21446
rect 16172 21210 16214 21446
rect 15894 19616 16214 21210
rect 15894 19552 15902 19616
rect 15966 19552 15982 19616
rect 16046 19552 16062 19616
rect 16126 19552 16142 19616
rect 16206 19552 16214 19616
rect 15894 18528 16214 19552
rect 15894 18464 15902 18528
rect 15966 18464 15982 18528
rect 16046 18464 16062 18528
rect 16126 18464 16142 18528
rect 16206 18464 16214 18528
rect 15894 17440 16214 18464
rect 15894 17376 15902 17440
rect 15966 17376 15982 17440
rect 16046 17376 16062 17440
rect 16126 17376 16142 17440
rect 16206 17376 16214 17440
rect 15894 17206 16214 17376
rect 15894 16970 15936 17206
rect 16172 16970 16214 17206
rect 15894 16352 16214 16970
rect 15894 16288 15902 16352
rect 15966 16288 15982 16352
rect 16046 16288 16062 16352
rect 16126 16288 16142 16352
rect 16206 16288 16214 16352
rect 15894 15264 16214 16288
rect 15894 15200 15902 15264
rect 15966 15200 15982 15264
rect 16046 15200 16062 15264
rect 16126 15200 16142 15264
rect 16206 15200 16214 15264
rect 15894 14176 16214 15200
rect 15894 14112 15902 14176
rect 15966 14112 15982 14176
rect 16046 14112 16062 14176
rect 16126 14112 16142 14176
rect 16206 14112 16214 14176
rect 15894 13088 16214 14112
rect 15894 13024 15902 13088
rect 15966 13024 15982 13088
rect 16046 13024 16062 13088
rect 16126 13024 16142 13088
rect 16206 13024 16214 13088
rect 15894 12000 16214 13024
rect 15894 11936 15902 12000
rect 15966 11936 15982 12000
rect 16046 11936 16062 12000
rect 16126 11936 16142 12000
rect 16206 11936 16214 12000
rect 15894 11222 16214 11936
rect 15894 10986 15936 11222
rect 16172 10986 16214 11222
rect 15894 10912 16214 10986
rect 15894 10848 15902 10912
rect 15966 10848 15982 10912
rect 16046 10848 16062 10912
rect 16126 10848 16142 10912
rect 16206 10848 16214 10912
rect 15894 9824 16214 10848
rect 15894 9760 15902 9824
rect 15966 9760 15982 9824
rect 16046 9760 16062 9824
rect 16126 9760 16142 9824
rect 16206 9760 16214 9824
rect 15894 8736 16214 9760
rect 15894 8672 15902 8736
rect 15966 8672 15982 8736
rect 16046 8672 16062 8736
rect 16126 8672 16142 8736
rect 16206 8672 16214 8736
rect 15894 7648 16214 8672
rect 15894 7584 15902 7648
rect 15966 7584 15982 7648
rect 16046 7584 16062 7648
rect 16126 7584 16142 7648
rect 16206 7584 16214 7648
rect 15894 6560 16214 7584
rect 15894 6496 15902 6560
rect 15966 6496 15982 6560
rect 16046 6496 16062 6560
rect 16126 6496 16142 6560
rect 16206 6496 16214 6560
rect 15894 5472 16214 6496
rect 15894 5408 15902 5472
rect 15966 5408 15982 5472
rect 16046 5408 16062 5472
rect 16126 5408 16142 5472
rect 16206 5408 16214 5472
rect 15894 5238 16214 5408
rect 15894 5002 15936 5238
rect 16172 5002 16214 5238
rect 15894 4384 16214 5002
rect 15894 4320 15902 4384
rect 15966 4320 15982 4384
rect 16046 4320 16062 4384
rect 16126 4320 16142 4384
rect 16206 4320 16214 4384
rect 15894 3296 16214 4320
rect 15894 3232 15902 3296
rect 15966 3232 15982 3296
rect 16046 3232 16062 3296
rect 16126 3232 16142 3296
rect 16206 3232 16214 3296
rect 15894 2208 16214 3232
rect 15894 2144 15902 2208
rect 15966 2144 15982 2208
rect 16046 2144 16062 2208
rect 16126 2144 16142 2208
rect 16206 2144 16214 2208
rect 15894 1094 16214 2144
rect 15894 858 15936 1094
rect 16172 858 16214 1094
rect 15894 156 16214 858
rect 20084 21446 20404 21488
rect 20084 21210 20126 21446
rect 20362 21210 20404 21446
rect 20084 17206 20404 21210
rect 20084 16970 20126 17206
rect 20362 16970 20404 17206
rect 20084 11222 20404 16970
rect 20084 10986 20126 11222
rect 20362 10986 20404 11222
rect 20084 5238 20404 10986
rect 20084 5002 20126 5238
rect 20362 5002 20404 5238
rect 20084 1094 20404 5002
rect 20084 858 20126 1094
rect 20362 858 20404 1094
rect 20084 816 20404 858
rect 20744 14214 21064 21870
rect 20744 13978 20786 14214
rect 21022 13978 21064 14214
rect 20744 8230 21064 13978
rect 20744 7994 20786 8230
rect 21022 7994 21064 8230
rect 20744 434 21064 7994
rect 20744 198 20786 434
rect 21022 198 21064 434
rect 20744 156 21064 198
<< via4 >>
rect -874 21870 -638 22106
rect -874 13978 -638 14214
rect -874 7994 -638 8230
rect -214 21210 22 21446
rect -214 16970 22 17206
rect -214 10986 22 11222
rect -214 5002 22 5238
rect -214 858 22 1094
rect 3976 21210 4212 21446
rect 3976 16970 4212 17206
rect 3976 10986 4212 11222
rect 3976 5002 4212 5238
rect 3976 858 4212 1094
rect -874 198 -638 434
rect 6966 21870 7202 22106
rect 6966 13978 7202 14214
rect 6966 8192 7202 8230
rect 6966 8128 6996 8192
rect 6996 8128 7012 8192
rect 7012 8128 7076 8192
rect 7076 8128 7092 8192
rect 7092 8128 7156 8192
rect 7156 8128 7172 8192
rect 7172 8128 7202 8192
rect 6966 7994 7202 8128
rect 6966 198 7202 434
rect 9956 21210 10192 21446
rect 9956 16970 10192 17206
rect 9956 10986 10192 11222
rect 9956 5002 10192 5238
rect 9956 858 10192 1094
rect 12946 21870 13182 22106
rect 12946 13978 13182 14214
rect 12946 8192 13182 8230
rect 12946 8128 12976 8192
rect 12976 8128 12992 8192
rect 12992 8128 13056 8192
rect 13056 8128 13072 8192
rect 13072 8128 13136 8192
rect 13136 8128 13152 8192
rect 13152 8128 13182 8192
rect 12946 7994 13182 8128
rect 12946 198 13182 434
rect 20786 21870 21022 22106
rect 15936 21210 16172 21446
rect 15936 16970 16172 17206
rect 15936 10986 16172 11222
rect 15936 5002 16172 5238
rect 15936 858 16172 1094
rect 20126 21210 20362 21446
rect 20126 16970 20362 17206
rect 20126 10986 20362 11222
rect 20126 5002 20362 5238
rect 20126 858 20362 1094
rect 20786 13978 21022 14214
rect 20786 7994 21022 8230
rect 20786 198 21022 434
<< metal5 >>
rect -916 22106 21064 22148
rect -916 21870 -874 22106
rect -638 21870 6966 22106
rect 7202 21870 12946 22106
rect 13182 21870 20786 22106
rect 21022 21870 21064 22106
rect -916 21828 21064 21870
rect -256 21446 20404 21488
rect -256 21210 -214 21446
rect 22 21210 3976 21446
rect 4212 21210 9956 21446
rect 10192 21210 15936 21446
rect 16172 21210 20126 21446
rect 20362 21210 20404 21446
rect -256 21168 20404 21210
rect -916 17206 21064 17248
rect -916 16970 -214 17206
rect 22 16970 3976 17206
rect 4212 16970 9956 17206
rect 10192 16970 15936 17206
rect 16172 16970 20126 17206
rect 20362 16970 21064 17206
rect -916 16928 21064 16970
rect -916 14214 21064 14256
rect -916 13978 -874 14214
rect -638 13978 6966 14214
rect 7202 13978 12946 14214
rect 13182 13978 20786 14214
rect 21022 13978 21064 14214
rect -916 13936 21064 13978
rect -916 11222 21064 11264
rect -916 10986 -214 11222
rect 22 10986 3976 11222
rect 4212 10986 9956 11222
rect 10192 10986 15936 11222
rect 16172 10986 20126 11222
rect 20362 10986 21064 11222
rect -916 10944 21064 10986
rect -916 8230 21064 8272
rect -916 7994 -874 8230
rect -638 7994 6966 8230
rect 7202 7994 12946 8230
rect 13182 7994 20786 8230
rect 21022 7994 21064 8230
rect -916 7952 21064 7994
rect -916 5238 21064 5280
rect -916 5002 -214 5238
rect 22 5002 3976 5238
rect 4212 5002 9956 5238
rect 10192 5002 15936 5238
rect 16172 5002 20126 5238
rect 20362 5002 21064 5238
rect -916 4960 21064 5002
rect -256 1094 20404 1136
rect -256 858 -214 1094
rect 22 858 3976 1094
rect 4212 858 9956 1094
rect 10192 858 15936 1094
rect 16172 858 20126 1094
rect 20362 858 20404 1094
rect -256 816 20404 858
rect -916 434 21064 476
rect -916 198 -874 434
rect -638 198 6966 434
rect 7202 198 12946 434
rect 13182 198 20786 434
rect 21022 198 21064 434
rect -916 156 21064 198
use sky130_fd_sc_hd__decap_8  FILLER_0_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 2208 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 2208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1618419204
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_18
timestamp 1618419204
transform 1 0 2760 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 2944 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 3404 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 1656 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrbp_2  idiv2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 3036 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1618419204
transform -1 0 4876 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25
timestamp 1618419204
transform 1 0 3404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30
timestamp 1618419204
transform 1 0 3864 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41
timestamp 1618419204
transform 1 0 4876 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1618419204
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_45
timestamp 1618419204
transform 1 0 5244 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_58
timestamp 1618419204
transform 1 0 6440 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1618419204
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1618419204
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1618419204
transform -1 0 6072 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1618419204
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1618419204
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_67 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 7268 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67
timestamp 1618419204
transform 1 0 7268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63
timestamp 1618419204
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1618419204
transform -1 0 7268 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  irb $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 6808 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 7820 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _369_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 7636 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _356_
timestamp 1618419204
transform -1 0 10396 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb0
timestamp 1618419204
transform 1 0 9936 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1618419204
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1618419204
transform 1 0 9200 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80
timestamp 1618419204
transform 1 0 8464 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86
timestamp 1618419204
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1618419204
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_80
timestamp 1618419204
transform 1 0 8464 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_92
timestamp 1618419204
transform 1 0 9568 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1618419204
transform 1 0 10580 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_108
timestamp 1618419204
transform 1 0 11040 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101
timestamp 1618419204
transform 1 0 10396 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 11224 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 10764 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_115
timestamp 1618419204
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1618419204
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117
timestamp 1618419204
transform 1 0 11868 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1618419204
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1618419204
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb1
timestamp 1618419204
transform -1 0 12696 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_1_132
timestamp 1618419204
transform 1 0 13248 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_126
timestamp 1618419204
transform 1 0 12696 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_128
timestamp 1618419204
transform 1 0 12880 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 14076 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb0
timestamp 1618419204
transform -1 0 13984 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1618419204
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_140
timestamp 1618419204
transform 1 0 13984 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1618419204
transform 1 0 14536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1618419204
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1618419204
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfrbp_1  idiv16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 16468 0 1 2720
box -38 -48 2154 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1618419204
transform 1 0 14904 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1618419204
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1618419204
transform 1 0 16100 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_159
timestamp 1618419204
transform 1 0 15732 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_167
timestamp 1618419204
transform 1 0 16468 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1618419204
transform 1 0 17020 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_167
timestamp 1618419204
transform 1 0 16468 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1618419204
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_179
timestamp 1618419204
transform 1 0 17572 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_175
timestamp 1618419204
transform 1 0 17204 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1618419204
transform 1 0 17296 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1618419204
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1618419204
transform 1 0 18400 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_191
timestamp 1618419204
transform 1 0 18676 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1618419204
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output43
timestamp 1618419204
transform -1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1618419204
transform -1 0 18400 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1618419204
transform -1 0 19044 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1618419204
transform -1 0 19044 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1618419204
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1618419204
transform -1 0 1656 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_6
timestamp 1618419204
transform 1 0 1656 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1618419204
transform 1 0 2760 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfrbp_2  idiv4
timestamp 1618419204
transform -1 0 6440 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1618419204
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_26
timestamp 1618419204
transform 1 0 3496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_30
timestamp 1618419204
transform 1 0 3864 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 7912 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1618419204
transform -1 0 7544 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_58
timestamp 1618419204
transform 1 0 6440 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_66
timestamp 1618419204
transform 1 0 7176 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_70
timestamp 1618419204
transform 1 0 7544 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1618419204
transform 1 0 9476 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1618419204
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_79
timestamp 1618419204
transform 1 0 8372 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1618419204
transform 1 0 8924 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1618419204
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_94
timestamp 1618419204
transform 1 0 9752 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen0
timestamp 1618419204
transform 1 0 10580 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen1
timestamp 1618419204
transform -1 0 12696 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1618419204
transform -1 0 11776 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_102
timestamp 1618419204
transform 1 0 10488 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1618419204
transform 1 0 11040 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_116
timestamp 1618419204
transform 1 0 11776 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_120
timestamp 1618419204
transform 1 0 12144 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1618419204
transform 1 0 13248 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen0
timestamp 1618419204
transform 1 0 14720 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1618419204
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_126
timestamp 1618419204
transform 1 0 12696 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_135
timestamp 1618419204
transform 1 0 13524 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_144
timestamp 1618419204
transform 1 0 14352 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrbp_2  idiv8
timestamp 1618419204
transform 1 0 15548 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_4  FILLER_2_153
timestamp 1618419204
transform 1 0 15180 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1618419204
transform -1 0 19044 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1618419204
transform 1 0 18124 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_181
timestamp 1618419204
transform 1 0 17756 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_188
timestamp 1618419204
transform 1 0 18400 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1618419204
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1618419204
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1618419204
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1618419204
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1618419204
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _368_
timestamp 1618419204
transform -1 0 7728 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1618419204
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1618419204
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_58
timestamp 1618419204
transform 1 0 6440 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_62
timestamp 1618419204
transform 1 0 6808 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_72
timestamp 1618419204
transform 1 0 7728 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1618419204
transform 1 0 9844 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb0
timestamp 1618419204
transform 1 0 8096 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1618419204
transform -1 0 9476 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_83
timestamp 1618419204
transform 1 0 8740 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_87
timestamp 1618419204
transform 1 0 9108 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_91
timestamp 1618419204
transform 1 0 9476 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp 1618419204
transform -1 0 12880 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1618419204
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1618419204
transform 1 0 10672 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_112
timestamp 1618419204
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1618419204
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1618419204
transform -1 0 14628 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb1
timestamp 1618419204
transform 1 0 13248 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_3_128
timestamp 1618419204
transform 1 0 12880 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_139
timestamp 1618419204
transform 1 0 13892 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_147
timestamp 1618419204
transform 1 0 14628 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1618419204
transform 1 0 14996 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1618419204
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_154
timestamp 1618419204
transform 1 0 15272 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_166
timestamp 1618419204
transform 1 0 16376 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_170
timestamp 1618419204
transform 1 0 16744 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_172
timestamp 1618419204
transform 1 0 16928 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1618419204
transform -1 0 19044 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_184
timestamp 1618419204
transform 1 0 18032 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  ringosc.ibufp11
timestamp 1618419204
transform -1 0 2484 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1618419204
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output41
timestamp 1618419204
transform -1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_7
timestamp 1618419204
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_11
timestamp 1618419204
transform 1 0 2116 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1618419204
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1618419204
transform 1 0 5612 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1618419204
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1618419204
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1618419204
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_42
timestamp 1618419204
transform 1 0 4968 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_48
timestamp 1618419204
transform 1 0 5520 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen0
timestamp 1618419204
transform -1 0 7728 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1618419204
transform -1 0 6624 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_52
timestamp 1618419204
transform 1 0 5888 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_60
timestamp 1618419204
transform 1 0 6624 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_66
timestamp 1618419204
transform 1 0 7176 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_72
timestamp 1618419204
transform 1 0 7728 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[11\].id.delayenb1
timestamp 1618419204
transform 1 0 10028 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1618419204
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1618419204
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_87
timestamp 1618419204
transform 1 0 9108 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_95
timestamp 1618419204
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  repeater46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 12512 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_104
timestamp 1618419204
transform 1 0 10672 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_124
timestamp 1618419204
transform 1 0 12512 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen1
timestamp 1618419204
transform 1 0 12880 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1618419204
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_133
timestamp 1618419204
transform 1 0 13340 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1618419204
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144
timestamp 1618419204
transform 1 0 14352 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1618419204
transform 1 0 16008 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_4_156
timestamp 1618419204
transform 1 0 15456 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_171
timestamp 1618419204
transform 1 0 16836 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1618419204
transform -1 0 19044 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1618419204
transform -1 0 18400 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_183
timestamp 1618419204
transform 1 0 17940 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_188
timestamp 1618419204
transform 1 0 18400 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1618419204
transform 1 0 3220 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  ringosc.ibufp10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 2852 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1618419204
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1618419204
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_15
timestamp 1618419204
transform 1 0 2484 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_19
timestamp 1618419204
transform 1 0 2852 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[5\].id.delayenb1
timestamp 1618419204
transform 1 0 4876 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1618419204
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_39
timestamp 1618419204
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_48
timestamp 1618419204
transform 1 0 5520 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 6808 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1618419204
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_56
timestamp 1618419204
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_58
timestamp 1618419204
transform 1 0 6440 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_67
timestamp 1618419204
transform 1 0 7268 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[11\].id.delayen1
timestamp 1618419204
transform 1 0 10120 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_5_79
timestamp 1618419204
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_91
timestamp 1618419204
transform 1 0 9476 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_97
timestamp 1618419204
transform 1 0 10028 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1618419204
transform 1 0 10948 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1618419204
transform -1 0 12788 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1618419204
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_103
timestamp 1618419204
transform 1 0 10580 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_110
timestamp 1618419204
transform 1 0 11224 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_115
timestamp 1618419204
transform 1 0 11684 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1618419204
transform 1 0 13156 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_127
timestamp 1618419204
transform 1 0 12788 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_134
timestamp 1618419204
transform 1 0 13432 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_146
timestamp 1618419204
transform 1 0 14536 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1618419204
transform -1 0 16468 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1618419204
transform 1 0 14996 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1618419204
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_150
timestamp 1618419204
transform 1 0 14904 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_160
timestamp 1618419204
transform 1 0 15824 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_167
timestamp 1618419204
transform 1 0 16468 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_172
timestamp 1618419204
transform 1 0 16928 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 17296 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1618419204
transform -1 0 19044 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_184
timestamp 1618419204
transform 1 0 18032 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1618419204
transform -1 0 3404 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1618419204
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1618419204
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1618419204
transform -1 0 1656 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1618419204
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_15
timestamp 1618419204
transform 1 0 2484 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_6
timestamp 1618419204
transform 1 0 1656 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_18
timestamp 1618419204
transform 1 0 2760 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_30
timestamp 1618419204
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_30
timestamp 1618419204
transform 1 0 3864 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_25
timestamp 1618419204
transform 1 0 3404 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1618419204
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 4232 0 -1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 4048 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_7_46
timestamp 1618419204
transform 1 0 5336 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_39
timestamp 1618419204
transform 1 0 4692 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_45
timestamp 1618419204
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1618419204
transform -1 0 5336 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[5\].id.delayen1
timestamp 1618419204
transform -1 0 6072 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1618419204
transform 1 0 6624 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.delayen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 6992 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1618419204
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_54
timestamp 1618419204
transform 1 0 6072 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_69
timestamp 1618419204
transform 1 0 7452 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_54
timestamp 1618419204
transform 1 0 6072 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_58
timestamp 1618419204
transform 1 0 6440 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_75
timestamp 1618419204
transform 1 0 8004 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_82
timestamp 1618419204
transform 1 0 8648 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1618419204
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb0
timestamp 1618419204
transform 1 0 8372 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.delayen1
timestamp 1618419204
transform 1 0 8188 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_7_98
timestamp 1618419204
transform 1 0 10120 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_90
timestamp 1618419204
transform 1 0 9384 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_94
timestamp 1618419204
transform 1 0 9752 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1618419204
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1618419204
transform 1 0 9476 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_4  ringosc.dstage\[11\].id.delayen0
timestamp 1618419204
transform 1 0 10212 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1618419204
transform 1 0 10672 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen0
timestamp 1618419204
transform 1 0 12328 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb0
timestamp 1618419204
transform 1 0 12052 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1618419204
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_102
timestamp 1618419204
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_107
timestamp 1618419204
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_110
timestamp 1618419204
transform 1 0 11224 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_115
timestamp 1618419204
transform 1 0 11684 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1618419204
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_2  _322_
timestamp 1618419204
transform -1 0 15364 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1618419204
transform -1 0 15548 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1618419204
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_126
timestamp 1618419204
transform 1 0 12696 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_138
timestamp 1618419204
transform 1 0 13800 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_142
timestamp 1618419204
transform 1 0 14168 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_144
timestamp 1618419204
transform 1 0 14352 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1618419204
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_139
timestamp 1618419204
transform 1 0 13892 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1618419204
transform 1 0 17020 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _323_
timestamp 1618419204
transform 1 0 15732 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _324_
timestamp 1618419204
transform -1 0 16652 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1618419204
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_157
timestamp 1618419204
transform 1 0 15548 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_169
timestamp 1618419204
transform 1 0 16652 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_155
timestamp 1618419204
transform 1 0 15364 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_167
timestamp 1618419204
transform 1 0 16468 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_172
timestamp 1618419204
transform 1 0 16928 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1618419204
transform -1 0 19044 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1618419204
transform -1 0 19044 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_176
timestamp 1618419204
transform 1 0 17296 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_188
timestamp 1618419204
transform 1 0 18400 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_184
timestamp 1618419204
transform 1 0 18032 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _360_
timestamp 1618419204
transform 1 0 1748 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen0
timestamp 1618419204
transform 1 0 2944 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1618419204
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1618419204
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_16
timestamp 1618419204
transform 1 0 2576 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _372_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 5428 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1618419204
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_25
timestamp 1618419204
transform 1 0 3404 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_30
timestamp 1618419204
transform 1 0 3864 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_47
timestamp 1618419204
transform 1 0 5428 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 6256 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.reseten0
timestamp 1618419204
transform -1 0 7636 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_8_56
timestamp 1618419204
transform 1 0 6256 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_71
timestamp 1618419204
transform 1 0 7636 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb0
timestamp 1618419204
transform 1 0 9936 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_2  ringosc.iss.delayenb1
timestamp 1618419204
transform 1 0 8004 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1618419204
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_82
timestamp 1618419204
transform 1 0 8648 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_87
timestamp 1618419204
transform 1 0 9108 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_95
timestamp 1618419204
transform 1 0 9844 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1618419204
transform -1 0 12512 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_107
timestamp 1618419204
transform 1 0 10948 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_124
timestamp 1618419204
transform 1 0 12512 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1618419204
transform 1 0 14720 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1618419204
transform 1 0 13616 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1618419204
transform -1 0 13248 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1618419204
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_128
timestamp 1618419204
transform 1 0 12880 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_132
timestamp 1618419204
transform 1 0 13248 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_139
timestamp 1618419204
transform 1 0 13892 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_144
timestamp 1618419204
transform 1 0 14352 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1618419204
transform -1 0 16652 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_157
timestamp 1618419204
transform 1 0 15548 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_169
timestamp 1618419204
transform 1 0 16652 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1618419204
transform -1 0 19044 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1618419204
transform 1 0 18124 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_181
timestamp 1618419204
transform 1 0 17756 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_188
timestamp 1618419204
transform 1 0 18400 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb0
timestamp 1618419204
transform 1 0 1748 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1618419204
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1618419204
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_14
timestamp 1618419204
transform 1 0 2392 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 5980 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 3772 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_9_26
timestamp 1618419204
transform 1 0 3496 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_35
timestamp 1618419204
transform 1 0 4324 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_43
timestamp 1618419204
transform 1 0 5060 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_8  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 8280 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1618419204
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_53
timestamp 1618419204
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_58
timestamp 1618419204
transform 1 0 6440 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1618419204
transform 1 0 8648 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_78
timestamp 1618419204
transform 1 0 8280 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_85
timestamp 1618419204
transform 1 0 8924 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_97
timestamp 1618419204
transform 1 0 10028 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0
timestamp 1618419204
transform 1 0 10764 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1618419204
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_109
timestamp 1618419204
transform 1 0 11132 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1618419204
transform 1 0 11500 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_115
timestamp 1618419204
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb1
timestamp 1618419204
transform 1 0 12788 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_9_134
timestamp 1618419204
transform 1 0 13432 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_146
timestamp 1618419204
transform 1 0 14536 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb0
timestamp 1618419204
transform 1 0 15732 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1618419204
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_158
timestamp 1618419204
transform 1 0 15640 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_166
timestamp 1618419204
transform 1 0 16376 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_170
timestamp 1618419204
transform 1 0 16744 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_172
timestamp 1618419204
transform 1 0 16928 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1618419204
transform -1 0 19044 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_184
timestamp 1618419204
transform 1 0 18032 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1618419204
transform -1 0 2760 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1618419204
transform 1 0 3128 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1618419204
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1618419204
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_18
timestamp 1618419204
transform 1 0 2760 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _354_
timestamp 1618419204
transform -1 0 5060 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1618419204
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_25
timestamp 1618419204
transform 1 0 3404 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_30
timestamp 1618419204
transform 1 0 3864 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_43
timestamp 1618419204
transform 1 0 5060 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 7544 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_10_55
timestamp 1618419204
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_70
timestamp 1618419204
transform 1 0 7544 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_1  _306_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 9476 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1618419204
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_82
timestamp 1618419204
transform 1 0 8648 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1618419204
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_96
timestamp 1618419204
transform 1 0 9936 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 10948 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1618419204
transform -1 0 12052 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_104
timestamp 1618419204
transform 1 0 10672 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_112
timestamp 1618419204
transform 1 0 11408 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_119
timestamp 1618419204
transform 1 0 12052 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen1
timestamp 1618419204
transform 1 0 12880 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1618419204
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_127
timestamp 1618419204
transform 1 0 12788 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_133
timestamp 1618419204
transform 1 0 13340 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1618419204
transform 1 0 14076 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_144
timestamp 1618419204
transform 1 0 14352 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen0
timestamp 1618419204
transform 1 0 16376 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_10_156
timestamp 1618419204
transform 1 0 15456 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_164
timestamp 1618419204
transform 1 0 16192 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_171
timestamp 1618419204
transform 1 0 16836 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1618419204
transform -1 0 17664 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1618419204
transform -1 0 19044 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_180
timestamp 1618419204
transform 1 0 17664 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen1
timestamp 1618419204
transform -1 0 3128 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb1
timestamp 1618419204
transform 1 0 1656 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1618419204
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1618419204
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_13
timestamp 1618419204
transform 1 0 2300 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_22
timestamp 1618419204
transform 1 0 3128 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1618419204
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _377_
timestamp 1618419204
transform -1 0 4600 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_28
timestamp 1618419204
transform 1 0 3680 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_38
timestamp 1618419204
transform 1 0 4600 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 7176 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1618419204
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_53
timestamp 1618419204
transform 1 0 5980 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_58
timestamp 1618419204
transform 1 0 6440 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_66
timestamp 1618419204
transform 1 0 7176 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_74
timestamp 1618419204
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_1  _312_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 9844 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1618419204
transform 1 0 8096 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_85
timestamp 1618419204
transform 1 0 8924 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_95
timestamp 1618419204
transform 1 0 9844 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen1
timestamp 1618419204
transform -1 0 12512 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb1
timestamp 1618419204
transform 1 0 10580 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1618419204
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_110
timestamp 1618419204
transform 1 0 11224 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115
timestamp 1618419204
transform 1 0 11684 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_124
timestamp 1618419204
transform 1 0 12512 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 1618419204
transform 1 0 12880 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb0
timestamp 1618419204
transform 1 0 14444 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_11_131
timestamp 1618419204
transform 1 0 13156 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_143
timestamp 1618419204
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen0
timestamp 1618419204
transform 1 0 15456 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1618419204
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_152
timestamp 1618419204
transform 1 0 15088 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_161
timestamp 1618419204
transform 1 0 15916 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1618419204
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_172
timestamp 1618419204
transform 1 0 16928 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb1
timestamp 1618419204
transform 1 0 17296 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1618419204
transform -1 0 19044 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_183
timestamp 1618419204
transform 1 0 17940 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_191
timestamp 1618419204
transform 1 0 18676 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _314_
timestamp 1618419204
transform 1 0 2852 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1618419204
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output39
timestamp 1618419204
transform -1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_7
timestamp 1618419204
transform 1 0 1748 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 4876 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1618419204
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_25
timestamp 1618419204
transform 1 0 3404 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_30
timestamp 1618419204
transform 1 0 3864 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_38
timestamp 1618419204
transform 1 0 4600 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_48
timestamp 1618419204
transform 1 0 5520 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1618419204
transform 1 0 5888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1618419204
transform 1 0 7268 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 6532 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_55
timestamp 1618419204
transform 1 0 6164 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_63
timestamp 1618419204
transform 1 0 6900 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_70
timestamp 1618419204
transform 1 0 7544 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 9476 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _319_
timestamp 1618419204
transform 1 0 8096 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1618419204
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_82
timestamp 1618419204
transform 1 0 8648 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1618419204
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_96
timestamp 1618419204
transform 1 0 9936 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1618419204
transform -1 0 11776 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb0
timestamp 1618419204
transform -1 0 13156 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_12_104
timestamp 1618419204
transform 1 0 10672 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_116
timestamp 1618419204
transform 1 0 11776 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1618419204
transform 1 0 14720 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1618419204
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_131
timestamp 1618419204
transform 1 0 13156 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_144
timestamp 1618419204
transform 1 0 14352 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1618419204
transform 1 0 15548 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1618419204
transform 1 0 16376 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_152
timestamp 1618419204
transform 1 0 15088 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_156
timestamp 1618419204
transform 1 0 15456 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_160
timestamp 1618419204
transform 1 0 15824 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1618419204
transform 1 0 16744 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1618419204
transform 1 0 18032 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen1
timestamp 1618419204
transform 1 0 17204 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1618419204
transform -1 0 19044 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_174
timestamp 1618419204
transform 1 0 17112 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_180
timestamp 1618419204
transform 1 0 17664 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_187
timestamp 1618419204
transform 1 0 18308 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_191
timestamp 1618419204
transform 1 0 18676 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_11
timestamp 1618419204
transform 1 0 2116 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1618419204
transform 1 0 1380 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1618419204
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1618419204
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1618419204
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb1
timestamp 1618419204
transform 1 0 2208 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1618419204
transform -1 0 2300 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp 1618419204
transform 1 0 2852 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_13
timestamp 1618419204
transform 1 0 2300 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1618419204
transform -1 0 3036 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_21
timestamp 1618419204
transform 1 0 3036 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_30
timestamp 1618419204
transform 1 0 3864 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1618419204
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_33
timestamp 1618419204
transform 1 0 4140 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1618419204
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _366_
timestamp 1618419204
transform 1 0 4232 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_43
timestamp 1618419204
transform 1 0 5060 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_43
timestamp 1618419204
transform 1 0 5060 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _308_
timestamp 1618419204
transform 1 0 4416 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _304_
timestamp 1618419204
transform 1 0 5428 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _296_
timestamp 1618419204
transform -1 0 5888 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_14_58
timestamp 1618419204
transform 1 0 6440 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_54
timestamp 1618419204
transform 1 0 6072 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_58
timestamp 1618419204
transform 1 0 6440 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_56
timestamp 1618419204
transform 1 0 6256 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1618419204
transform 1 0 5888 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1618419204
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_63
timestamp 1618419204
transform 1 0 6900 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_64
timestamp 1618419204
transform 1 0 6992 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _302_
timestamp 1618419204
transform 1 0 7268 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _300_
timestamp 1618419204
transform -1 0 6900 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _298_
timestamp 1618419204
transform -1 0 7728 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_14_71
timestamp 1618419204
transform 1 0 7636 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_72
timestamp 1618419204
transform 1 0 7728 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1618419204
transform 1 0 8924 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_81
timestamp 1618419204
transform 1 0 8556 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_75
timestamp 1618419204
transform 1 0 8004 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_86
timestamp 1618419204
transform 1 0 9016 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1618419204
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _321_
timestamp 1618419204
transform 1 0 8464 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _310_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 8556 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_14_97
timestamp 1618419204
transform 1 0 10028 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_87
timestamp 1618419204
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _317_
timestamp 1618419204
transform -1 0 10028 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1618419204
transform 1 0 9384 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1618419204
transform 1 0 9660 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _347_
timestamp 1618419204
transform -1 0 12512 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _365_
timestamp 1618419204
transform 1 0 10764 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1618419204
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_105
timestamp 1618419204
transform 1 0 10764 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1618419204
transform 1 0 11500 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_115
timestamp 1618419204
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_114
timestamp 1618419204
transform 1 0 11592 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_120
timestamp 1618419204
transform 1 0 12144 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_124
timestamp 1618419204
transform 1 0 12512 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _357_
timestamp 1618419204
transform 1 0 12880 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen0
timestamp 1618419204
transform -1 0 13340 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1618419204
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_127
timestamp 1618419204
transform 1 0 12788 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_133
timestamp 1618419204
transform 1 0 13340 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_145
timestamp 1618419204
transform 1 0 14444 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_137
timestamp 1618419204
transform 1 0 13708 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_144
timestamp 1618419204
transform 1 0 14352 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_161
timestamp 1618419204
transform 1 0 15916 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_156
timestamp 1618419204
transform 1 0 15456 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen1
timestamp 1618419204
transform 1 0 14996 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1618419204
transform 1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp 1618419204
transform 1 0 15088 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_169
timestamp 1618419204
transform 1 0 16652 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_163
timestamp 1618419204
transform 1 0 16100 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1618419204
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _373_
timestamp 1618419204
transform -1 0 17572 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1618419204
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1618419204
transform -1 0 19044 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1618419204
transform -1 0 19044 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1618419204
transform 1 0 18124 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_184
timestamp 1618419204
transform 1 0 18032 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_188
timestamp 1618419204
transform 1 0 18400 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_179
timestamp 1618419204
transform 1 0 17572 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_191
timestamp 1618419204
transform 1 0 18676 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1618419204
transform 1 0 3220 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen1
timestamp 1618419204
transform 1 0 2392 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1618419204
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1618419204
transform 1 0 1380 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_11
timestamp 1618419204
transform 1 0 2116 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_19
timestamp 1618419204
transform 1 0 2852 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _248_
timestamp 1618419204
transform 1 0 4600 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_15_26
timestamp 1618419204
transform 1 0 3496 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_43
timestamp 1618419204
transform 1 0 5060 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_49
timestamp 1618419204
transform 1 0 5612 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1618419204
transform 1 0 5704 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _254_
timestamp 1618419204
transform 1 0 6808 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1618419204
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_53
timestamp 1618419204
transform 1 0 5980 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_58
timestamp 1618419204
transform 1 0 6440 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_69
timestamp 1618419204
transform 1 0 7452 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 8280 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 10304 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_77
timestamp 1618419204
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_87
timestamp 1618419204
transform 1 0 9108 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _290_
timestamp 1618419204
transform 1 0 10672 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 12512 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1618419204
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_100
timestamp 1618419204
transform 1 0 10304 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_109
timestamp 1618419204
transform 1 0 11132 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1618419204
transform 1 0 11500 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_115
timestamp 1618419204
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_124
timestamp 1618419204
transform 1 0 12512 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1618419204
transform 1 0 12972 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb1
timestamp 1618419204
transform 1 0 14812 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_15_128
timestamp 1618419204
transform 1 0 12880 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_138
timestamp 1618419204
transform 1 0 13800 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_146
timestamp 1618419204
transform 1 0 14536 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1618419204
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_156
timestamp 1618419204
transform 1 0 15456 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_168
timestamp 1618419204
transform 1 0 16560 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_172
timestamp 1618419204
transform 1 0 16928 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1618419204
transform -1 0 19044 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1618419204
transform -1 0 18400 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_184
timestamp 1618419204
transform 1 0 18032 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_188
timestamp 1618419204
transform 1 0 18400 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1618419204
transform 1 0 2760 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1618419204
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output40
timestamp 1618419204
transform -1 0 1748 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_7
timestamp 1618419204
transform 1 0 1748 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_15
timestamp 1618419204
transform 1 0 2484 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_21
timestamp 1618419204
transform 1 0 3036 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1618419204
transform -1 0 5336 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _293_
timestamp 1618419204
transform -1 0 4692 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1618419204
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_30
timestamp 1618419204
transform 1 0 3864 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_39
timestamp 1618419204
transform 1 0 4692 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_46
timestamp 1618419204
transform 1 0 5336 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1618419204
transform 1 0 7544 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1618419204
transform 1 0 6900 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _294_
timestamp 1618419204
transform 1 0 6072 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_16_59
timestamp 1618419204
transform 1 0 6532 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_66
timestamp 1618419204
transform 1 0 7176 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_73
timestamp 1618419204
transform 1 0 7820 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _309_
timestamp 1618419204
transform 1 0 8188 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1618419204
transform -1 0 10672 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1618419204
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_82
timestamp 1618419204
transform 1 0 8648 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_87
timestamp 1618419204
transform 1 0 9108 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _292_
timestamp 1618419204
transform 1 0 12420 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _371_
timestamp 1618419204
transform -1 0 11868 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_104
timestamp 1618419204
transform 1 0 10672 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_117
timestamp 1618419204
transform 1 0 11868 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1618419204
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_128
timestamp 1618419204
transform 1 0 12880 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_140
timestamp 1618419204
transform 1 0 13984 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_144
timestamp 1618419204
transform 1 0 14352 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _385_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 16100 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_16_156
timestamp 1618419204
transform 1 0 15456 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_162
timestamp 1618419204
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1618419204
transform -1 0 19044 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_184
timestamp 1618419204
transform 1 0 18032 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _364_
timestamp 1618419204
transform -1 0 2300 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen0
timestamp 1618419204
transform 1 0 2668 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1618419204
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1618419204
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1618419204
transform 1 0 2300 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_22
timestamp 1618419204
transform 1 0 3128 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _305_
timestamp 1618419204
transform 1 0 4508 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1618419204
transform 1 0 5520 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_34
timestamp 1618419204
transform 1 0 4232 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_44
timestamp 1618419204
transform 1 0 5152 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _394_
timestamp 1618419204
transform 1 0 6808 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1618419204
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_51
timestamp 1618419204
transform 1 0 5796 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_58
timestamp 1618419204
transform 1 0 6440 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _320_
timestamp 1618419204
transform -1 0 9936 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_83
timestamp 1618419204
transform 1 0 8740 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_96
timestamp 1618419204
transform 1 0 9936 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 10580 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1618419204
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_102
timestamp 1618419204
transform 1 0 10488 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_106
timestamp 1618419204
transform 1 0 10856 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_115
timestamp 1618419204
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1618419204
transform 1 0 13340 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _386_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 14168 0 1 11424
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_6  FILLER_17_127
timestamp 1618419204
transform 1 0 12788 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_136
timestamp 1618419204
transform 1 0 13616 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1618419204
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_165
timestamp 1618419204
transform 1 0 16284 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_172
timestamp 1618419204
transform 1 0 16928 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1618419204
transform 1 0 17940 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1618419204
transform 1 0 17296 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1618419204
transform -1 0 19044 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1618419204
transform 1 0 17572 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_186
timestamp 1618419204
transform 1 0 18216 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb0
timestamp 1618419204
transform 1 0 1748 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1618419204
transform 1 0 2852 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1618419204
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1618419204
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_14
timestamp 1618419204
transform 1 0 2392 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_18
timestamp 1618419204
transform 1 0 2760 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_23
timestamp 1618419204
transform 1 0 3220 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_2  _392_
timestamp 1618419204
transform 1 0 4232 0 -1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1618419204
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_30
timestamp 1618419204
transform 1 0 3864 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1618419204
transform 1 0 6532 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp 1618419204
transform -1 0 7728 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_55
timestamp 1618419204
transform 1 0 6164 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_62
timestamp 1618419204
transform 1 0 6808 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_68
timestamp 1618419204
transform 1 0 7360 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_72
timestamp 1618419204
transform 1 0 7728 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1618419204
transform -1 0 8556 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _258_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 9476 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1618419204
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_81
timestamp 1618419204
transform 1 0 8556 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1618419204
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1618419204
transform 1 0 9108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1618419204
transform 1 0 10120 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1618419204
transform 1 0 10488 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1618419204
transform -1 0 11408 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _401_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 12052 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_18_105
timestamp 1618419204
transform 1 0 10764 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_112
timestamp 1618419204
transform 1 0 11408 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_118
timestamp 1618419204
transform 1 0 11960 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1618419204
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_139
timestamp 1618419204
transform 1 0 13892 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_144
timestamp 1618419204
transform 1 0 14352 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _341_
timestamp 1618419204
transform -1 0 15364 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _400_
timestamp 1618419204
transform 1 0 16560 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_18_155
timestamp 1618419204
transform 1 0 15364 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_167
timestamp 1618419204
transform 1 0 16468 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1618419204
transform -1 0 19044 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_188
timestamp 1618419204
transform 1 0 18400 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1618419204
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1618419204
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1618419204
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1618419204
transform 1 0 1472 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1618419204
transform 1 0 3312 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_13
timestamp 1618419204
transform 1 0 2300 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_21
timestamp 1618419204
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_15
timestamp 1618419204
transform 1 0 2484 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb1
timestamp 1618419204
transform -1 0 3312 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1618419204
transform 1 0 3128 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1618419204
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_30
timestamp 1618419204
transform 1 0 3864 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_28
timestamp 1618419204
transform 1 0 3680 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_37
timestamp 1618419204
transform 1 0 4508 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1618419204
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_44
timestamp 1618419204
transform 1 0 5152 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_38
timestamp 1618419204
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_43
timestamp 1618419204
transform 1 0 5060 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _273_
timestamp 1618419204
transform -1 0 5152 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1618419204
transform 1 0 5520 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _246_
timestamp 1618419204
transform 1 0 5152 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_19_25
timestamp 1618419204
transform 1 0 3404 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_58
timestamp 1618419204
transform 1 0 6440 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_51
timestamp 1618419204
transform 1 0 5796 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1618419204
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_68
timestamp 1618419204
transform 1 0 7360 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_63
timestamp 1618419204
transform 1 0 6900 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_66
timestamp 1618419204
transform 1 0 7176 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _266_
timestamp 1618419204
transform -1 0 7360 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1618419204
transform 1 0 7728 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _252_
timestamp 1618419204
transform -1 0 8096 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_20_51
timestamp 1618419204
transform 1 0 5796 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_83
timestamp 1618419204
transform 1 0 8740 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_75
timestamp 1618419204
transform 1 0 8004 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_76
timestamp 1618419204
transform 1 0 8096 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1618419204
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _363_
timestamp 1618419204
transform 1 0 8832 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_94
timestamp 1618419204
transform 1 0 9752 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_87
timestamp 1618419204
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_93
timestamp 1618419204
transform 1 0 9660 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1618419204
transform 1 0 9476 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _395_
timestamp 1618419204
transform 1 0 10120 0 -1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1618419204
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_4  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 11224 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_19_115
timestamp 1618419204
transform 1 0 11684 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_110
timestamp 1618419204
transform 1 0 11224 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1618419204
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_123
timestamp 1618419204
transform 1 0 12420 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_119
timestamp 1618419204
transform 1 0 12052 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_123
timestamp 1618419204
transform 1 0 12420 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 12512 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 13156 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 13616 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _279_
timestamp 1618419204
transform -1 0 15180 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _285_
timestamp 1618419204
transform -1 0 15180 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1618419204
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_131
timestamp 1618419204
transform 1 0 13156 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_143
timestamp 1618419204
transform 1 0 14260 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_132
timestamp 1618419204
transform 1 0 13248 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_139
timestamp 1618419204
transform 1 0 13892 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_144
timestamp 1618419204
transform 1 0 14352 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_153
timestamp 1618419204
transform 1 0 15180 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1618419204
transform 1 0 15180 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 16376 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1618419204
transform -1 0 15824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_166
timestamp 1618419204
transform 1 0 16376 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_168
timestamp 1618419204
transform 1 0 16560 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp 1618419204
transform 1 0 15824 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_173
timestamp 1618419204
transform 1 0 17020 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_172
timestamp 1618419204
transform 1 0 16928 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1618419204
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1618419204
transform -1 0 17020 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _200_
timestamp 1618419204
transform -1 0 17940 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _209_
timestamp 1618419204
transform 1 0 17480 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1618419204
transform -1 0 19044 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1618419204
transform -1 0 19044 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_183
timestamp 1618419204
transform 1 0 17940 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_191
timestamp 1618419204
transform 1 0 18676 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_177
timestamp 1618419204
transform 1 0 17388 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_186
timestamp 1618419204
transform 1 0 18216 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1618419204
transform 1 0 2024 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen1
timestamp 1618419204
transform -1 0 3496 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1618419204
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1618419204
transform -1 0 1656 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_6
timestamp 1618419204
transform 1 0 1656 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_17
timestamp 1618419204
transform 1 0 2668 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1618419204
transform -1 0 4324 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 5428 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_26
timestamp 1618419204
transform 1 0 3496 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_35
timestamp 1618419204
transform 1 0 4324 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1618419204
transform 1 0 5428 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _265_
timestamp 1618419204
transform -1 0 7728 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1618419204
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_55
timestamp 1618419204
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_58
timestamp 1618419204
transform 1 0 6440 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_72
timestamp 1618419204
transform 1 0 7728 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1618419204
transform 1 0 8096 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _260_
timestamp 1618419204
transform 1 0 8924 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _261_
timestamp 1618419204
transform -1 0 10396 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_79
timestamp 1618419204
transform 1 0 8372 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_93
timestamp 1618419204
transform 1 0 9660 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1618419204
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_101
timestamp 1618419204
transform 1 0 10396 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1618419204
transform 1 0 11500 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_115
timestamp 1618419204
transform 1 0 11684 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1618419204
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_1  _223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 13708 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 12604 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _286_
timestamp 1618419204
transform 1 0 14720 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_21_133
timestamp 1618419204
transform 1 0 13340 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_141
timestamp 1618419204
transform 1 0 14076 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_147
timestamp 1618419204
transform 1 0 14628 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _288_
timestamp 1618419204
transform 1 0 15916 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1618419204
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_155
timestamp 1618419204
transform 1 0 15364 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_166
timestamp 1618419204
transform 1 0 16376 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_170
timestamp 1618419204
transform 1 0 16744 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_172
timestamp 1618419204
transform 1 0 16928 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _210_
timestamp 1618419204
transform 1 0 17296 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1618419204
transform -1 0 19044 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_183
timestamp 1618419204
transform 1 0 17940 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_191
timestamp 1618419204
transform 1 0 18676 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb0
timestamp 1618419204
transform 1 0 1472 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1618419204
transform -1 0 3128 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1618419204
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1618419204
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_11
timestamp 1618419204
transform 1 0 2116 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_22
timestamp 1618419204
transform 1 0 3128 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 5888 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _270_
timestamp 1618419204
transform -1 0 4784 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1618419204
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_28
timestamp 1618419204
transform 1 0 3680 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_30
timestamp 1618419204
transform 1 0 3864 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_40
timestamp 1618419204
transform 1 0 4784 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _256_
timestamp 1618419204
transform -1 0 8372 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _263_
timestamp 1618419204
transform 1 0 6900 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_52
timestamp 1618419204
transform 1 0 5888 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_60
timestamp 1618419204
transform 1 0 6624 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_67
timestamp 1618419204
transform 1 0 7268 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1618419204
transform 1 0 9476 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1618419204
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_79
timestamp 1618419204
transform 1 0 8372 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1618419204
transform 1 0 8924 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_87
timestamp 1618419204
transform 1 0 9108 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1618419204
transform 1 0 9752 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__o2bb2a_1  _220_
timestamp 1618419204
transform 1 0 10948 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_106
timestamp 1618419204
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_115
timestamp 1618419204
transform 1 0 11684 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1618419204
transform -1 0 13432 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1618419204
transform -1 0 15088 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1618419204
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_127
timestamp 1618419204
transform 1 0 12788 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_134
timestamp 1618419204
transform 1 0 13432 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_142
timestamp 1618419204
transform 1 0 14168 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_144
timestamp 1618419204
transform 1 0 14352 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_148
timestamp 1618419204
transform 1 0 14720 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1618419204
transform 1 0 16100 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 17388 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_22_152
timestamp 1618419204
transform 1 0 15088 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_160
timestamp 1618419204
transform 1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_166
timestamp 1618419204
transform 1 0 16376 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1618419204
transform -1 0 19044 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1618419204
transform -1 0 18400 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_177
timestamp 1618419204
transform 1 0 17388 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_188
timestamp 1618419204
transform 1 0 18400 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1618419204
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1618419204
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1618419204
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _244_
timestamp 1618419204
transform 1 0 4692 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1618419204
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_46
timestamp 1618419204
transform 1 0 5336 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1618419204
transform 1 0 5704 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _251_
timestamp 1618419204
transform 1 0 7268 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1618419204
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_53
timestamp 1618419204
transform 1 0 5980 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_58
timestamp 1618419204
transform 1 0 6440 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_66
timestamp 1618419204
transform 1 0 7176 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_74
timestamp 1618419204
transform 1 0 7912 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 10396 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _262_
timestamp 1618419204
transform 1 0 8280 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_23_83
timestamp 1618419204
transform 1 0 8740 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_91
timestamp 1618419204
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_1  _219_
timestamp 1618419204
transform 1 0 12052 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _221_
timestamp 1618419204
transform -1 0 11224 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1618419204
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_101
timestamp 1618419204
transform 1 0 10396 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_110
timestamp 1618419204
transform 1 0 11224 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_115
timestamp 1618419204
transform 1 0 11684 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 14444 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1618419204
transform 1 0 12604 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_137
timestamp 1618419204
transform 1 0 13708 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1618419204
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_152
timestamp 1618419204
transform 1 0 15088 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_164
timestamp 1618419204
transform 1 0 16192 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_170
timestamp 1618419204
transform 1 0 16744 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_172
timestamp 1618419204
transform 1 0 16928 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _208_
timestamp 1618419204
transform 1 0 17296 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1618419204
transform 1 0 18124 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1618419204
transform -1 0 19044 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_181
timestamp 1618419204
transform 1 0 17756 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_188
timestamp 1618419204
transform 1 0 18400 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1618419204
transform -1 0 3036 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1618419204
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1618419204
transform -1 0 1656 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_6
timestamp 1618419204
transform 1 0 1656 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_21
timestamp 1618419204
transform 1 0 3036 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _269_
timestamp 1618419204
transform -1 0 5796 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 4232 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1618419204
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_30
timestamp 1618419204
transform 1 0 3864 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_42
timestamp 1618419204
transform 1 0 4968 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1618419204
transform 1 0 6164 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _267_
timestamp 1618419204
transform -1 0 7728 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_51
timestamp 1618419204
transform 1 0 5796 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_58
timestamp 1618419204
transform 1 0 6440 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_66
timestamp 1618419204
transform 1 0 7176 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_72
timestamp 1618419204
transform 1 0 7728 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_1  _237_
timestamp 1618419204
transform 1 0 9660 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1618419204
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1618419204
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_87
timestamp 1618419204
transform 1 0 9108 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_98
timestamp 1618419204
transform 1 0 10120 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _213_
timestamp 1618419204
transform -1 0 11592 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _402_
timestamp 1618419204
transform -1 0 13800 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_24_114
timestamp 1618419204
transform 1 0 11592 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _384_
timestamp 1618419204
transform 1 0 14720 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1618419204
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_138
timestamp 1618419204
transform 1 0 13800 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_142
timestamp 1618419204
transform 1 0 14168 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_144
timestamp 1618419204
transform 1 0 14352 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _201_
timestamp 1618419204
transform -1 0 17572 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_24_168
timestamp 1618419204
transform 1 0 16560 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1618419204
transform -1 0 18216 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1618419204
transform -1 0 19044 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_179
timestamp 1618419204
transform 1 0 17572 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_186
timestamp 1618419204
transform 1 0 18216 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_2  _391_
timestamp 1618419204
transform 1 0 1840 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1618419204
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1618419204
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1618419204
transform 1 0 1748 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _274_
timestamp 1618419204
transform -1 0 5060 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_25_29
timestamp 1618419204
transform 1 0 3772 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_37
timestamp 1618419204
transform 1 0 4508 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_43
timestamp 1618419204
transform 1 0 5060 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_49
timestamp 1618419204
transform 1 0 5612 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1618419204
transform 1 0 5704 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _268_
timestamp 1618419204
transform 1 0 6900 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1618419204
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_53
timestamp 1618419204
transform 1 0 5980 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_58
timestamp 1618419204
transform 1 0 6440 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_62
timestamp 1618419204
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_71
timestamp 1618419204
transform 1 0 7636 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1618419204
transform 1 0 8556 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_2  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 10304 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_79
timestamp 1618419204
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_84
timestamp 1618419204
transform 1 0 8832 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _198_
timestamp 1618419204
transform 1 0 12052 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1618419204
transform -1 0 10948 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1618419204
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_100
timestamp 1618419204
transform 1 0 10304 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_107
timestamp 1618419204
transform 1 0 10948 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1618419204
transform 1 0 11500 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_115
timestamp 1618419204
transform 1 0 11684 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _289_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 14996 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_126
timestamp 1618419204
transform 1 0 12696 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_138
timestamp 1618419204
transform 1 0 13800 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_142
timestamp 1618419204
transform 1 0 14168 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _343_
timestamp 1618419204
transform -1 0 15640 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1618419204
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1618419204
transform -1 0 16468 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_151
timestamp 1618419204
transform 1 0 14996 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_158
timestamp 1618419204
transform 1 0 15640 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_167
timestamp 1618419204
transform 1 0 16468 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_172
timestamp 1618419204
transform 1 0 16928 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _227_
timestamp 1618419204
transform 1 0 17296 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1618419204
transform -1 0 19044 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_182
timestamp 1618419204
transform 1 0 17848 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_190
timestamp 1618419204
transform 1 0 18584 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _390_
timestamp 1618419204
transform 1 0 1564 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1618419204
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1618419204
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1618419204
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1618419204
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1618419204
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_25
timestamp 1618419204
transform 1 0 3404 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_30
timestamp 1618419204
transform 1 0 3864 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1618419204
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1618419204
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_1  _277_
timestamp 1618419204
transform 1 0 3772 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_37
timestamp 1618419204
transform 1 0 4508 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_38
timestamp 1618419204
transform 1 0 4600 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _242_
timestamp 1618419204
transform -1 0 5060 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _240_
timestamp 1618419204
transform -1 0 5520 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1618419204
transform 1 0 5520 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_43
timestamp 1618419204
transform 1 0 5060 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1618419204
transform 1 0 5428 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_58
timestamp 1618419204
transform 1 0 6440 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_56
timestamp 1618419204
transform 1 0 6256 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_58
timestamp 1618419204
transform 1 0 6440 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_50
timestamp 1618419204
transform 1 0 5704 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1618419204
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _241_
timestamp 1618419204
transform -1 0 7084 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_65
timestamp 1618419204
transform 1 0 7084 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1618419204
transform -1 0 7728 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_72
timestamp 1618419204
transform 1 0 7728 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _393_
timestamp 1618419204
transform 1 0 6532 0 -1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__a41o_2  _234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 9292 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_4  _238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 9476 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1618419204
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_80
timestamp 1618419204
transform 1 0 8464 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1618419204
transform 1 0 9108 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_84
timestamp 1618419204
transform 1 0 8832 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_88
timestamp 1618419204
transform 1 0 9200 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_98
timestamp 1618419204
transform 1 0 10120 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_106
timestamp 1618419204
transform 1 0 10856 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_108
timestamp 1618419204
transform 1 0 11040 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _236_
timestamp 1618419204
transform -1 0 10856 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_115
timestamp 1618419204
transform 1 0 11684 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_26_116
timestamp 1618419204
transform 1 0 11776 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1618419204
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _206_
timestamp 1618419204
transform -1 0 12328 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1618419204
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_122
timestamp 1618419204
transform 1 0 12328 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _283_
timestamp 1618419204
transform 1 0 12328 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1618419204
transform -1 0 13616 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _387_
timestamp 1618419204
transform 1 0 13524 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1618419204
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_130
timestamp 1618419204
transform 1 0 13064 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_136
timestamp 1618419204
transform 1 0 13616 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_142
timestamp 1618419204
transform 1 0 14168 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_144
timestamp 1618419204
transform 1 0 14352 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_131
timestamp 1618419204
transform 1 0 13156 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_156
timestamp 1618419204
transform 1 0 15456 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_157
timestamp 1618419204
transform 1 0 15548 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_152
timestamp 1618419204
transform 1 0 15088 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__a21boi_1  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 15824 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1618419204
transform -1 0 15548 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _229_
timestamp 1618419204
transform -1 0 16192 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_172
timestamp 1618419204
transform 1 0 16928 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_170
timestamp 1618419204
transform 1 0 16744 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_166
timestamp 1618419204
transform 1 0 16376 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_164
timestamp 1618419204
transform 1 0 16192 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1618419204
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _399_
timestamp 1618419204
transform 1 0 16560 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__o221a_1  _231_
timestamp 1618419204
transform 1 0 17296 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1618419204
transform -1 0 19044 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1618419204
transform -1 0 19044 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_188
timestamp 1618419204
transform 1 0 18400 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_185
timestamp 1618419204
transform 1 0 18124 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_191
timestamp 1618419204
transform 1 0 18676 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1618419204
transform 1 0 2576 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1618419204
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1618419204
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_6
timestamp 1618419204
transform 1 0 1656 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_14
timestamp 1618419204
transform 1 0 2392 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1618419204
transform 1 0 2852 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _276_
timestamp 1618419204
transform -1 0 4692 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _398_
timestamp 1618419204
transform 1 0 5612 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1618419204
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1618419204
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_30
timestamp 1618419204
transform 1 0 3864 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_39
timestamp 1618419204
transform 1 0 4692 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_47
timestamp 1618419204
transform 1 0 5428 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_69
timestamp 1618419204
transform 1 0 7452 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1618419204
transform 1 0 9752 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1618419204
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_81
timestamp 1618419204
transform 1 0 8556 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 1618419204
transform 1 0 8924 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_87
timestamp 1618419204
transform 1 0 9108 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_93
timestamp 1618419204
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_97
timestamp 1618419204
transform 1 0 10028 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _214_
timestamp 1618419204
transform 1 0 12512 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _216_
timestamp 1618419204
transform -1 0 12144 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _218_
timestamp 1618419204
transform -1 0 10948 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_103
timestamp 1618419204
transform 1 0 10580 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_107
timestamp 1618419204
transform 1 0 10948 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_120
timestamp 1618419204
transform 1 0 12144 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1618419204
transform -1 0 13616 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp 1618419204
transform 1 0 14720 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1618419204
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_129
timestamp 1618419204
transform 1 0 12972 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_136
timestamp 1618419204
transform 1 0 13616 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_142
timestamp 1618419204
transform 1 0 14168 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_144
timestamp 1618419204
transform 1 0 14352 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _382_
timestamp 1618419204
transform 1 0 15732 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_28_151
timestamp 1618419204
transform 1 0 14996 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp 1618419204
transform 1 0 17940 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1618419204
transform -1 0 19044 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1618419204
transform 1 0 17572 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_186
timestamp 1618419204
transform 1 0 18216 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1618419204
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1618419204
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1618419204
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1618419204
transform -1 0 4968 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _278_
timestamp 1618419204
transform 1 0 3680 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_29_27
timestamp 1618419204
transform 1 0 3588 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_35
timestamp 1618419204
transform 1 0 4324 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_42
timestamp 1618419204
transform 1 0 4968 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4_2  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 7728 0 1 17952
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1618419204
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1618419204
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_54
timestamp 1618419204
transform 1 0 6072 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_58
timestamp 1618419204
transform 1 0 6440 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_65
timestamp 1618419204
transform 1 0 7084 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_71
timestamp 1618419204
transform 1 0 7636 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1618419204
transform 1 0 9016 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_82
timestamp 1618419204
transform 1 0 8648 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_89
timestamp 1618419204
transform 1 0 9292 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1618419204
transform -1 0 11224 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _215_
timestamp 1618419204
transform -1 0 12788 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1618419204
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_101
timestamp 1618419204
transform 1 0 10396 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_110
timestamp 1618419204
transform 1 0 11224 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_115
timestamp 1618419204
transform 1 0 11684 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _205_
timestamp 1618419204
transform -1 0 13800 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _383_
timestamp 1618419204
transform 1 0 14628 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_29_127
timestamp 1618419204
transform 1 0 12788 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_138
timestamp 1618419204
transform 1 0 13800 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_146
timestamp 1618419204
transform 1 0 14536 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1618419204
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_167
timestamp 1618419204
transform 1 0 16468 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_172
timestamp 1618419204
transform 1 0 16928 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1618419204
transform -1 0 19044 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output42
timestamp 1618419204
transform 1 0 18032 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_188
timestamp 1618419204
transform 1 0 18400 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _338_
timestamp 1618419204
transform -1 0 3404 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1618419204
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1618419204
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_15
timestamp 1618419204
transform 1 0 2484 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_21
timestamp 1618419204
transform 1 0 3036 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1618419204
transform -1 0 4508 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _396_
timestamp 1618419204
transform 1 0 4968 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1618419204
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_25
timestamp 1618419204
transform 1 0 3404 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_30
timestamp 1618419204
transform 1 0 3864 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_37
timestamp 1618419204
transform 1 0 4508 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_41
timestamp 1618419204
transform 1 0 4876 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _202_
timestamp 1618419204
transform -1 0 8280 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_30_62
timestamp 1618419204
transform 1 0 6808 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_70
timestamp 1618419204
transform 1 0 7544 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _403_
timestamp 1618419204
transform 1 0 9660 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1618419204
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_78
timestamp 1618419204
transform 1 0 8280 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_87
timestamp 1618419204
transform 1 0 9108 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _195_
timestamp 1618419204
transform -1 0 12512 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_30_113
timestamp 1618419204
transform 1 0 11500 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_124
timestamp 1618419204
transform 1 0 12512 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _282_
timestamp 1618419204
transform -1 0 13248 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _339_
timestamp 1618419204
transform -1 0 13892 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _381_
timestamp 1618419204
transform 1 0 14720 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1618419204
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_132
timestamp 1618419204
transform 1 0 13248 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_139
timestamp 1618419204
transform 1 0 13892 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_144
timestamp 1618419204
transform 1 0 14352 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 16928 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_168
timestamp 1618419204
transform 1 0 16560 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1618419204
transform -1 0 19044 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_188
timestamp 1618419204
transform 1 0 18400 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _349_
timestamp 1618419204
transform 1 0 1656 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _389_
timestamp 1618419204
transform 1 0 2392 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1618419204
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1618419204
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_9
timestamp 1618419204
transform 1 0 1932 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_13
timestamp 1618419204
transform 1 0 2300 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_34
timestamp 1618419204
transform 1 0 4232 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_46
timestamp 1618419204
transform 1 0 5336 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _204_
timestamp 1618419204
transform -1 0 7360 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 1618419204
transform -1 0 5980 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _397_
timestamp 1618419204
transform 1 0 7728 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1618419204
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_53
timestamp 1618419204
transform 1 0 5980 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_58
timestamp 1618419204
transform 1 0 6440 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_62
timestamp 1618419204
transform 1 0 6808 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_68
timestamp 1618419204
transform 1 0 7360 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_92
timestamp 1618419204
transform 1 0 9568 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp 1618419204
transform -1 0 10672 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1618419204
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_100
timestamp 1618419204
transform 1 0 10304 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 1618419204
transform 1 0 10672 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_112
timestamp 1618419204
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_115
timestamp 1618419204
transform 1 0 11684 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _388_
timestamp 1618419204
transform 1 0 12788 0 1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_31_148
timestamp 1618419204
transform 1 0 14720 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp 1618419204
transform -1 0 15548 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1618419204
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_157
timestamp 1618419204
transform 1 0 15548 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1618419204
transform 1 0 16652 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_172
timestamp 1618419204
transform 1 0 16928 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _345_
timestamp 1618419204
transform 1 0 17296 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1618419204
transform -1 0 19044 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1618419204
transform 1 0 17940 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1618419204
transform 1 0 17572 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_186
timestamp 1618419204
transform 1 0 18216 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1618419204
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1618419204
transform 1 0 2300 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1618419204
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output44
timestamp 1618419204
transform -1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_7
timestamp 1618419204
transform 1 0 1748 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_16
timestamp 1618419204
transform 1 0 2576 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_23
timestamp 1618419204
transform 1 0 3220 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1618419204
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1618419204
transform 1 0 4232 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1618419204
transform 1 0 5520 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_30
timestamp 1618419204
transform 1 0 3864 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_37
timestamp 1618419204
transform 1 0 4508 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_45
timestamp 1618419204
transform 1 0 5244 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _203_
timestamp 1618419204
transform 1 0 7544 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1618419204
transform 1 0 6440 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1618419204
transform 1 0 6900 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_51
timestamp 1618419204
transform 1 0 5796 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_57
timestamp 1618419204
transform 1 0 6348 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_59
timestamp 1618419204
transform 1 0 6532 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_66
timestamp 1618419204
transform 1 0 7176 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1618419204
transform 1 0 9108 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1618419204
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_77
timestamp 1618419204
transform 1 0 8188 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1618419204
transform 1 0 8924 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_88
timestamp 1618419204
transform 1 0 9200 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_92
timestamp 1618419204
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_96
timestamp 1618419204
transform 1 0 9936 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1618419204
transform 1 0 11776 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1618419204
transform -1 0 12512 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1618419204
transform -1 0 10580 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_103
timestamp 1618419204
transform 1 0 10580 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_115
timestamp 1618419204
transform 1 0 11684 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_117
timestamp 1618419204
transform 1 0 11868 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_124
timestamp 1618419204
transform 1 0 12512 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1618419204
transform 1 0 14444 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1618419204
transform 1 0 12880 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_131
timestamp 1618419204
transform 1 0 13156 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_143
timestamp 1618419204
transform 1 0 14260 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1618419204
transform 1 0 14536 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1618419204
transform 1 0 14904 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1618419204
transform -1 0 16744 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1618419204
transform 1 0 15640 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_153
timestamp 1618419204
transform 1 0 15180 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_157
timestamp 1618419204
transform 1 0 15548 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_161
timestamp 1618419204
transform 1 0 15916 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_170
timestamp 1618419204
transform 1 0 16744 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1618419204
transform -1 0 19044 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1618419204
transform 1 0 17112 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1618419204
transform -1 0 18400 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_175
timestamp 1618419204
transform 1 0 17204 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_183
timestamp 1618419204
transform 1 0 17940 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_188
timestamp 1618419204
transform 1 0 18400 0 -1 20128
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 8848 800 8968 6 clockc
port 0 nsew signal tristate
rlabel metal3 s 0 11568 800 11688 6 clockd[0]
port 1 nsew signal tristate
rlabel metal3 s 0 4768 800 4888 6 clockd[1]
port 2 nsew signal tristate
rlabel metal3 s 19396 18368 20196 18488 6 clockd[2]
port 3 nsew signal tristate
rlabel metal2 s 17958 0 18014 800 6 clockd[3]
port 4 nsew signal tristate
rlabel metal3 s 0 20408 800 20528 6 clockp[0]
port 5 nsew signal tristate
rlabel metal2 s 1858 0 1914 800 6 clockp[1]
port 6 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 dco
port 7 nsew signal input
rlabel metal3 s 19396 13608 20196 13728 6 div[0]
port 8 nsew signal input
rlabel metal2 s 17498 21540 17554 22340 6 div[1]
port 9 nsew signal input
rlabel metal2 s 6918 21540 6974 22340 6 div[2]
port 10 nsew signal input
rlabel metal2 s 478 0 534 800 6 div[3]
port 11 nsew signal input
rlabel metal2 s 12898 21540 12954 22340 6 div[4]
port 12 nsew signal input
rlabel metal2 s 14278 21540 14334 22340 6 ext_trim[0]
port 13 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 ext_trim[10]
port 14 nsew signal input
rlabel metal2 s 2318 21540 2374 22340 6 ext_trim[11]
port 15 nsew signal input
rlabel metal3 s 19396 4768 20196 4888 6 ext_trim[12]
port 16 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 ext_trim[13]
port 17 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 ext_trim[14]
port 18 nsew signal input
rlabel metal3 s 19396 15648 20196 15768 6 ext_trim[15]
port 19 nsew signal input
rlabel metal2 s 3698 21540 3754 22340 6 ext_trim[16]
port 20 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 ext_trim[17]
port 21 nsew signal input
rlabel metal2 s 5538 21540 5594 22340 6 ext_trim[18]
port 22 nsew signal input
rlabel metal3 s 19396 9528 20196 9648 6 ext_trim[19]
port 23 nsew signal input
rlabel metal2 s 11518 21540 11574 22340 6 ext_trim[1]
port 24 nsew signal input
rlabel metal2 s 9678 21540 9734 22340 6 ext_trim[20]
port 25 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 ext_trim[21]
port 26 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 ext_trim[22]
port 27 nsew signal input
rlabel metal3 s 19396 20408 20196 20528 6 ext_trim[23]
port 28 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 ext_trim[24]
port 29 nsew signal input
rlabel metal2 s 8298 21540 8354 22340 6 ext_trim[25]
port 30 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 ext_trim[2]
port 31 nsew signal input
rlabel metal3 s 19396 6808 20196 6928 6 ext_trim[3]
port 32 nsew signal input
rlabel metal3 s 19396 688 20196 808 6 ext_trim[4]
port 33 nsew signal input
rlabel metal3 s 19396 11568 20196 11688 6 ext_trim[5]
port 34 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 ext_trim[6]
port 35 nsew signal input
rlabel metal2 s 938 21540 994 22340 6 ext_trim[7]
port 36 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 ext_trim[8]
port 37 nsew signal input
rlabel metal3 s 19396 2728 20196 2848 6 ext_trim[9]
port 38 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 extclk_sel
port 39 nsew signal input
rlabel metal2 s 15658 21540 15714 22340 6 osc
port 40 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 reset
port 41 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 sel[0]
port 42 nsew signal input
rlabel metal2 s 18878 21540 18934 22340 6 sel[1]
port 43 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 sel[2]
port 44 nsew signal input
rlabel metal4 s 15894 156 16214 22148 6 VPWR
port 45 nsew power bidirectional
rlabel metal4 s 9914 156 10234 22148 6 VPWR
port 46 nsew power bidirectional
rlabel metal4 s 3934 156 4254 22148 6 VPWR
port 47 nsew power bidirectional
rlabel metal4 s 20084 816 20404 21488 6 VPWR
port 48 nsew power bidirectional
rlabel metal4 s -256 816 64 21488 4 VPWR
port 49 nsew power bidirectional
rlabel metal5 s -256 21168 20404 21488 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s -916 16928 21064 17248 6 VPWR
port 51 nsew power bidirectional
rlabel metal5 s -916 10944 21064 11264 6 VPWR
port 52 nsew power bidirectional
rlabel metal5 s -916 4960 21064 5280 6 VPWR
port 53 nsew power bidirectional
rlabel metal5 s -256 816 20404 1136 6 VPWR
port 54 nsew power bidirectional
rlabel metal4 s 20744 156 21064 22148 6 VGND
port 55 nsew ground bidirectional
rlabel metal4 s 12904 156 13224 22148 6 VGND
port 56 nsew ground bidirectional
rlabel metal4 s 6924 156 7244 22148 6 VGND
port 57 nsew ground bidirectional
rlabel metal4 s -916 156 -596 22148 4 VGND
port 58 nsew ground bidirectional
rlabel metal5 s -916 21828 21064 22148 6 VGND
port 59 nsew ground bidirectional
rlabel metal5 s -916 13936 21064 14256 6 VGND
port 60 nsew ground bidirectional
rlabel metal5 s -916 7952 21064 8272 6 VGND
port 61 nsew ground bidirectional
rlabel metal5 s -916 156 21064 476 6 VGND
port 62 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20196 22340
<< end >>
