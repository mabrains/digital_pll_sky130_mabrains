* NGSPICE file created from digital_pll.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_1 abstract view
.subckt sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_2 abstract view
.subckt sky130_fd_sc_hd__einvn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvn_4 abstract view
.subckt sky130_fd_sc_hd__einvn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_4 abstract view
.subckt sky130_fd_sc_hd__einvp_4 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrbp_1 abstract view
.subckt sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_2 abstract view
.subckt sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrbp_2 abstract view
.subckt sky130_fd_sc_hd__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

.subckt digital_pll clockc clockd[0] clockd[1] clockd[2] clockd[3] clockp[0] clockp[1]
+ dco div[0] div[1] div[2] div[3] div[4] ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12]
+ ext_trim[13] ext_trim[14] ext_trim[15] ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19]
+ ext_trim[1] ext_trim[20] ext_trim[21] ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25]
+ ext_trim[2] ext_trim[3] ext_trim[4] ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8]
+ ext_trim[9] extclk_sel osc reset sel[0] sel[1] sel[2] VPWR VGND
XFILLER_22_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_363_ _320_/X _363_/A1 _376_/S VGND VGND VPWR VPWR _363_/X sky130_fd_sc_hd__mux2_2
X_294_ _294_/A _294_/B VGND VGND VPWR VPWR _309_/C sky130_fd_sc_hd__or2_1
XFILLER_13_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[1\].id.delayint0 ringosc.dstage\[1\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_346_ _348_/A VGND VGND VPWR VPWR _346_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_277_ _235_/Y _241_/Y _276_/X _390_/Q _235_/A VGND VGND VPWR VPWR _390_/D sky130_fd_sc_hd__a32o_1
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_200_ _400_/Q _284_/D _385_/Q _233_/B VGND VGND VPWR VPWR _400_/D sky130_fd_sc_hd__a22o_1
X_329_ _348_/A VGND VGND VPWR VPWR _329_/X sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[11\].id.delayen1 ringosc.dstage\[11\].id.delayen1/A _355_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[11\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[10\].id.delayenb0 ringosc.dstage\[10\].id.delayenb1/A _356_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
XFILLER_19_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[9\].id.delayenb0 ringosc.dstage\[9\].id.delayenb1/A _358_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[9\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
XFILLER_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput42 idiv8/D VGND VGND VPWR VPWR clockd[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_22_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_362_ _305_/X _362_/A1 _379_/S VGND VGND VPWR VPWR _362_/X sky130_fd_sc_hd__mux2_1
X_293_ _395_/Q _392_/Q _315_/B VGND VGND VPWR VPWR _293_/X sky130_fd_sc_hd__or3_1
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_345_ _348_/A VGND VGND VPWR VPWR _345_/X sky130_fd_sc_hd__clkbuf_1
X_276_ _389_/Q _276_/B VGND VGND VPWR VPWR _276_/X sky130_fd_sc_hd__or2_1
X_328_ _348_/A VGND VGND VPWR VPWR _328_/X sky130_fd_sc_hd__clkbuf_1
X_259_ _259_/A VGND VGND VPWR VPWR _259_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[10\].id.delayenb1 ringosc.dstage\[10\].id.delayenb1/A _357_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
Xringosc.dstage\[9\].id.delayenb1 ringosc.dstage\[9\].id.delayenb1/A _359_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[9\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput43 idiv16/D VGND VGND VPWR VPWR clockd[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_292_ _395_/Q _292_/B VGND VGND VPWR VPWR _292_/X sky130_fd_sc_hd__or2_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_361_ _314_/X _361_/A1 _379_/S VGND VGND VPWR VPWR _361_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_344_ _348_/A VGND VGND VPWR VPWR _344_/X sky130_fd_sc_hd__clkbuf_1
X_275_ _235_/Y _269_/X _274_/X _391_/Q _235_/A VGND VGND VPWR VPWR _391_/D sky130_fd_sc_hd__a32o_1
XFILLER_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[4\].id.delayen0 ringosc.dstage\[4\].id.delayen0/A _368_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XFILLER_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_258_ _395_/Q _239_/Y _313_/A _239_/A VGND VGND VPWR VPWR _259_/A sky130_fd_sc_hd__o22a_1
X_327_ _348_/A VGND VGND VPWR VPWR _327_/X sky130_fd_sc_hd__clkbuf_1
X_189_ _189_/A VGND VGND VPWR VPWR _221_/A sky130_fd_sc_hd__inv_2
XFILLER_18_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput44 _349_/X VGND VGND VPWR VPWR clockp[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[10\].id.delaybuf0 ringosc.dstage\[9\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[9\].id.delaybuf0 ringosc.dstage\[8\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[5\].id.delayenb0 ringosc.dstage\[5\].id.delayenb1/A _366_/X VGND
+ VGND VPWR VPWR ringosc.ibufp10/A sky130_fd_sc_hd__einvn_4
X_291_ _395_/Q _315_/B VGND VGND VPWR VPWR _291_/X sky130_fd_sc_hd__or2_1
XFILLER_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_360_ _303_/X _360_/A1 _379_/S VGND VGND VPWR VPWR _360_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_343_ _348_/A VGND VGND VPWR VPWR _343_/X sky130_fd_sc_hd__clkbuf_1
X_274_ _274_/A _274_/B VGND VGND VPWR VPWR _274_/X sky130_fd_sc_hd__or2_1
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[4\].id.delayen1 ringosc.dstage\[4\].id.delayen1/A _369_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[4\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_188_ _389_/Q VGND VGND VPWR VPWR _188_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_257_ _257_/A VGND VGND VPWR VPWR _257_/Y sky130_fd_sc_hd__inv_2
X_326_ _348_/A VGND VGND VPWR VPWR _326_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_309_ _309_/A _311_/C _309_/C VGND VGND VPWR VPWR _313_/B sky130_fd_sc_hd__or3_1
XFILLER_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput45 idiv2/CLK VGND VGND VPWR VPWR clockp[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_31_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[10\].id.delaybuf1 ringosc.dstage\[10\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[9\].id.delaybuf1 ringosc.dstage\[9\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[5\].id.delayenb1 ringosc.dstage\[5\].id.delayenb1/A _367_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[5\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
XFILLER_22_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_290_ _290_/A _315_/B VGND VGND VPWR VPWR _292_/B sky130_fd_sc_hd__or2_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_273_ _294_/A _235_/Y _272_/X VGND VGND VPWR VPWR _392_/D sky130_fd_sc_hd__o21ai_1
X_342_ _348_/A VGND VGND VPWR VPWR _342_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_187_ _390_/Q VGND VGND VPWR VPWR _187_/Y sky130_fd_sc_hd__inv_2
X_256_ _267_/B _253_/A _267_/A _239_/A _310_/B VGND VGND VPWR VPWR _257_/A sky130_fd_sc_hd__o32a_1
X_325_ _325_/A _325_/B _325_/C VGND VGND VPWR VPWR _350_/S sky130_fd_sc_hd__nor3_2
XFILLER_9_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_239_ _239_/A VGND VGND VPWR VPWR _239_/Y sky130_fd_sc_hd__inv_2
X_308_ _393_/Q _392_/Q _394_/Q _395_/Q VGND VGND VPWR VPWR _308_/X sky130_fd_sc_hd__a31o_1
XFILLER_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[5\].id.delaybuf0 ringosc.dstage\[4\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_272_ _247_/Y _271_/A _247_/A _271_/Y _235_/A VGND VGND VPWR VPWR _272_/X sky130_fd_sc_hd__a221o_1
X_341_ _348_/A VGND VGND VPWR VPWR _341_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[1\].id.delayenb0 ringosc.dstage\[1\].id.delayenb1/A _374_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[1\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
XFILLER_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[8\].id.delayint0 ringosc.dstage\[8\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_23_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_255_ _315_/B VGND VGND VPWR VPWR _310_/B sky130_fd_sc_hd__inv_2
X_186_ _391_/Q VGND VGND VPWR VPWR _294_/B sky130_fd_sc_hd__inv_2
XFILLER_2_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_324_ _325_/A _325_/B _324_/C VGND VGND VPWR VPWR _351_/S sky130_fd_sc_hd__nor3_2
XFILLER_18_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_238_ _218_/Y _221_/X _237_/X _236_/Y _217_/Y VGND VGND VPWR VPWR _239_/A sky130_fd_sc_hd__a41o_4
X_307_ _392_/Q _391_/Q _297_/A _299_/Y VGND VGND VPWR VPWR _307_/X sky130_fd_sc_hd__a31o_1
XFILLER_29_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[1\].id.delayenb1 ringosc.dstage\[1\].id.delayenb1/A _375_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[1\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
XFILLER_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[5\].id.delaybuf1 ringosc.dstage\[5\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_340_ _348_/A VGND VGND VPWR VPWR _340_/X sky130_fd_sc_hd__clkbuf_1
X_271_ _271_/A VGND VGND VPWR VPWR _271_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[1\].id.delayen0 ringosc.dstage\[1\].id.delayen0/A _374_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XFILLER_4_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_185_ _392_/Q VGND VGND VPWR VPWR _294_/A sky130_fd_sc_hd__inv_2
X_254_ _394_/Q _393_/Q VGND VGND VPWR VPWR _315_/B sky130_fd_sc_hd__or2_4
XFILLER_2_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_323_ _325_/A _323_/B _325_/C VGND VGND VPWR VPWR _352_/S sky130_fd_sc_hd__nor3_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_237_ _237_/A _237_/B _237_/C VGND VGND VPWR VPWR _237_/X sky130_fd_sc_hd__or3_1
X_306_ _315_/B _306_/B _395_/Q VGND VGND VPWR VPWR _306_/X sky130_fd_sc_hd__or3_1
XFILLER_29_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_270_ _294_/B _239_/A _269_/X VGND VGND VPWR VPWR _271_/A sky130_fd_sc_hd__o21ai_1
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_399_ _349_/A _399_/D _328_/X VGND VGND VPWR VPWR _399_/Q sky130_fd_sc_hd__dfrtp_1
Xringosc.dstage\[1\].id.delayen1 ringosc.dstage\[1\].id.delayen1/A _375_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[1\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_4_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[1\].id.delaybuf0 ringosc.dstage\[0\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
X_322_ _325_/A _323_/B _324_/C VGND VGND VPWR VPWR _353_/S sky130_fd_sc_hd__nor3_2
X_253_ _253_/A VGND VGND VPWR VPWR _253_/Y sky130_fd_sc_hd__inv_2
X_184_ _393_/Q VGND VGND VPWR VPWR _311_/C sky130_fd_sc_hd__inv_2
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[4\].id.delayint0 ringosc.dstage\[4\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_236_ _230_/Y _231_/X _226_/Y VGND VGND VPWR VPWR _236_/Y sky130_fd_sc_hd__o21ai_1
X_305_ _394_/Q _393_/Q _290_/A _395_/Q VGND VGND VPWR VPWR _305_/X sky130_fd_sc_hd__a31o_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_219_ _387_/Q _402_/Q _206_/Y VGND VGND VPWR VPWR _219_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.dstage\[9\].id.delayen0 ringosc.dstage\[9\].id.delayen0/A _358_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater46 _376_/S VGND VGND VPWR VPWR _379_/S sky130_fd_sc_hd__buf_8
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_398_ _349_/A _398_/D _329_/X VGND VGND VPWR VPWR _398_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[1\].id.delaybuf1 ringosc.dstage\[1\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[1\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_252_ _309_/A _239_/Y _394_/Q _239_/A VGND VGND VPWR VPWR _253_/A sky130_fd_sc_hd__o22a_1
X_183_ _394_/Q VGND VGND VPWR VPWR _309_/A sky130_fd_sc_hd__inv_2
X_321_ _315_/B _306_/B _395_/Q VGND VGND VPWR VPWR _321_/X sky130_fd_sc_hd__o21a_1
XFILLER_13_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_235_ _235_/A VGND VGND VPWR VPWR _235_/Y sky130_fd_sc_hd__inv_2
X_304_ _392_/Q _391_/Q _393_/Q _297_/A VGND VGND VPWR VPWR _304_/X sky130_fd_sc_hd__a31o_1
XFILLER_1_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_218_ _218_/A _218_/B VGND VGND VPWR VPWR _218_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput39 _353_/X VGND VGND VPWR VPWR clockc sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[9\].id.delayen1 ringosc.dstage\[9\].id.delayen1/A _359_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[9\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_397_ _349_/A _397_/D _330_/X VGND VGND VPWR VPWR _397_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_251_ _393_/Q _239_/Y _311_/C _239_/A VGND VGND VPWR VPWR _267_/B sky130_fd_sc_hd__a22o_1
X_182_ _395_/Q VGND VGND VPWR VPWR _313_/A sky130_fd_sc_hd__inv_2
X_320_ _309_/A _393_/Q _313_/A _392_/Q _315_/X VGND VGND VPWR VPWR _320_/X sky130_fd_sc_hd__o41a_1
XFILLER_18_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_234_ _218_/Y _232_/Y _226_/Y _217_/A _233_/Y VGND VGND VPWR VPWR _235_/A sky130_fd_sc_hd__a41o_2
XFILLER_24_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_303_ _391_/Q _315_/B _300_/Y VGND VGND VPWR VPWR _303_/X sky130_fd_sc_hd__a21o_1
Xringosc.dstage\[0\].id.delayint0 ringosc.dstage\[0\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.iss.reseten0 ringosc.iss.const1/HI _197_/B VGND VGND VPWR VPWR ringosc.ibufp00/A
+ sky130_fd_sc_hd__einvp_4
X_217_ _217_/A VGND VGND VPWR VPWR _217_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_396_ _349_/A _396_/D _331_/X VGND VGND VPWR VPWR _396_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_27_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[8\].id.delayenb0 ringosc.dstage\[8\].id.delayenb1/A _360_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[8\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_181_ _399_/Q VGND VGND VPWR VPWR _208_/B sky130_fd_sc_hd__inv_2
X_250_ _269_/B _247_/A _269_/A _239_/A _249_/Y VGND VGND VPWR VPWR _267_/A sky130_fd_sc_hd__o32a_1
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_379_ _321_/X _379_/A1 _379_/S VGND VGND VPWR VPWR _379_/X sky130_fd_sc_hd__mux2_1
X_233_ _397_/Q _233_/B _398_/Q _396_/Q VGND VGND VPWR VPWR _233_/Y sky130_fd_sc_hd__nand4_2
XFILLER_24_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_302_ _294_/A _297_/Y _299_/A VGND VGND VPWR VPWR _302_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_216_ _176_/Y _177_/Y _218_/A _218_/B _214_/X VGND VGND VPWR VPWR _217_/A sky130_fd_sc_hd__o221a_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xringosc.iss.delayint0 ringosc.iss.delayen1/Z VGND VGND VPWR VPWR ringosc.iss.delayen0/A
+ sky130_fd_sc_hd__clkinv_1
XFILLER_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_395_ _349_/A _395_/D _332_/X VGND VGND VPWR VPWR _395_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[8\].id.delayenb1 ringosc.dstage\[8\].id.delayenb1/A _361_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[8\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_180_ _384_/Q VGND VGND VPWR VPWR _279_/B sky130_fd_sc_hd__inv_2
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_378_ _300_/Y _378_/A1 _379_/S VGND VGND VPWR VPWR _378_/X sky130_fd_sc_hd__mux2_1
X_232_ input2/X _227_/X _231_/X VGND VGND VPWR VPWR _232_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_301_ _249_/Y _297_/Y _299_/A VGND VGND VPWR VPWR _301_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_1_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_215_ _214_/A _214_/B _214_/X VGND VGND VPWR VPWR _218_/B sky130_fd_sc_hd__a21bo_1
Xringosc.dstage\[6\].id.delayen0 ringosc.dstage\[6\].id.delayen0/A _364_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_394_ _349_/A _394_/D _333_/X VGND VGND VPWR VPWR _394_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_377_ _308_/X _377_/A1 _379_/S VGND VGND VPWR VPWR _377_/X sky130_fd_sc_hd__mux2_2
XFILLER_1_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[8\].id.delaybuf0 ringosc.dstage\[7\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[4\].id.delayenb0 ringosc.dstage\[4\].id.delayenb1/A _368_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[4\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
X_231_ _229_/A _229_/B input2/X _227_/X _230_/A VGND VGND VPWR VPWR _231_/X sky130_fd_sc_hd__o221a_1
XFILLER_24_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_300_ _311_/C _294_/A _297_/Y VGND VGND VPWR VPWR _300_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 dco VGND VGND VPWR VPWR _376_/S sky130_fd_sc_hd__buf_6
Xringosc.dstage\[10\].id.delayen0 ringosc.dstage\[10\].id.delayen0/A _356_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XFILLER_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_214_ _214_/A _214_/B VGND VGND VPWR VPWR _214_/X sky130_fd_sc_hd__or2_1
Xringosc.dstage\[6\].id.delayen1 ringosc.dstage\[6\].id.delayen1/A _365_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[6\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_393_ _349_/A _393_/D _334_/X VGND VGND VPWR VPWR _393_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_376_ _292_/X input7/X _376_/S VGND VGND VPWR VPWR _376_/X sky130_fd_sc_hd__mux2_1
Xringosc.dstage\[4\].id.delayenb1 ringosc.dstage\[4\].id.delayenb1/A _369_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[4\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
Xringosc.dstage\[8\].id.delaybuf1 ringosc.dstage\[8\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[8\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
X_230_ _230_/A VGND VGND VPWR VPWR _230_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_359_ _312_/X _359_/A1 _376_/S VGND VGND VPWR VPWR _359_/X sky130_fd_sc_hd__mux2_1
Xinput2 div[0] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__buf_1
Xringosc.dstage\[10\].id.delayen1 ringosc.dstage\[10\].id.delayen1/A _357_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[10\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_213_ _387_/Q _402_/Q _206_/Y _212_/X VGND VGND VPWR VPWR _214_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_392_ _349_/A _392_/D _335_/X VGND VGND VPWR VPWR _392_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_13_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_375_ _316_/X _375_/A1 _376_/S VGND VGND VPWR VPWR _375_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_358_ _301_/Y _358_/A1 _376_/S VGND VGND VPWR VPWR _358_/X sky130_fd_sc_hd__mux2_1
Xinput3 div[1] VGND VGND VPWR VPWR _229_/A sky130_fd_sc_hd__clkbuf_1
X_289_ _387_/Q _284_/B _388_/Q _279_/B _233_/B VGND VGND VPWR VPWR _384_/D sky130_fd_sc_hd__a311o_1
Xringosc.dstage\[4\].id.delaybuf0 ringosc.dstage\[3\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[7\].id.delayint0 ringosc.dstage\[7\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
X_212_ _386_/Q _401_/Q _207_/Y _211_/Y VGND VGND VPWR VPWR _212_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[0\].id.delayenb0 ringosc.dstage\[0\].id.delayenb1/A _376_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[0\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xirb irb/A VGND VGND VPWR VPWR irb/Y sky130_fd_sc_hd__inv_4
XFILLER_27_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_391_ _349_/A _391_/D _336_/X VGND VGND VPWR VPWR _391_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_374_ _299_/Y _374_/A1 _376_/S VGND VGND VPWR VPWR _374_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput4 div[2] VGND VGND VPWR VPWR _190_/A sky130_fd_sc_hd__buf_1
X_288_ _288_/A _288_/B VGND VGND VPWR VPWR _385_/D sky130_fd_sc_hd__or2_1
X_357_ _347_/X _357_/A1 _376_/S VGND VGND VPWR VPWR _357_/X sky130_fd_sc_hd__mux2_2
Xringosc.dstage\[3\].id.delayen0 ringosc.dstage\[3\].id.delayen0/A _370_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_211_ _211_/A VGND VGND VPWR VPWR _211_/Y sky130_fd_sc_hd__inv_2
Xringosc.dstage\[0\].id.delayenb1 ringosc.dstage\[0\].id.delayenb1/A _377_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[0\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
Xringosc.dstage\[4\].id.delaybuf1 ringosc.dstage\[4\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[4\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.iss.delayenb0 ringosc.iss.delayenb1/A ringosc.iss.ctrlen0/X VGND VGND VPWR
+ VPWR ringosc.ibufp00/A sky130_fd_sc_hd__einvn_4
XFILLER_15_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_390_ _349_/A _390_/D _337_/X VGND VGND VPWR VPWR _390_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_373_ _317_/X _373_/A1 _376_/S VGND VGND VPWR VPWR _373_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_287_ _279_/A _279_/B _385_/Q _384_/Q _284_/D VGND VGND VPWR VPWR _288_/B sky130_fd_sc_hd__o221a_1
X_356_ _306_/X input8/X _379_/S VGND VGND VPWR VPWR _356_/X sky130_fd_sc_hd__mux2_1
Xinput5 div[3] VGND VGND VPWR VPWR _189_/A sky130_fd_sc_hd__buf_1
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[3\].id.delayen1 ringosc.dstage\[3\].id.delayen1/A _371_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[3\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
X_210_ _385_/Q _400_/Q _208_/Y _209_/X VGND VGND VPWR VPWR _211_/A sky130_fd_sc_hd__a22o_1
XFILLER_18_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_339_ _348_/A VGND VGND VPWR VPWR _339_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.iss.delayenb1 ringosc.iss.delayenb1/A _379_/X VGND VGND VPWR VPWR ringosc.iss.delayen1/Z
+ sky130_fd_sc_hd__einvn_2
Xringosc.dstage\[0\].id.delaybuf0 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.dstage\[0\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
Xinput30 ext_trim[7] VGND VGND VPWR VPWR _362_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[3\].id.delayint0 ringosc.dstage\[3\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_32_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_372_ _297_/A _372_/A1 _379_/S VGND VGND VPWR VPWR _372_/X sky130_fd_sc_hd__mux2_2
XFILLER_24_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_286_ _284_/D _280_/A _285_/Y _288_/A VGND VGND VPWR VPWR _386_/D sky130_fd_sc_hd__a31o_1
XFILLER_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_355_ _315_/X _355_/A1 _379_/S VGND VGND VPWR VPWR _355_/X sky130_fd_sc_hd__mux2_1
Xinput6 div[4] VGND VGND VPWR VPWR _218_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_19_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xidiv16 idiv8/D idiv16/D irb/Y VGND VGND VPWR VPWR idiv16/Q idiv16/D sky130_fd_sc_hd__dfrbp_1
X_338_ _348_/A VGND VGND VPWR VPWR _338_/X sky130_fd_sc_hd__clkbuf_1
X_269_ _269_/A _269_/B VGND VGND VPWR VPWR _269_/X sky130_fd_sc_hd__or2_1
XFILLER_2_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[0\].id.delaybuf1 ringosc.dstage\[0\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[0\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xinput20 ext_trim[21] VGND VGND VPWR VPWR _361_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput31 ext_trim[8] VGND VGND VPWR VPWR _360_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.iss.delaybuf0 ringosc.iss.delayenb1/A VGND VGND VPWR VPWR ringosc.iss.delayen1/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_371_ _318_/X _371_/A1 _376_/S VGND VGND VPWR VPWR _371_/X sky130_fd_sc_hd__mux2_1
X_285_ _279_/A _279_/B _279_/C VGND VGND VPWR VPWR _285_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_354_ _307_/X input9/X _379_/S VGND VGND VPWR VPWR _354_/X sky130_fd_sc_hd__mux2_2
Xinput7 ext_trim[0] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_337_ _348_/A VGND VGND VPWR VPWR _337_/X sky130_fd_sc_hd__clkbuf_1
X_268_ _235_/Y _262_/X _267_/Y _393_/Q _235_/A VGND VGND VPWR VPWR _393_/D sky130_fd_sc_hd__a32o_1
X_199_ _401_/Q _284_/D _386_/Q _233_/B VGND VGND VPWR VPWR _401_/D sky130_fd_sc_hd__a22o_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput32 ext_trim[9] VGND VGND VPWR VPWR _358_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput10 ext_trim[12] VGND VGND VPWR VPWR _378_/A1 sky130_fd_sc_hd__buf_1
Xinput21 ext_trim[22] VGND VGND VPWR VPWR _359_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_370_ _291_/X _370_/A1 _376_/S VGND VGND VPWR VPWR _370_/X sky130_fd_sc_hd__mux2_1
X_284_ _387_/Q _284_/B _388_/Q _284_/D VGND VGND VPWR VPWR _288_/A sky130_fd_sc_hd__and4_1
Xringosc.dstage\[0\].id.delayen0 ringosc.dstage\[0\].id.delayen0/A _376_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XFILLER_14_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_353_ _352_/X _349_/A _353_/S VGND VGND VPWR VPWR _353_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 ext_trim[10] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_198_ _402_/Q _284_/D _387_/Q _233_/B VGND VGND VPWR VPWR _402_/D sky130_fd_sc_hd__a22o_1
X_267_ _267_/A _267_/B VGND VGND VPWR VPWR _267_/Y sky130_fd_sc_hd__nand2_1
X_336_ _348_/A VGND VGND VPWR VPWR _336_/X sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[7\].id.delayenb0 ringosc.dstage\[7\].id.delayenb1/A _362_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[7\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput22 ext_trim[23] VGND VGND VPWR VPWR _357_/A1 sky130_fd_sc_hd__buf_1
Xinput33 extclk_sel VGND VGND VPWR VPWR _196_/A sky130_fd_sc_hd__buf_1
XFILLER_16_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_319_ _306_/B _315_/C _310_/Y VGND VGND VPWR VPWR _319_/X sky130_fd_sc_hd__o21a_1
Xinput11 ext_trim[13] VGND VGND VPWR VPWR _377_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_32_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[0\].id.delayen1 ringosc.dstage\[0\].id.delayen1/A _377_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[0\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
Xinput9 ext_trim[11] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__buf_1
X_283_ _387_/Q _284_/B _388_/Q _281_/Y _284_/D VGND VGND VPWR VPWR _387_/D sky130_fd_sc_hd__o221a_1
X_352_ _351_/X idiv2/D _352_/S VGND VGND VPWR VPWR _352_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_266_ _309_/A _235_/Y _265_/X VGND VGND VPWR VPWR _394_/D sky130_fd_sc_hd__o21ai_1
Xringosc.dstage\[7\].id.delayenb1 ringosc.dstage\[7\].id.delayenb1/A _363_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[7\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
X_335_ _348_/A VGND VGND VPWR VPWR _335_/X sky130_fd_sc_hd__clkbuf_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_197_ _379_/S _197_/B VGND VGND VPWR VPWR _348_/A sky130_fd_sc_hd__nor2_8
XFILLER_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput34 osc VGND VGND VPWR VPWR _381_/D sky130_fd_sc_hd__clkbuf_1
X_318_ _380_/X _318_/B VGND VGND VPWR VPWR _318_/X sky130_fd_sc_hd__and2_1
X_249_ _290_/A VGND VGND VPWR VPWR _249_/Y sky130_fd_sc_hd__inv_2
Xinput12 ext_trim[14] VGND VGND VPWR VPWR _375_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput23 ext_trim[24] VGND VGND VPWR VPWR _355_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[8\].id.delayen0 ringosc.dstage\[8\].id.delayen0/A _360_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[8\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_282_ _176_/Y _281_/Y _233_/B VGND VGND VPWR VPWR _388_/D sky130_fd_sc_hd__a21oi_1
X_351_ _350_/X idiv4/D _351_/S VGND VGND VPWR VPWR _351_/X sky130_fd_sc_hd__mux2_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_403_ _349_/A _403_/D _348_/X VGND VGND VPWR VPWR _403_/Q sky130_fd_sc_hd__dfrtp_1
X_334_ _348_/A VGND VGND VPWR VPWR _334_/X sky130_fd_sc_hd__clkbuf_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_265_ _253_/Y _264_/A _253_/A _264_/Y _235_/A VGND VGND VPWR VPWR _265_/X sky130_fd_sc_hd__a221o_1
XFILLER_2_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_196_ _196_/A irb/A VGND VGND VPWR VPWR _197_/B sky130_fd_sc_hd__or2_4
XFILLER_23_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput24 ext_trim[25] VGND VGND VPWR VPWR _379_/A1 sky130_fd_sc_hd__buf_1
Xinput13 ext_trim[15] VGND VGND VPWR VPWR _373_/A1 sky130_fd_sc_hd__clkbuf_1
X_179_ _385_/Q VGND VGND VPWR VPWR _279_/A sky130_fd_sc_hd__inv_2
X_248_ _392_/Q _391_/Q VGND VGND VPWR VPWR _290_/A sky130_fd_sc_hd__or2_2
X_317_ _290_/A _315_/C _310_/Y VGND VGND VPWR VPWR _317_/X sky130_fd_sc_hd__o21a_1
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput35 reset VGND VGND VPWR VPWR irb/A sky130_fd_sc_hd__buf_1
XFILLER_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[7\].id.delaybuf0 ringosc.dstage\[6\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[3\].id.delayenb0 ringosc.dstage\[3\].id.delayenb1/A _370_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[3\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
XFILLER_22_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[11\].id.delayint0 ringosc.dstage\[11\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_7_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[8\].id.delayen1 ringosc.dstage\[8\].id.delayen1/A _361_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[8\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_281_ _387_/Q _284_/B VGND VGND VPWR VPWR _281_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_350_ idiv16/D idiv8/D _350_/S VGND VGND VPWR VPWR _350_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_195_ _403_/Q _284_/D _388_/Q _233_/B VGND VGND VPWR VPWR _403_/D sky130_fd_sc_hd__a22o_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_402_ _349_/A _402_/D _348_/A VGND VGND VPWR VPWR _402_/Q sky130_fd_sc_hd__dfrtp_1
X_264_ _264_/A VGND VGND VPWR VPWR _264_/Y sky130_fd_sc_hd__inv_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_333_ _348_/A VGND VGND VPWR VPWR _333_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput14 ext_trim[16] VGND VGND VPWR VPWR _371_/A1 sky130_fd_sc_hd__buf_1
X_247_ _247_/A VGND VGND VPWR VPWR _247_/Y sky130_fd_sc_hd__inv_2
X_316_ _309_/A _393_/Q _313_/A _290_/A _315_/X VGND VGND VPWR VPWR _316_/X sky130_fd_sc_hd__o41a_1
XFILLER_14_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput36 sel[0] VGND VGND VPWR VPWR _324_/C sky130_fd_sc_hd__clkbuf_2
Xinput25 ext_trim[2] VGND VGND VPWR VPWR _372_/A1 sky130_fd_sc_hd__clkbuf_1
X_178_ _386_/Q VGND VGND VPWR VPWR _279_/C sky130_fd_sc_hd__inv_2
XFILLER_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[7\].id.delaybuf1 ringosc.dstage\[7\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[7\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[3\].id.delayenb1 ringosc.dstage\[3\].id.delayenb1/A _371_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[3\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_280_ _280_/A VGND VGND VPWR VPWR _284_/B sky130_fd_sc_hd__inv_2
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_263_ _311_/C _239_/A _262_/X VGND VGND VPWR VPWR _264_/A sky130_fd_sc_hd__o21ai_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_194_ _284_/D VGND VGND VPWR VPWR _233_/B sky130_fd_sc_hd__clkinv_4
XFILLER_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_401_ _349_/A _401_/D _326_/X VGND VGND VPWR VPWR _401_/Q sky130_fd_sc_hd__dfrtp_1
X_332_ _348_/A VGND VGND VPWR VPWR _332_/X sky130_fd_sc_hd__clkbuf_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput37 sel[1] VGND VGND VPWR VPWR _323_/B sky130_fd_sc_hd__clkbuf_2
X_177_ _403_/Q VGND VGND VPWR VPWR _177_/Y sky130_fd_sc_hd__inv_2
X_246_ _294_/A _239_/Y _392_/Q _239_/A VGND VGND VPWR VPWR _247_/A sky130_fd_sc_hd__o22a_1
X_315_ _395_/Q _315_/B _315_/C VGND VGND VPWR VPWR _315_/X sky130_fd_sc_hd__and3_1
Xinput15 ext_trim[17] VGND VGND VPWR VPWR _369_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput26 ext_trim[3] VGND VGND VPWR VPWR _370_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_229_ _229_/A _229_/B VGND VGND VPWR VPWR _230_/A sky130_fd_sc_hd__nand2_1
Xringosc.dstage\[3\].id.delaybuf0 ringosc.dstage\[2\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[6\].id.delayint0 ringosc.dstage\[6\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.ibufp10 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.ibufp11/A sky130_fd_sc_hd__inv_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_331_ _348_/A VGND VGND VPWR VPWR _331_/X sky130_fd_sc_hd__clkbuf_1
X_193_ _383_/D _383_/Q _383_/D _383_/Q VGND VGND VPWR VPWR _284_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_262_ _267_/A _267_/B VGND VGND VPWR VPWR _262_/X sky130_fd_sc_hd__or2_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_400_ _349_/A _400_/D _327_/X VGND VGND VPWR VPWR _400_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput16 ext_trim[18] VGND VGND VPWR VPWR _367_/A1 sky130_fd_sc_hd__buf_1
X_176_ _388_/Q VGND VGND VPWR VPWR _176_/Y sky130_fd_sc_hd__inv_2
X_245_ _274_/B VGND VGND VPWR VPWR _269_/B sky130_fd_sc_hd__inv_2
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_314_ _392_/Q _315_/B _395_/Q VGND VGND VPWR VPWR _314_/X sky130_fd_sc_hd__o21a_1
Xinput27 ext_trim[4] VGND VGND VPWR VPWR _368_/A1 sky130_fd_sc_hd__buf_1
Xinput38 sel[2] VGND VGND VPWR VPWR _325_/A sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[5\].id.delayen0 ringosc.dstage\[5\].id.delayen0/A _366_/X VGND VGND
+ VPWR VPWR ringosc.ibufp10/A sky130_fd_sc_hd__einvp_2
XFILLER_9_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_228_ _208_/Y _209_/X _208_/Y _209_/X VGND VGND VPWR VPWR _229_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_10_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.dstage\[3\].id.delaybuf1 ringosc.dstage\[3\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[3\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_3_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.ibufp00 ringosc.ibufp00/A VGND VGND VPWR VPWR ringosc.ibufp01/A sky130_fd_sc_hd__clkinv_2
Xidiv2 idiv2/CLK idiv2/D irb/Y VGND VGND VPWR VPWR idiv2/Q idiv2/D sky130_fd_sc_hd__dfrbp_2
Xringosc.ibufp11 ringosc.ibufp11/A VGND VGND VPWR VPWR idiv2/CLK sky130_fd_sc_hd__inv_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ _348_/A VGND VGND VPWR VPWR _330_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ _313_/A _235_/Y _260_/X VGND VGND VPWR VPWR _395_/D sky130_fd_sc_hd__o21ai_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_192_ _324_/C VGND VGND VPWR VPWR _325_/C sky130_fd_sc_hd__inv_2
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_244_ _294_/B _239_/A _391_/Q _239_/Y VGND VGND VPWR VPWR _274_/B sky130_fd_sc_hd__o22a_1
X_313_ _313_/A _313_/B VGND VGND VPWR VPWR _318_/B sky130_fd_sc_hd__nand2_1
Xinput28 ext_trim[5] VGND VGND VPWR VPWR _366_/A1 sky130_fd_sc_hd__buf_1
Xinput17 ext_trim[19] VGND VGND VPWR VPWR _365_/A1 sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[5\].id.delayen1 ringosc.dstage\[5\].id.delayen1/A _367_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[5\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_22_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_227_ _279_/B _208_/B _208_/Y VGND VGND VPWR VPWR _227_/X sky130_fd_sc_hd__a21o_1
XFILLER_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[2\].id.delayint0 ringosc.dstage\[2\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xringosc.ibufp01 ringosc.ibufp01/A VGND VGND VPWR VPWR _349_/A sky130_fd_sc_hd__clkinv_8
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ _257_/Y _259_/A _257_/A _259_/Y _235_/A VGND VGND VPWR VPWR _260_/X sky130_fd_sc_hd__a221o_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_389_ _349_/A _389_/D _338_/X VGND VGND VPWR VPWR _389_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_191_ _323_/B VGND VGND VPWR VPWR _325_/B sky130_fd_sc_hd__inv_2
XFILLER_11_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 ext_trim[1] VGND VGND VPWR VPWR _374_/A1 sky130_fd_sc_hd__buf_1
X_243_ _274_/A VGND VGND VPWR VPWR _269_/A sky130_fd_sc_hd__inv_2
Xinput29 ext_trim[6] VGND VGND VPWR VPWR _364_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_312_ _392_/Q _315_/C _310_/Y VGND VGND VPWR VPWR _312_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_226_ _237_/A _237_/B _190_/A _225_/A _237_/C VGND VGND VPWR VPWR _226_/Y sky130_fd_sc_hd__a221oi_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[11\].id.delayenb0 ringosc.dstage\[11\].id.delayenb1/A _354_/X VGND
+ VGND VPWR VPWR ringosc.iss.delayenb1/A sky130_fd_sc_hd__einvn_4
XFILLER_17_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_209_ _385_/Q _400_/Q _385_/Q _400_/Q VGND VGND VPWR VPWR _209_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xidiv4 idiv2/D idiv4/D irb/Y VGND VGND VPWR VPWR idiv4/Q idiv4/D sky130_fd_sc_hd__dfrbp_2
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_190_ _190_/A VGND VGND VPWR VPWR _237_/A sky130_fd_sc_hd__inv_2
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_388_ _349_/A _388_/D _339_/X VGND VGND VPWR VPWR _388_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput19 ext_trim[20] VGND VGND VPWR VPWR _363_/A1 sky130_fd_sc_hd__clkbuf_1
X_242_ _187_/Y _239_/A _241_/Y VGND VGND VPWR VPWR _274_/A sky130_fd_sc_hd__o21ai_1
X_311_ _313_/A _394_/Q _311_/C VGND VGND VPWR VPWR _315_/C sky130_fd_sc_hd__or3_4
XFILLER_14_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_225_ _225_/A VGND VGND VPWR VPWR _237_/B sky130_fd_sc_hd__inv_2
Xringosc.dstage\[11\].id.delayenb1 ringosc.dstage\[11\].id.delayenb1/A _355_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[11\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
XFILLER_6_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_208_ _279_/B _208_/B VGND VGND VPWR VPWR _208_/Y sky130_fd_sc_hd__nor2_2
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_387_ _349_/A _387_/D _340_/X VGND VGND VPWR VPWR _387_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_310_ _313_/A _310_/B VGND VGND VPWR VPWR _310_/Y sky130_fd_sc_hd__nor2_2
X_241_ _389_/Q _276_/B VGND VGND VPWR VPWR _241_/Y sky130_fd_sc_hd__nand2_1
Xringosc.dstage\[2\].id.delayen0 ringosc.dstage\[2\].id.delayen0/A _372_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen0/Z sky130_fd_sc_hd__einvp_1
Xringosc.iss.const1 VGND VGND VPWR VPWR ringosc.iss.const1/HI ringosc.iss.const1/LO
+ sky130_fd_sc_hd__conb_1
X_224_ _211_/A _223_/Y _211_/A _223_/Y VGND VGND VPWR VPWR _225_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_207_ _386_/Q _401_/Q VGND VGND VPWR VPWR _207_/Y sky130_fd_sc_hd__nor2_1
Xringosc.dstage\[6\].id.delayenb0 ringosc.dstage\[6\].id.delayenb1/A _364_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[6\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
Xringosc.dstage\[11\].id.delaybuf0 ringosc.dstage\[10\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_386_ _349_/A _386_/D _341_/X VGND VGND VPWR VPWR _386_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_240_ _187_/Y _239_/A _390_/Q _239_/Y VGND VGND VPWR VPWR _276_/B sky130_fd_sc_hd__o22a_1
XFILLER_22_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[2\].id.delayen1 ringosc.dstage\[2\].id.delayen1/A _373_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[2\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_20_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_369_ _319_/X _369_/A1 _379_/S VGND VGND VPWR VPWR _369_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_223_ _386_/Q _401_/Q _207_/Y VGND VGND VPWR VPWR _223_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_206_ _387_/Q _402_/Q VGND VGND VPWR VPWR _206_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xringosc.dstage\[6\].id.delayenb1 ringosc.dstage\[6\].id.delayenb1/A _365_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[6\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
XFILLER_2_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[11\].id.delaybuf1 ringosc.dstage\[11\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[11\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_28_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_385_ _349_/A _385_/D _342_/X VGND VGND VPWR VPWR _385_/Q sky130_fd_sc_hd__dfrtp_2
Xringosc.iss.delayen0 ringosc.iss.delayen0/A _378_/X VGND VGND VPWR VPWR ringosc.ibufp00/A
+ sky130_fd_sc_hd__einvp_4
XFILLER_31_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_299_ _299_/A VGND VGND VPWR VPWR _299_/Y sky130_fd_sc_hd__inv_2
X_368_ _302_/Y _368_/A1 _379_/S VGND VGND VPWR VPWR _368_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_222_ _221_/A _221_/B _221_/X VGND VGND VPWR VPWR _237_/C sky130_fd_sc_hd__a21bo_1
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_205_ _388_/Q _403_/Q _176_/Y _177_/Y VGND VGND VPWR VPWR _214_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xringosc.dstage\[6\].id.delaybuf0 ringosc.ibufp10/A VGND VGND VPWR VPWR ringosc.dstage\[6\].id.delayenb1/A
+ sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[2\].id.delayenb0 ringosc.dstage\[2\].id.delayenb1/A _372_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[2\].id.delayen0/Z sky130_fd_sc_hd__einvn_2
Xringosc.dstage\[10\].id.delayint0 ringosc.dstage\[10\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[10\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
Xidiv8 idiv4/D idiv8/D irb/Y VGND VGND VPWR VPWR idiv8/Q idiv8/D sky130_fd_sc_hd__dfrbp_2
Xringosc.dstage\[9\].id.delayint0 ringosc.dstage\[9\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[9\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_25_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_384_ _349_/A _384_/D _343_/X VGND VGND VPWR VPWR _384_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xringosc.iss.delayen1 ringosc.iss.delayen1/A _379_/X VGND VGND VPWR VPWR ringosc.iss.delayen1/Z
+ sky130_fd_sc_hd__einvp_1
XFILLER_31_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_298_ _394_/Q _311_/C _313_/A _297_/Y VGND VGND VPWR VPWR _299_/A sky130_fd_sc_hd__a31o_1
X_367_ _310_/Y _367_/A1 _379_/S VGND VGND VPWR VPWR _367_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_221_ _221_/A _221_/B VGND VGND VPWR VPWR _221_/X sky130_fd_sc_hd__or2_1
XFILLER_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_204_ _396_/Q _233_/B VGND VGND VPWR VPWR _396_/D sky130_fd_sc_hd__or2_1
XFILLER_3_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xringosc.dstage\[6\].id.delaybuf1 ringosc.dstage\[6\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[6\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[2\].id.delayenb1 ringosc.dstage\[2\].id.delayenb1/A _373_/X VGND
+ VGND VPWR VPWR ringosc.dstage\[2\].id.delayen1/Z sky130_fd_sc_hd__einvn_2
XFILLER_29_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_383_ _349_/A _383_/D _344_/X VGND VGND VPWR VPWR _383_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_366_ _304_/X _366_/A1 _379_/S VGND VGND VPWR VPWR _366_/X sky130_fd_sc_hd__mux2_2
X_297_ _297_/A VGND VGND VPWR VPWR _297_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_220_ _212_/X _219_/X _212_/X _219_/X VGND VGND VPWR VPWR _221_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_349_ _349_/A VGND VGND VPWR VPWR _349_/X sky130_fd_sc_hd__clkbuf_1
X_203_ _397_/Q _284_/D _396_/Q _233_/B VGND VGND VPWR VPWR _397_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.iss.ctrlen0 _197_/B _378_/X VGND VGND VPWR VPWR ringosc.iss.ctrlen0/X sky130_fd_sc_hd__or2_2
XFILLER_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[2\].id.delaybuf0 ringosc.dstage\[1\].id.delayen0/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayenb1/A sky130_fd_sc_hd__clkbuf_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_382_ _349_/A _382_/D _345_/X VGND VGND VPWR VPWR _383_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[5\].id.delayint0 ringosc.dstage\[5\].id.delayen1/Z VGND VGND VPWR
+ VPWR ringosc.dstage\[5\].id.delayen0/A sky130_fd_sc_hd__clkinv_1
XFILLER_31_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_365_ _318_/B _365_/A1 _376_/S VGND VGND VPWR VPWR _365_/X sky130_fd_sc_hd__mux2_2
X_296_ _395_/Q _394_/Q VGND VGND VPWR VPWR _297_/A sky130_fd_sc_hd__or2_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_348_ _348_/A VGND VGND VPWR VPWR _348_/X sky130_fd_sc_hd__clkbuf_1
X_279_ _279_/A _279_/B _279_/C VGND VGND VPWR VPWR _280_/A sky130_fd_sc_hd__or3_1
XFILLER_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_202_ _397_/Q _233_/B _398_/Q _284_/D VGND VGND VPWR VPWR _398_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[7\].id.delayen0 ringosc.dstage\[7\].id.delayen0/A _362_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[7\].id.delayen0/Z sky130_fd_sc_hd__einvp_2
XFILLER_18_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[2\].id.delaybuf1 ringosc.dstage\[2\].id.delayenb1/A VGND VGND VPWR
+ VPWR ringosc.dstage\[2\].id.delayen1/A sky130_fd_sc_hd__clkbuf_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_381_ _349_/A _381_/D _346_/X VGND VGND VPWR VPWR _382_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_25_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput40 idiv2/D VGND VGND VPWR VPWR clockd[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_364_ _293_/X _364_/A1 _379_/S VGND VGND VPWR VPWR _364_/X sky130_fd_sc_hd__mux2_1
X_295_ _309_/C VGND VGND VPWR VPWR _306_/B sky130_fd_sc_hd__inv_2
XFILLER_9_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_278_ _389_/Q _235_/Y _188_/Y _235_/A VGND VGND VPWR VPWR _389_/D sky130_fd_sc_hd__o22a_1
X_347_ _395_/Q VGND VGND VPWR VPWR _347_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_201_ _399_/Q _284_/D _384_/Q _233_/B VGND VGND VPWR VPWR _399_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xringosc.dstage\[11\].id.delayen0 ringosc.dstage\[11\].id.delayen0/A _354_/X VGND
+ VGND VPWR VPWR ringosc.iss.delayenb1/A sky130_fd_sc_hd__einvp_4
XFILLER_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[7\].id.delayen1 ringosc.dstage\[7\].id.delayen1/A _363_/X VGND VGND
+ VPWR VPWR ringosc.dstage\[7\].id.delayen1/Z sky130_fd_sc_hd__einvp_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_380_ _313_/B _292_/B _395_/Q VGND VGND VPWR VPWR _380_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput41 idiv4/D VGND VGND VPWR VPWR clockd[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_31_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

