VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_pll
  CLASS BLOCK ;
  FOREIGN digital_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.135 BY 100.855 ;
  PIN clockp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END clockp[0]
  PIN clockp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 96.855 34.870 100.855 ;
    END
  END clockp[1]
  PIN dco
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 96.855 50.970 100.855 ;
    END
  END dco
  PIN div[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 96.855 69.370 100.855 ;
    END
  END div[0]
  PIN div[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 86.135 17.040 90.135 17.640 ;
    END
  END div[1]
  PIN div[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END div[2]
  PIN div[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END div[3]
  PIN div[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END div[4]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 96.855 85.470 100.855 ;
    END
  END enable
  PIN ext_trim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 96.855 44.070 100.855 ;
    END
  END ext_trim[0]
  PIN ext_trim[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END ext_trim[10]
  PIN ext_trim[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END ext_trim[11]
  PIN ext_trim[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 96.855 18.770 100.855 ;
    END
  END ext_trim[12]
  PIN ext_trim[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 96.855 27.970 100.855 ;
    END
  END ext_trim[13]
  PIN ext_trim[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END ext_trim[14]
  PIN ext_trim[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END ext_trim[15]
  PIN ext_trim[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 86.135 54.440 90.135 55.040 ;
    END
  END ext_trim[16]
  PIN ext_trim[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END ext_trim[17]
  PIN ext_trim[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 86.135 6.840 90.135 7.440 ;
    END
  END ext_trim[18]
  PIN ext_trim[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 96.855 76.270 100.855 ;
    END
  END ext_trim[19]
  PIN ext_trim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END ext_trim[1]
  PIN ext_trim[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END ext_trim[20]
  PIN ext_trim[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END ext_trim[21]
  PIN ext_trim[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 86.135 78.240 90.135 78.840 ;
    END
  END ext_trim[22]
  PIN ext_trim[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 96.855 11.870 100.855 ;
    END
  END ext_trim[23]
  PIN ext_trim[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 96.855 2.670 100.855 ;
    END
  END ext_trim[24]
  PIN ext_trim[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END ext_trim[25]
  PIN ext_trim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END ext_trim[2]
  PIN ext_trim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 96.855 60.170 100.855 ;
    END
  END ext_trim[3]
  PIN ext_trim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END ext_trim[4]
  PIN ext_trim[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END ext_trim[5]
  PIN ext_trim[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END ext_trim[6]
  PIN ext_trim[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 86.135 68.040 90.135 68.640 ;
    END
  END ext_trim[7]
  PIN ext_trim[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 86.135 30.640 90.135 31.240 ;
    END
  END ext_trim[8]
  PIN ext_trim[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 86.135 91.840 90.135 92.440 ;
    END
  END ext_trim[9]
  PIN osc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 86.135 40.840 90.135 41.440 ;
    END
  END osc
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END resetb
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 70.270 10.640 71.870 90.000 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 44.050 10.640 45.650 90.000 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 17.830 10.640 19.430 90.000 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 75.575 84.180 77.175 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 49.280 84.180 50.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 22.985 84.180 24.585 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 57.160 10.640 58.760 90.000 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.640 32.540 90.000 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 62.425 84.180 64.025 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 36.135 84.180 37.735 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 84.180 89.845 ;
      LAYER met1 ;
        RECT 2.370 10.240 85.490 90.000 ;
      LAYER met2 ;
        RECT 2.950 96.575 11.310 96.855 ;
        RECT 12.150 96.575 18.210 96.855 ;
        RECT 19.050 96.575 27.410 96.855 ;
        RECT 28.250 96.575 34.310 96.855 ;
        RECT 35.150 96.575 43.510 96.855 ;
        RECT 44.350 96.575 50.410 96.855 ;
        RECT 51.250 96.575 59.610 96.855 ;
        RECT 60.450 96.575 68.810 96.855 ;
        RECT 69.650 96.575 75.710 96.855 ;
        RECT 76.550 96.575 84.910 96.855 ;
        RECT 2.400 4.280 85.460 96.575 ;
        RECT 2.950 4.000 9.010 4.280 ;
        RECT 9.850 4.000 18.210 4.280 ;
        RECT 19.050 4.000 25.110 4.280 ;
        RECT 25.950 4.000 34.310 4.280 ;
        RECT 35.150 4.000 41.210 4.280 ;
        RECT 42.050 4.000 50.410 4.280 ;
        RECT 51.250 4.000 57.310 4.280 ;
        RECT 58.150 4.000 66.510 4.280 ;
        RECT 67.350 4.000 75.710 4.280 ;
        RECT 76.550 4.000 82.610 4.280 ;
        RECT 83.450 4.000 85.460 4.280 ;
      LAYER met3 ;
        RECT 4.000 91.440 85.735 92.305 ;
        RECT 4.000 86.040 86.135 91.440 ;
        RECT 4.400 84.640 86.135 86.040 ;
        RECT 4.000 79.240 86.135 84.640 ;
        RECT 4.000 77.840 85.735 79.240 ;
        RECT 4.000 75.840 86.135 77.840 ;
        RECT 4.400 74.440 86.135 75.840 ;
        RECT 4.000 69.040 86.135 74.440 ;
        RECT 4.000 67.640 85.735 69.040 ;
        RECT 4.000 62.240 86.135 67.640 ;
        RECT 4.400 60.840 86.135 62.240 ;
        RECT 4.000 55.440 86.135 60.840 ;
        RECT 4.000 54.040 85.735 55.440 ;
        RECT 4.000 52.040 86.135 54.040 ;
        RECT 4.400 50.640 86.135 52.040 ;
        RECT 4.000 41.840 86.135 50.640 ;
        RECT 4.000 40.440 85.735 41.840 ;
        RECT 4.000 38.440 86.135 40.440 ;
        RECT 4.400 37.040 86.135 38.440 ;
        RECT 4.000 31.640 86.135 37.040 ;
        RECT 4.000 30.240 85.735 31.640 ;
        RECT 4.000 28.240 86.135 30.240 ;
        RECT 4.400 26.840 86.135 28.240 ;
        RECT 4.000 18.040 86.135 26.840 ;
        RECT 4.000 16.640 85.735 18.040 ;
        RECT 4.000 14.640 86.135 16.640 ;
        RECT 4.400 13.240 86.135 14.640 ;
        RECT 4.000 7.840 86.135 13.240 ;
        RECT 4.000 6.975 85.735 7.840 ;
      LAYER met5 ;
        RECT 5.520 65.625 84.180 73.975 ;
        RECT 5.520 52.480 84.180 60.825 ;
        RECT 5.520 39.335 84.180 47.680 ;
  END
END digital_pll
END LIBRARY

