VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_pll
  CLASS BLOCK ;
  FOREIGN digital_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 114.895 BY 125.615 ;
  PIN clockc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END clockc
  PIN clockd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END clockd[0]
  PIN clockd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END clockd[1]
  PIN clockd[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.895 102.040 114.895 102.640 ;
    END
  END clockd[2]
  PIN clockd[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END clockd[3]
  PIN clockp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END clockp[0]
  PIN clockp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END clockp[1]
  PIN dco
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END dco
  PIN div[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.895 78.240 114.895 78.840 ;
    END
  END div[0]
  PIN div[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 121.615 99.270 125.615 ;
    END
  END div[1]
  PIN div[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 121.615 39.470 125.615 ;
    END
  END div[2]
  PIN div[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END div[3]
  PIN div[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 121.615 73.970 125.615 ;
    END
  END div[4]
  PIN ext_trim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 121.615 83.170 125.615 ;
    END
  END ext_trim[0]
  PIN ext_trim[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END ext_trim[10]
  PIN ext_trim[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 121.615 14.170 125.615 ;
    END
  END ext_trim[11]
  PIN ext_trim[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.895 27.240 114.895 27.840 ;
    END
  END ext_trim[12]
  PIN ext_trim[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END ext_trim[13]
  PIN ext_trim[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END ext_trim[14]
  PIN ext_trim[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.895 88.440 114.895 89.040 ;
    END
  END ext_trim[15]
  PIN ext_trim[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 121.615 23.370 125.615 ;
    END
  END ext_trim[16]
  PIN ext_trim[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END ext_trim[17]
  PIN ext_trim[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 121.615 30.270 125.615 ;
    END
  END ext_trim[18]
  PIN ext_trim[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.895 51.040 114.895 51.640 ;
    END
  END ext_trim[19]
  PIN ext_trim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 121.615 64.770 125.615 ;
    END
  END ext_trim[1]
  PIN ext_trim[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 121.615 57.870 125.615 ;
    END
  END ext_trim[20]
  PIN ext_trim[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END ext_trim[21]
  PIN ext_trim[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END ext_trim[22]
  PIN ext_trim[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.895 115.640 114.895 116.240 ;
    END
  END ext_trim[23]
  PIN ext_trim[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END ext_trim[24]
  PIN ext_trim[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 121.615 48.670 125.615 ;
    END
  END ext_trim[25]
  PIN ext_trim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END ext_trim[2]
  PIN ext_trim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.895 40.840 114.895 41.440 ;
    END
  END ext_trim[3]
  PIN ext_trim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END ext_trim[4]
  PIN ext_trim[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.895 64.640 114.895 65.240 ;
    END
  END ext_trim[5]
  PIN ext_trim[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END ext_trim[6]
  PIN ext_trim[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 121.615 4.970 125.615 ;
    END
  END ext_trim[7]
  PIN ext_trim[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END ext_trim[8]
  PIN ext_trim[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.895 13.640 114.895 14.240 ;
    END
  END ext_trim[9]
  PIN extclk_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END extclk_sel
  PIN osc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 121.615 90.070 125.615 ;
    END
  END osc
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END reset
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END sel[0]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 121.615 108.470 125.615 ;
    END
  END sel[1]
  PIN sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END sel[2]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 90.970 10.640 92.570 114.480 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 56.470 10.640 58.070 114.480 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.970 10.640 23.570 114.480 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 95.975 109.020 97.575 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 61.520 109.020 63.120 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 27.065 109.020 28.665 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 73.720 10.640 75.320 114.480 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.220 10.640 40.820 114.480 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 78.745 109.020 80.345 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 44.295 109.020 45.895 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 109.020 114.325 ;
      LAYER met1 ;
        RECT 2.370 10.640 110.790 114.480 ;
      LAYER met2 ;
        RECT 2.400 121.335 4.410 121.615 ;
        RECT 5.250 121.335 13.610 121.615 ;
        RECT 14.450 121.335 22.810 121.615 ;
        RECT 23.650 121.335 29.710 121.615 ;
        RECT 30.550 121.335 38.910 121.615 ;
        RECT 39.750 121.335 48.110 121.615 ;
        RECT 48.950 121.335 57.310 121.615 ;
        RECT 58.150 121.335 64.210 121.615 ;
        RECT 65.050 121.335 73.410 121.615 ;
        RECT 74.250 121.335 82.610 121.615 ;
        RECT 83.450 121.335 89.510 121.615 ;
        RECT 90.350 121.335 98.710 121.615 ;
        RECT 99.550 121.335 107.910 121.615 ;
        RECT 108.750 121.335 110.760 121.615 ;
        RECT 2.400 4.280 110.760 121.335 ;
        RECT 2.950 4.000 9.010 4.280 ;
        RECT 9.850 4.000 18.210 4.280 ;
        RECT 19.050 4.000 27.410 4.280 ;
        RECT 28.250 4.000 34.310 4.280 ;
        RECT 35.150 4.000 43.510 4.280 ;
        RECT 44.350 4.000 52.710 4.280 ;
        RECT 53.550 4.000 59.610 4.280 ;
        RECT 60.450 4.000 68.810 4.280 ;
        RECT 69.650 4.000 78.010 4.280 ;
        RECT 78.850 4.000 84.910 4.280 ;
        RECT 85.750 4.000 94.110 4.280 ;
        RECT 94.950 4.000 103.310 4.280 ;
        RECT 104.150 4.000 110.210 4.280 ;
      LAYER met3 ;
        RECT 4.400 115.240 110.495 116.105 ;
        RECT 4.000 103.040 110.895 115.240 ;
        RECT 4.400 101.640 110.495 103.040 ;
        RECT 4.000 89.440 110.895 101.640 ;
        RECT 4.400 88.040 110.495 89.440 ;
        RECT 4.000 79.240 110.895 88.040 ;
        RECT 4.400 77.840 110.495 79.240 ;
        RECT 4.000 65.640 110.895 77.840 ;
        RECT 4.400 64.240 110.495 65.640 ;
        RECT 4.000 52.040 110.895 64.240 ;
        RECT 4.400 50.640 110.495 52.040 ;
        RECT 4.000 41.840 110.895 50.640 ;
        RECT 4.400 40.440 110.495 41.840 ;
        RECT 4.000 28.240 110.895 40.440 ;
        RECT 4.400 26.840 110.495 28.240 ;
        RECT 4.000 14.640 110.895 26.840 ;
        RECT 4.400 13.240 110.495 14.640 ;
        RECT 4.000 10.715 110.895 13.240 ;
      LAYER met5 ;
        RECT 5.520 81.945 109.020 94.375 ;
        RECT 5.520 64.720 109.020 77.145 ;
        RECT 5.520 47.495 109.020 59.920 ;
  END
END digital_pll
END LIBRARY

