magic
tech sky130A
magscale 1 2
timestamp 1619516433
<< locali >>
rect 14565 17527 14599 17629
rect 5181 13855 5215 13957
rect 10517 13855 10551 13957
rect 4353 12631 4387 12937
rect 9321 9435 9355 9673
rect 8953 7735 8987 7905
rect 6561 2295 6595 2465
<< viali >>
rect 1501 17833 1535 17867
rect 2145 17833 2179 17867
rect 1593 17765 1627 17799
rect 15025 17765 15059 17799
rect 16497 17765 16531 17799
rect 2329 17697 2363 17731
rect 3157 17697 3191 17731
rect 4629 17697 4663 17731
rect 5457 17697 5491 17731
rect 5641 17697 5675 17731
rect 7021 17697 7055 17731
rect 7665 17697 7699 17731
rect 8493 17697 8527 17731
rect 9597 17697 9631 17731
rect 9781 17697 9815 17731
rect 10517 17697 10551 17731
rect 11161 17697 11195 17731
rect 12357 17697 12391 17731
rect 13001 17697 13035 17731
rect 13829 17697 13863 17731
rect 14749 17697 14783 17731
rect 14841 17697 14875 17731
rect 15669 17697 15703 17731
rect 14565 17629 14599 17663
rect 3341 17561 3375 17595
rect 7205 17561 7239 17595
rect 10701 17561 10735 17595
rect 16313 17561 16347 17595
rect 4813 17493 4847 17527
rect 5273 17493 5307 17527
rect 7849 17493 7883 17527
rect 8401 17493 8435 17527
rect 9689 17493 9723 17527
rect 11345 17493 11379 17527
rect 12541 17493 12575 17527
rect 13185 17493 13219 17527
rect 14013 17493 14047 17527
rect 14565 17493 14599 17527
rect 15025 17493 15059 17527
rect 15761 17493 15795 17527
rect 14638 17289 14672 17323
rect 2881 17221 2915 17255
rect 5181 17221 5215 17255
rect 3709 17153 3743 17187
rect 8033 17153 8067 17187
rect 13645 17153 13679 17187
rect 1777 17085 1811 17119
rect 2605 17085 2639 17119
rect 2743 17085 2777 17119
rect 2973 17085 3007 17119
rect 3433 17085 3467 17119
rect 5825 17085 5859 17119
rect 7297 17085 7331 17119
rect 9781 17085 9815 17119
rect 10425 17085 10459 17119
rect 10517 17085 10551 17119
rect 10793 17085 10827 17119
rect 13921 17085 13955 17119
rect 14381 17085 14415 17119
rect 2421 17017 2455 17051
rect 9505 17017 9539 17051
rect 10609 17017 10643 17051
rect 1961 16949 1995 16983
rect 5641 16949 5675 16983
rect 7481 16949 7515 16983
rect 10241 16949 10275 16983
rect 12173 16949 12207 16983
rect 16129 16949 16163 16983
rect 5825 16745 5859 16779
rect 9781 16745 9815 16779
rect 12173 16745 12207 16779
rect 12817 16745 12851 16779
rect 1685 16677 1719 16711
rect 4721 16677 4755 16711
rect 5457 16677 5491 16711
rect 6561 16677 6595 16711
rect 11161 16677 11195 16711
rect 4629 16609 4663 16643
rect 5273 16609 5307 16643
rect 5549 16609 5583 16643
rect 5641 16609 5675 16643
rect 11069 16609 11103 16643
rect 11253 16609 11287 16643
rect 11437 16609 11471 16643
rect 12081 16609 12115 16643
rect 12725 16609 12759 16643
rect 12909 16609 12943 16643
rect 13369 16609 13403 16643
rect 1409 16541 1443 16575
rect 6285 16541 6319 16575
rect 9965 16541 9999 16575
rect 10057 16541 10091 16575
rect 10425 16541 10459 16575
rect 14749 16541 14783 16575
rect 15025 16541 15059 16575
rect 10885 16473 10919 16507
rect 3157 16405 3191 16439
rect 8033 16405 8067 16439
rect 13553 16405 13587 16439
rect 16497 16405 16531 16439
rect 2881 16201 2915 16235
rect 11069 16201 11103 16235
rect 14197 16201 14231 16235
rect 3893 16065 3927 16099
rect 7481 16065 7515 16099
rect 8677 16065 8711 16099
rect 8861 16065 8895 16099
rect 10057 16065 10091 16099
rect 10149 16065 10183 16099
rect 16313 16065 16347 16099
rect 1501 15997 1535 16031
rect 2145 15997 2179 16031
rect 2973 15997 3007 16031
rect 6837 15997 6871 16031
rect 7021 15997 7055 16031
rect 7297 15997 7331 16031
rect 7665 15997 7699 16031
rect 8401 15997 8435 16031
rect 8493 15997 8527 16031
rect 9781 15997 9815 16031
rect 9965 15997 9999 16031
rect 10333 15997 10367 16031
rect 10977 15997 11011 16031
rect 11989 15997 12023 16031
rect 12449 15997 12483 16031
rect 15485 15997 15519 16031
rect 15669 15997 15703 16031
rect 16221 15997 16255 16031
rect 4169 15929 4203 15963
rect 8217 15929 8251 15963
rect 8769 15929 8803 15963
rect 12725 15929 12759 15963
rect 15117 15929 15151 15963
rect 1685 15861 1719 15895
rect 2329 15861 2363 15895
rect 5641 15861 5675 15895
rect 10517 15861 10551 15895
rect 11805 15861 11839 15895
rect 5825 15657 5859 15691
rect 10425 15657 10459 15691
rect 12725 15657 12759 15691
rect 16589 15657 16623 15691
rect 2789 15589 2823 15623
rect 6193 15589 6227 15623
rect 10057 15589 10091 15623
rect 10241 15589 10275 15623
rect 15117 15589 15151 15623
rect 1869 15521 1903 15555
rect 2697 15521 2731 15555
rect 2881 15521 2915 15555
rect 3019 15521 3053 15555
rect 4261 15521 4295 15555
rect 5365 15521 5399 15555
rect 6009 15521 6043 15555
rect 6105 15521 6139 15555
rect 6377 15521 6411 15555
rect 7021 15521 7055 15555
rect 7205 15521 7239 15555
rect 7573 15521 7607 15555
rect 7941 15521 7975 15555
rect 11161 15521 11195 15555
rect 11989 15521 12023 15555
rect 12173 15521 12207 15555
rect 12265 15521 12299 15555
rect 12357 15521 12391 15555
rect 12541 15521 12575 15555
rect 13829 15521 13863 15555
rect 3157 15453 3191 15487
rect 7757 15453 7791 15487
rect 8033 15453 8067 15487
rect 10885 15453 10919 15487
rect 14841 15453 14875 15487
rect 10977 15385 11011 15419
rect 13737 15385 13771 15419
rect 2053 15317 2087 15351
rect 2513 15317 2547 15351
rect 4353 15317 4387 15351
rect 5273 15317 5307 15351
rect 11069 15317 11103 15351
rect 4077 15113 4111 15147
rect 5825 15113 5859 15147
rect 10149 15113 10183 15147
rect 13093 15113 13127 15147
rect 1685 14977 1719 15011
rect 3157 14977 3191 15011
rect 4629 14977 4663 15011
rect 4813 14977 4847 15011
rect 7389 14977 7423 15011
rect 10793 14977 10827 15011
rect 12173 14977 12207 15011
rect 13645 14977 13679 15011
rect 14565 14977 14599 15011
rect 1409 14909 1443 14943
rect 3801 14909 3835 14943
rect 3893 14909 3927 14943
rect 4169 14909 4203 14943
rect 4905 14909 4939 14943
rect 5733 14909 5767 14943
rect 6929 14909 6963 14943
rect 8401 14909 8435 14943
rect 8585 14909 8619 14943
rect 8769 14909 8803 14943
rect 8953 14909 8987 14943
rect 9321 14909 9355 14943
rect 10330 14909 10364 14943
rect 10701 14909 10735 14943
rect 12081 14909 12115 14943
rect 12265 14909 12299 14943
rect 13001 14909 13035 14943
rect 13185 14909 13219 14943
rect 13829 14909 13863 14943
rect 14105 14909 14139 14943
rect 14749 14909 14783 14943
rect 14933 14909 14967 14943
rect 15025 14909 15059 14943
rect 15117 14909 15151 14943
rect 15301 14909 15335 14943
rect 15761 14909 15795 14943
rect 7941 14841 7975 14875
rect 3617 14773 3651 14807
rect 4629 14773 4663 14807
rect 10333 14773 10367 14807
rect 14013 14773 14047 14807
rect 15853 14773 15887 14807
rect 2513 14569 2547 14603
rect 2973 14569 3007 14603
rect 7757 14569 7791 14603
rect 8585 14569 8619 14603
rect 10149 14569 10183 14603
rect 12449 14569 12483 14603
rect 16405 14569 16439 14603
rect 3341 14501 3375 14535
rect 8401 14501 8435 14535
rect 10977 14501 11011 14535
rect 13277 14501 13311 14535
rect 15209 14501 15243 14535
rect 1685 14433 1719 14467
rect 2329 14433 2363 14467
rect 2513 14433 2547 14467
rect 3157 14433 3191 14467
rect 7389 14433 7423 14467
rect 8217 14433 8251 14467
rect 9965 14433 9999 14467
rect 10241 14433 10275 14467
rect 13093 14433 13127 14467
rect 13185 14433 13219 14467
rect 13461 14433 13495 14467
rect 13553 14433 13587 14467
rect 15117 14433 15151 14467
rect 15301 14433 15335 14467
rect 15485 14433 15519 14467
rect 15945 14433 15979 14467
rect 16037 14433 16071 14467
rect 16221 14433 16255 14467
rect 4537 14365 4571 14399
rect 4813 14365 4847 14399
rect 7481 14365 7515 14399
rect 10701 14365 10735 14399
rect 1869 14297 1903 14331
rect 6285 14229 6319 14263
rect 7389 14229 7423 14263
rect 9781 14229 9815 14263
rect 12909 14229 12943 14263
rect 14933 14229 14967 14263
rect 5273 14025 5307 14059
rect 6929 14025 6963 14059
rect 8125 14025 8159 14059
rect 9965 14025 9999 14059
rect 11161 14025 11195 14059
rect 14105 14025 14139 14059
rect 16405 14025 16439 14059
rect 2053 13957 2087 13991
rect 3801 13957 3835 13991
rect 5181 13957 5215 13991
rect 9413 13957 9447 13991
rect 10517 13957 10551 13991
rect 7113 13889 7147 13923
rect 8309 13889 8343 13923
rect 8401 13889 8435 13923
rect 8769 13889 8803 13923
rect 10057 13889 10091 13923
rect 12357 13889 12391 13923
rect 12633 13889 12667 13923
rect 14933 13889 14967 13923
rect 1869 13821 1903 13855
rect 2697 13821 2731 13855
rect 3525 13821 3559 13855
rect 3617 13821 3651 13855
rect 3893 13821 3927 13855
rect 4353 13821 4387 13855
rect 5181 13821 5215 13855
rect 5457 13821 5491 13855
rect 5917 13821 5951 13855
rect 6837 13821 6871 13855
rect 9594 13821 9628 13855
rect 10517 13821 10551 13855
rect 10609 13821 10643 13855
rect 10793 13821 10827 13855
rect 10977 13821 11011 13855
rect 14657 13821 14691 13855
rect 2881 13753 2915 13787
rect 4445 13753 4479 13787
rect 5549 13753 5583 13787
rect 5641 13753 5675 13787
rect 5779 13753 5813 13787
rect 10885 13753 10919 13787
rect 2513 13685 2547 13719
rect 3341 13685 3375 13719
rect 7113 13685 7147 13719
rect 9597 13685 9631 13719
rect 4261 13481 4295 13515
rect 7205 13481 7239 13515
rect 7941 13481 7975 13515
rect 10701 13481 10735 13515
rect 10885 13481 10919 13515
rect 12909 13481 12943 13515
rect 15025 13481 15059 13515
rect 16037 13481 16071 13515
rect 2973 13413 3007 13447
rect 3203 13413 3237 13447
rect 4445 13413 4479 13447
rect 5181 13413 5215 13447
rect 6193 13413 6227 13447
rect 12633 13413 12667 13447
rect 12817 13413 12851 13447
rect 13737 13413 13771 13447
rect 15209 13413 15243 13447
rect 1409 13345 1443 13379
rect 2053 13345 2087 13379
rect 2881 13345 2915 13379
rect 3065 13345 3099 13379
rect 4629 13345 4663 13379
rect 5089 13345 5123 13379
rect 5963 13345 5997 13379
rect 6101 13345 6135 13379
rect 6377 13345 6411 13379
rect 6837 13345 6871 13379
rect 7021 13345 7055 13379
rect 8217 13345 8251 13379
rect 9505 13345 9539 13379
rect 10882 13345 10916 13379
rect 11989 13345 12023 13379
rect 13001 13345 13035 13379
rect 13645 13345 13679 13379
rect 14749 13345 14783 13379
rect 14933 13345 14967 13379
rect 15301 13345 15335 13379
rect 15853 13345 15887 13379
rect 16129 13345 16163 13379
rect 3341 13277 3375 13311
rect 7941 13277 7975 13311
rect 8125 13277 8159 13311
rect 11345 13277 11379 13311
rect 1593 13209 1627 13243
rect 9597 13209 9631 13243
rect 2237 13141 2271 13175
rect 2697 13141 2731 13175
rect 5825 13141 5859 13175
rect 11253 13141 11287 13175
rect 11805 13141 11839 13175
rect 13185 13141 13219 13175
rect 3157 12937 3191 12971
rect 4353 12937 4387 12971
rect 4445 12937 4479 12971
rect 7849 12937 7883 12971
rect 11069 12937 11103 12971
rect 12081 12937 12115 12971
rect 12909 12937 12943 12971
rect 14657 12937 14691 12971
rect 16221 12937 16255 12971
rect 1409 12801 1443 12835
rect 1685 12801 1719 12835
rect 3709 12733 3743 12767
rect 3801 12733 3835 12767
rect 15209 12869 15243 12903
rect 4813 12801 4847 12835
rect 4905 12801 4939 12835
rect 8585 12801 8619 12835
rect 12725 12801 12759 12835
rect 4629 12733 4663 12767
rect 4721 12733 4755 12767
rect 5089 12733 5123 12767
rect 5917 12733 5951 12767
rect 7205 12733 7239 12767
rect 7353 12733 7387 12767
rect 7670 12733 7704 12767
rect 8309 12733 8343 12767
rect 10977 12733 11011 12767
rect 12081 12733 12115 12767
rect 12265 12733 12299 12767
rect 13001 12733 13035 12767
rect 13921 12733 13955 12767
rect 14565 12733 14599 12767
rect 15393 12733 15427 12767
rect 15577 12733 15611 12767
rect 15761 12733 15795 12767
rect 16405 12733 16439 12767
rect 7481 12665 7515 12699
rect 7573 12665 7607 12699
rect 13737 12665 13771 12699
rect 15485 12665 15519 12699
rect 4353 12597 4387 12631
rect 5825 12597 5859 12631
rect 10057 12597 10091 12631
rect 12725 12597 12759 12631
rect 14105 12597 14139 12631
rect 3341 12393 3375 12427
rect 7481 12393 7515 12427
rect 10701 12393 10735 12427
rect 16405 12393 16439 12427
rect 11805 12325 11839 12359
rect 15393 12325 15427 12359
rect 1869 12257 1903 12291
rect 2513 12257 2547 12291
rect 3157 12257 3191 12291
rect 3341 12257 3375 12291
rect 4537 12257 4571 12291
rect 5181 12257 5215 12291
rect 5917 12257 5951 12291
rect 6561 12257 6595 12291
rect 7021 12257 7055 12291
rect 7665 12257 7699 12291
rect 7757 12257 7791 12291
rect 8033 12257 8067 12291
rect 9505 12257 9539 12291
rect 10885 12257 10919 12291
rect 10977 12257 11011 12291
rect 11253 12257 11287 12291
rect 11989 12257 12023 12291
rect 12081 12257 12115 12291
rect 12817 12257 12851 12291
rect 12909 12257 12943 12291
rect 13093 12257 13127 12291
rect 13645 12257 13679 12291
rect 15301 12257 15335 12291
rect 15485 12257 15519 12291
rect 15669 12257 15703 12291
rect 16589 12257 16623 12291
rect 4261 12189 4295 12223
rect 4445 12189 4479 12223
rect 6745 12189 6779 12223
rect 6854 12189 6888 12223
rect 9597 12189 9631 12223
rect 11345 12189 11379 12223
rect 13001 12189 13035 12223
rect 6377 12121 6411 12155
rect 6653 12121 6687 12155
rect 11805 12121 11839 12155
rect 2053 12053 2087 12087
rect 2697 12053 2731 12087
rect 4353 12053 4387 12087
rect 5089 12053 5123 12087
rect 5825 12053 5859 12087
rect 7941 12053 7975 12087
rect 12633 12053 12667 12087
rect 13737 12053 13771 12087
rect 15117 12053 15151 12087
rect 5365 11849 5399 11883
rect 5825 11849 5859 11883
rect 12265 11849 12299 11883
rect 13093 11849 13127 11883
rect 13553 11849 13587 11883
rect 15393 11849 15427 11883
rect 12725 11781 12759 11815
rect 2605 11713 2639 11747
rect 13001 11713 13035 11747
rect 14013 11713 14047 11747
rect 3801 11645 3835 11679
rect 4261 11645 4295 11679
rect 4354 11645 4388 11679
rect 4629 11645 4663 11679
rect 4726 11645 4760 11679
rect 5549 11645 5583 11679
rect 5641 11645 5675 11679
rect 5917 11645 5951 11679
rect 6837 11645 6871 11679
rect 6985 11645 7019 11679
rect 7302 11645 7336 11679
rect 8493 11645 8527 11679
rect 10977 11645 11011 11679
rect 12081 11645 12115 11679
rect 13093 11645 13127 11679
rect 13737 11645 13771 11679
rect 13921 11645 13955 11679
rect 14105 11645 14139 11679
rect 14289 11645 14323 11679
rect 14933 11645 14967 11679
rect 15574 11645 15608 11679
rect 15945 11645 15979 11679
rect 16037 11645 16071 11679
rect 2053 11577 2087 11611
rect 2789 11577 2823 11611
rect 3709 11577 3743 11611
rect 4537 11577 4571 11611
rect 7113 11577 7147 11611
rect 7205 11577 7239 11611
rect 8769 11577 8803 11611
rect 14841 11577 14875 11611
rect 2145 11509 2179 11543
rect 4905 11509 4939 11543
rect 7481 11509 7515 11543
rect 10241 11509 10275 11543
rect 10793 11509 10827 11543
rect 15577 11509 15611 11543
rect 2513 11305 2547 11339
rect 8033 11305 8067 11339
rect 11345 11305 11379 11339
rect 16589 11305 16623 11339
rect 1961 11237 1995 11271
rect 13829 11237 13863 11271
rect 15117 11237 15151 11271
rect 1501 11169 1535 11203
rect 2053 11169 2087 11203
rect 2513 11169 2547 11203
rect 7205 11169 7239 11203
rect 7297 11169 7331 11203
rect 7573 11169 7607 11203
rect 8217 11169 8251 11203
rect 8309 11169 8343 11203
rect 9597 11169 9631 11203
rect 14841 11169 14875 11203
rect 2881 11101 2915 11135
rect 4261 11101 4295 11135
rect 4537 11101 4571 11135
rect 7481 11101 7515 11135
rect 8033 11101 8067 11135
rect 9873 11101 9907 11135
rect 11805 11101 11839 11135
rect 12081 11101 12115 11135
rect 7021 11033 7055 11067
rect 6009 10965 6043 10999
rect 2145 10761 2179 10795
rect 3801 10761 3835 10795
rect 4445 10761 4479 10795
rect 5181 10761 5215 10795
rect 7205 10761 7239 10795
rect 10609 10761 10643 10795
rect 12081 10761 12115 10795
rect 12909 10761 12943 10795
rect 2789 10693 2823 10727
rect 8217 10693 8251 10727
rect 1593 10625 1627 10659
rect 3157 10625 3191 10659
rect 4353 10625 4387 10659
rect 4537 10625 4571 10659
rect 8677 10625 8711 10659
rect 8769 10625 8803 10659
rect 14105 10625 14139 10659
rect 15853 10625 15887 10659
rect 3617 10557 3651 10591
rect 4261 10557 4295 10591
rect 5273 10557 5307 10591
rect 5733 10557 5767 10591
rect 7113 10557 7147 10591
rect 9965 10557 9999 10591
rect 10793 10557 10827 10591
rect 10885 10557 10919 10591
rect 11161 10557 11195 10591
rect 12265 10557 12299 10591
rect 13093 10557 13127 10591
rect 13829 10557 13863 10591
rect 1685 10489 1719 10523
rect 10977 10489 11011 10523
rect 1777 10421 1811 10455
rect 2789 10421 2823 10455
rect 5825 10421 5859 10455
rect 8585 10421 8619 10455
rect 10057 10421 10091 10455
rect 1501 10217 1535 10251
rect 6101 10217 6135 10251
rect 9505 10217 9539 10251
rect 14933 10217 14967 10251
rect 15945 10217 15979 10251
rect 16405 10217 16439 10251
rect 2697 10149 2731 10183
rect 4537 10149 4571 10183
rect 4905 10149 4939 10183
rect 10885 10149 10919 10183
rect 11069 10149 11103 10183
rect 12265 10149 12299 10183
rect 1593 10081 1627 10115
rect 2605 10081 2639 10115
rect 3157 10081 3191 10115
rect 4721 10081 4755 10115
rect 5641 10081 5675 10115
rect 6285 10081 6319 10115
rect 7389 10081 7423 10115
rect 7481 10081 7515 10115
rect 8033 10081 8067 10115
rect 8217 10081 8251 10115
rect 9781 10081 9815 10115
rect 10241 10081 10275 10115
rect 10701 10081 10735 10115
rect 11529 10081 11563 10115
rect 11713 10081 11747 10115
rect 12449 10081 12483 10115
rect 13277 10081 13311 10115
rect 14749 10081 14783 10115
rect 16589 10081 16623 10115
rect 6377 10013 6411 10047
rect 6469 10013 6503 10047
rect 6561 10013 6595 10047
rect 9873 10013 9907 10047
rect 15577 10013 15611 10047
rect 7297 9945 7331 9979
rect 9965 9945 9999 9979
rect 15945 9945 15979 9979
rect 5549 9877 5583 9911
rect 8033 9877 8067 9911
rect 8401 9877 8435 9911
rect 10057 9877 10091 9911
rect 11621 9877 11655 9911
rect 12633 9877 12667 9911
rect 13093 9877 13127 9911
rect 3709 9673 3743 9707
rect 9321 9673 9355 9707
rect 15669 9673 15703 9707
rect 16221 9673 16255 9707
rect 2605 9605 2639 9639
rect 2053 9537 2087 9571
rect 4261 9537 4295 9571
rect 3617 9469 3651 9503
rect 4813 9469 4847 9503
rect 4997 9469 5031 9503
rect 8125 9469 8159 9503
rect 8217 9469 8251 9503
rect 8401 9469 8435 9503
rect 9965 9537 9999 9571
rect 10517 9537 10551 9571
rect 10701 9537 10735 9571
rect 12725 9537 12759 9571
rect 12909 9537 12943 9571
rect 15025 9537 15059 9571
rect 9597 9469 9631 9503
rect 10793 9469 10827 9503
rect 12173 9469 12207 9503
rect 13001 9469 13035 9503
rect 13829 9469 13863 9503
rect 14197 9469 14231 9503
rect 16405 9469 16439 9503
rect 1777 9401 1811 9435
rect 2789 9401 2823 9435
rect 6837 9401 6871 9435
rect 7021 9401 7055 9435
rect 7205 9401 7239 9435
rect 9321 9401 9355 9435
rect 9413 9401 9447 9435
rect 15301 9401 15335 9435
rect 1409 9333 1443 9367
rect 1869 9333 1903 9367
rect 8585 9333 8619 9367
rect 11161 9333 11195 9367
rect 11989 9333 12023 9367
rect 13369 9333 13403 9367
rect 14197 9333 14231 9367
rect 15209 9333 15243 9367
rect 2237 9129 2271 9163
rect 5733 9129 5767 9163
rect 8585 9129 8619 9163
rect 12357 9129 12391 9163
rect 12725 9129 12759 9163
rect 14749 9129 14783 9163
rect 5089 9061 5123 9095
rect 11345 9061 11379 9095
rect 13737 9061 13771 9095
rect 15945 9061 15979 9095
rect 5917 8993 5951 9027
rect 6101 8993 6135 9027
rect 6745 8993 6779 9027
rect 6929 8993 6963 9027
rect 7389 8993 7423 9027
rect 8401 8993 8435 9027
rect 9505 8993 9539 9027
rect 9781 8993 9815 9027
rect 9965 8993 9999 9027
rect 12265 8993 12299 9027
rect 13277 8993 13311 9027
rect 13829 8993 13863 9027
rect 14933 8993 14967 9027
rect 15485 8993 15519 9027
rect 16037 8993 16071 9027
rect 1869 8925 1903 8959
rect 2789 8925 2823 8959
rect 3157 8925 3191 8959
rect 5089 8925 5123 8959
rect 5181 8925 5215 8959
rect 7665 8925 7699 8959
rect 8125 8925 8159 8959
rect 11345 8925 11379 8959
rect 11437 8925 11471 8959
rect 12173 8925 12207 8959
rect 2237 8857 2271 8891
rect 6561 8857 6595 8891
rect 8217 8857 8251 8891
rect 9873 8857 9907 8891
rect 10241 8857 10275 8891
rect 2789 8789 2823 8823
rect 4629 8789 4663 8823
rect 6009 8789 6043 8823
rect 7481 8789 7515 8823
rect 7573 8789 7607 8823
rect 9689 8789 9723 8823
rect 10885 8789 10919 8823
rect 2605 8585 2639 8619
rect 5365 8585 5399 8619
rect 12449 8585 12483 8619
rect 14657 8585 14691 8619
rect 11805 8517 11839 8551
rect 4629 8449 4663 8483
rect 4813 8449 4847 8483
rect 5641 8449 5675 8483
rect 5825 8449 5859 8483
rect 7665 8449 7699 8483
rect 10057 8449 10091 8483
rect 10333 8449 10367 8483
rect 13001 8449 13035 8483
rect 2605 8381 2639 8415
rect 3157 8381 3191 8415
rect 4537 8381 4571 8415
rect 5549 8381 5583 8415
rect 5733 8381 5767 8415
rect 7481 8381 7515 8415
rect 7573 8381 7607 8415
rect 7757 8381 7791 8415
rect 8769 8381 8803 8415
rect 10241 8381 10275 8415
rect 10425 8381 10459 8415
rect 10517 8381 10551 8415
rect 11989 8381 12023 8415
rect 14105 8381 14139 8415
rect 14841 8381 14875 8415
rect 15301 8381 15335 8415
rect 15669 8381 15703 8415
rect 16221 8381 16255 8415
rect 1409 8313 1443 8347
rect 1593 8313 1627 8347
rect 9413 8313 9447 8347
rect 12909 8313 12943 8347
rect 13921 8313 13955 8347
rect 16129 8313 16163 8347
rect 4169 8245 4203 8279
rect 7941 8245 7975 8279
rect 12817 8245 12851 8279
rect 15669 8245 15703 8279
rect 2697 8041 2731 8075
rect 3157 8041 3191 8075
rect 5825 8041 5859 8075
rect 11437 8041 11471 8075
rect 12725 8041 12759 8075
rect 14657 8041 14691 8075
rect 16405 8041 16439 8075
rect 1869 7973 1903 8007
rect 2513 7973 2547 8007
rect 8401 7973 8435 8007
rect 9657 7973 9691 8007
rect 9873 7973 9907 8007
rect 15761 7973 15795 8007
rect 1409 7905 1443 7939
rect 1961 7905 1995 7939
rect 3341 7905 3375 7939
rect 4261 7905 4295 7939
rect 5181 7905 5215 7939
rect 7113 7905 7147 7939
rect 7573 7905 7607 7939
rect 8493 7905 8527 7939
rect 8953 7905 8987 7939
rect 10333 7905 10367 7939
rect 11161 7905 11195 7939
rect 11253 7905 11287 7939
rect 12081 7905 12115 7939
rect 12541 7905 12575 7939
rect 13185 7905 13219 7939
rect 13737 7905 13771 7939
rect 14841 7905 14875 7939
rect 15289 7905 15323 7939
rect 15853 7905 15887 7939
rect 16589 7905 16623 7939
rect 5733 7837 5767 7871
rect 5917 7837 5951 7871
rect 6837 7837 6871 7871
rect 7665 7837 7699 7871
rect 7849 7837 7883 7871
rect 5089 7769 5123 7803
rect 7021 7769 7055 7803
rect 9505 7769 9539 7803
rect 11897 7769 11931 7803
rect 4353 7701 4387 7735
rect 6285 7701 6319 7735
rect 6929 7701 6963 7735
rect 7757 7701 7791 7735
rect 8953 7701 8987 7735
rect 9689 7701 9723 7735
rect 10425 7701 10459 7735
rect 13737 7701 13771 7735
rect 2513 7497 2547 7531
rect 6837 7497 6871 7531
rect 8493 7497 8527 7531
rect 10333 7497 10367 7531
rect 13277 7497 13311 7531
rect 16221 7497 16255 7531
rect 5825 7429 5859 7463
rect 12173 7429 12207 7463
rect 15025 7429 15059 7463
rect 5457 7361 5491 7395
rect 7021 7361 7055 7395
rect 7297 7361 7331 7395
rect 12541 7361 12575 7395
rect 13829 7361 13863 7395
rect 1409 7293 1443 7327
rect 3709 7293 3743 7327
rect 4261 7293 4295 7327
rect 7113 7293 7147 7327
rect 7205 7293 7239 7327
rect 8309 7293 8343 7327
rect 8585 7293 8619 7327
rect 9045 7293 9079 7327
rect 10885 7293 10919 7327
rect 15209 7293 15243 7327
rect 16405 7293 16439 7327
rect 2605 7225 2639 7259
rect 4169 7225 4203 7259
rect 5273 7225 5307 7259
rect 9781 7225 9815 7259
rect 9873 7225 9907 7259
rect 10057 7225 10091 7259
rect 12725 7225 12759 7259
rect 1593 7157 1627 7191
rect 5365 7157 5399 7191
rect 8125 7157 8159 7191
rect 9137 7157 9171 7191
rect 11069 7157 11103 7191
rect 12633 7157 12667 7191
rect 13645 7157 13679 7191
rect 13737 7157 13771 7191
rect 2053 6953 2087 6987
rect 8217 6953 8251 6987
rect 12909 6953 12943 6987
rect 13829 6953 13863 6987
rect 16405 6953 16439 6987
rect 1961 6885 1995 6919
rect 12725 6885 12759 6919
rect 2973 6817 3007 6851
rect 4813 6817 4847 6851
rect 5733 6817 5767 6851
rect 5917 6817 5951 6851
rect 6009 6817 6043 6851
rect 6653 6817 6687 6851
rect 7389 6817 7423 6851
rect 9689 6817 9723 6851
rect 11161 6817 11195 6851
rect 11345 6817 11379 6851
rect 12081 6817 12115 6851
rect 12541 6817 12575 6851
rect 13461 6817 13495 6851
rect 13829 6817 13863 6851
rect 14841 6817 14875 6851
rect 15669 6817 15703 6851
rect 16313 6817 16347 6851
rect 2237 6749 2271 6783
rect 3341 6749 3375 6783
rect 4261 6749 4295 6783
rect 8033 6749 8067 6783
rect 8125 6749 8159 6783
rect 10149 6749 10183 6783
rect 10701 6749 10735 6783
rect 4353 6681 4387 6715
rect 6469 6681 6503 6715
rect 10241 6681 10275 6715
rect 15025 6681 15059 6715
rect 1593 6613 1627 6647
rect 3341 6613 3375 6647
rect 5549 6613 5583 6647
rect 7205 6613 7239 6647
rect 8585 6613 8619 6647
rect 9505 6613 9539 6647
rect 15485 6613 15519 6647
rect 4445 6409 4479 6443
rect 5457 6409 5491 6443
rect 8401 6409 8435 6443
rect 9045 6409 9079 6443
rect 13461 6409 13495 6443
rect 14197 6409 14231 6443
rect 15393 6409 15427 6443
rect 16221 6409 16255 6443
rect 12081 6341 12115 6375
rect 1777 6273 1811 6307
rect 5917 6273 5951 6307
rect 7297 6273 7331 6307
rect 7481 6273 7515 6307
rect 12449 6273 12483 6307
rect 15853 6273 15887 6307
rect 1961 6205 1995 6239
rect 3249 6205 3283 6239
rect 3893 6205 3927 6239
rect 4629 6205 4663 6239
rect 5641 6205 5675 6239
rect 5825 6205 5859 6239
rect 8309 6205 8343 6239
rect 8493 6205 8527 6239
rect 8953 6205 8987 6239
rect 9229 6205 9263 6239
rect 9873 6205 9907 6239
rect 10425 6205 10459 6239
rect 10977 6205 11011 6239
rect 13553 6205 13587 6239
rect 14381 6205 14415 6239
rect 14841 6205 14875 6239
rect 15393 6205 15427 6239
rect 16221 6205 16255 6239
rect 1869 6137 1903 6171
rect 2973 6137 3007 6171
rect 10333 6137 10367 6171
rect 2329 6069 2363 6103
rect 6837 6069 6871 6103
rect 7205 6069 7239 6103
rect 8125 6069 8159 6103
rect 9413 6069 9447 6103
rect 11161 6069 11195 6103
rect 12081 6069 12115 6103
rect 2237 5865 2271 5899
rect 4537 5865 4571 5899
rect 6285 5865 6319 5899
rect 13645 5865 13679 5899
rect 6377 5797 6411 5831
rect 13001 5797 13035 5831
rect 1869 5729 1903 5763
rect 2697 5729 2731 5763
rect 4629 5729 4663 5763
rect 4813 5729 4847 5763
rect 7481 5729 7515 5763
rect 8217 5729 8251 5763
rect 9505 5729 9539 5763
rect 11161 5729 11195 5763
rect 11621 5729 11655 5763
rect 12173 5729 12207 5763
rect 13829 5729 13863 5763
rect 14749 5729 14783 5763
rect 15209 5729 15243 5763
rect 5273 5661 5307 5695
rect 6469 5661 6503 5695
rect 7757 5661 7791 5695
rect 10149 5661 10183 5695
rect 10517 5661 10551 5695
rect 13093 5661 13127 5695
rect 14381 5661 14415 5695
rect 15853 5661 15887 5695
rect 16221 5661 16255 5695
rect 2237 5593 2271 5627
rect 2881 5593 2915 5627
rect 8309 5593 8343 5627
rect 10977 5593 11011 5627
rect 15393 5593 15427 5627
rect 5917 5525 5951 5559
rect 7297 5525 7331 5559
rect 7665 5525 7699 5559
rect 9689 5525 9723 5559
rect 10149 5525 10183 5559
rect 12173 5525 12207 5559
rect 14381 5525 14415 5559
rect 15853 5525 15887 5559
rect 2329 5321 2363 5355
rect 2789 5321 2823 5355
rect 7389 5321 7423 5355
rect 10241 5321 10275 5355
rect 12725 5321 12759 5355
rect 9781 5253 9815 5287
rect 4445 5185 4479 5219
rect 8033 5185 8067 5219
rect 9137 5185 9171 5219
rect 14381 5185 14415 5219
rect 15485 5185 15519 5219
rect 1777 5117 1811 5151
rect 2329 5117 2363 5151
rect 2973 5117 3007 5151
rect 3985 5117 4019 5151
rect 5273 5117 5307 5151
rect 6837 5117 6871 5151
rect 7389 5117 7423 5151
rect 8217 5117 8251 5151
rect 9413 5117 9447 5151
rect 10241 5117 10275 5151
rect 10793 5117 10827 5151
rect 12265 5117 12299 5151
rect 12725 5117 12759 5151
rect 13277 5117 13311 5151
rect 14473 5117 14507 5151
rect 14749 5117 14783 5151
rect 15301 5117 15335 5151
rect 15853 5117 15887 5151
rect 5089 5049 5123 5083
rect 14197 5049 14231 5083
rect 3801 4981 3835 5015
rect 8125 4981 8159 5015
rect 8585 4981 8619 5015
rect 9321 4981 9355 5015
rect 12081 4981 12115 5015
rect 9413 4777 9447 4811
rect 10241 4777 10275 4811
rect 12081 4777 12115 4811
rect 15025 4777 15059 4811
rect 15485 4777 15519 4811
rect 16313 4777 16347 4811
rect 4629 4709 4663 4743
rect 11253 4709 11287 4743
rect 15117 4709 15151 4743
rect 1777 4641 1811 4675
rect 2329 4641 2363 4675
rect 3157 4641 3191 4675
rect 4905 4641 4939 4675
rect 5549 4641 5583 4675
rect 6009 4641 6043 4675
rect 6837 4641 6871 4675
rect 7573 4641 7607 4675
rect 8033 4641 8067 4675
rect 8585 4641 8619 4675
rect 9597 4641 9631 4675
rect 11069 4641 11103 4675
rect 11713 4641 11747 4675
rect 12081 4641 12115 4675
rect 13277 4641 13311 4675
rect 13553 4641 13587 4675
rect 16221 4641 16255 4675
rect 2789 4573 2823 4607
rect 6745 4573 6779 4607
rect 12909 4573 12943 4607
rect 13093 4573 13127 4607
rect 14841 4573 14875 4607
rect 2329 4437 2363 4471
rect 2789 4437 2823 4471
rect 7389 4437 7423 4471
rect 8033 4437 8067 4471
rect 10149 4437 10183 4471
rect 16297 4233 16331 4267
rect 7205 4165 7239 4199
rect 7849 4165 7883 4199
rect 1409 4097 1443 4131
rect 2697 4097 2731 4131
rect 4721 4097 4755 4131
rect 5273 4097 5307 4131
rect 6837 4097 6871 4131
rect 8585 4097 8619 4131
rect 8953 4097 8987 4131
rect 11161 4097 11195 4131
rect 12541 4097 12575 4131
rect 12725 4097 12759 4131
rect 14565 4097 14599 4131
rect 2605 4029 2639 4063
rect 4169 4029 4203 4063
rect 5457 4029 5491 4063
rect 5641 4029 5675 4063
rect 8033 4029 8067 4063
rect 9597 4029 9631 4063
rect 10241 4029 10275 4063
rect 13737 4029 13771 4063
rect 14289 4029 14323 4063
rect 1593 3961 1627 3995
rect 10977 3961 11011 3995
rect 7205 3893 7239 3927
rect 8953 3893 8987 3927
rect 9413 3893 9447 3927
rect 10057 3893 10091 3927
rect 12081 3893 12115 3927
rect 12449 3893 12483 3927
rect 13645 3893 13679 3927
rect 1777 3689 1811 3723
rect 11437 3689 11471 3723
rect 12449 3689 12483 3723
rect 16037 3689 16071 3723
rect 3157 3621 3191 3655
rect 3341 3621 3375 3655
rect 7481 3621 7515 3655
rect 7757 3621 7791 3655
rect 11345 3621 11379 3655
rect 12909 3621 12943 3655
rect 1593 3553 1627 3587
rect 2386 3553 2420 3587
rect 6837 3553 6871 3587
rect 8217 3553 8251 3587
rect 8585 3553 8619 3587
rect 9505 3553 9539 3587
rect 10057 3553 10091 3587
rect 12817 3553 12851 3587
rect 13645 3553 13679 3587
rect 15117 3553 15151 3587
rect 15945 3553 15979 3587
rect 16221 3553 16255 3587
rect 16405 3553 16439 3587
rect 6101 3485 6135 3519
rect 6377 3485 6411 3519
rect 9873 3485 9907 3519
rect 11621 3485 11655 3519
rect 13001 3485 13035 3519
rect 15209 3485 15243 3519
rect 15393 3485 15427 3519
rect 13737 3417 13771 3451
rect 2283 3349 2317 3383
rect 4369 3349 4403 3383
rect 8585 3349 8619 3383
rect 10977 3349 11011 3383
rect 14749 3349 14783 3383
rect 9597 3145 9631 3179
rect 10793 3145 10827 3179
rect 13185 3145 13219 3179
rect 5181 3077 5215 3111
rect 1777 3009 1811 3043
rect 2513 3009 2547 3043
rect 5825 3009 5859 3043
rect 8861 3009 8895 3043
rect 9045 3009 9079 3043
rect 10057 3009 10091 3043
rect 10149 3009 10183 3043
rect 10793 3009 10827 3043
rect 11161 3009 11195 3043
rect 12265 3009 12299 3043
rect 13737 3009 13771 3043
rect 14381 3009 14415 3043
rect 1869 2941 1903 2975
rect 6837 2941 6871 2975
rect 7481 2941 7515 2975
rect 7573 2941 7607 2975
rect 12449 2941 12483 2975
rect 12725 2941 12759 2975
rect 13553 2941 13587 2975
rect 2789 2873 2823 2907
rect 5273 2873 5307 2907
rect 9965 2873 9999 2907
rect 13645 2873 13679 2907
rect 14657 2873 14691 2907
rect 4513 2805 4547 2839
rect 5917 2805 5951 2839
rect 8401 2805 8435 2839
rect 8769 2805 8803 2839
rect 12633 2805 12667 2839
rect 16405 2805 16439 2839
rect 2237 2601 2271 2635
rect 2789 2601 2823 2635
rect 4169 2601 4203 2635
rect 5089 2601 5123 2635
rect 6653 2601 6687 2635
rect 9965 2601 9999 2635
rect 13921 2601 13955 2635
rect 15025 2601 15059 2635
rect 15669 2601 15703 2635
rect 1593 2533 1627 2567
rect 10517 2533 10551 2567
rect 12909 2533 12943 2567
rect 16405 2533 16439 2567
rect 2329 2465 2363 2499
rect 2973 2465 3007 2499
rect 4353 2465 4387 2499
rect 4905 2465 4939 2499
rect 5825 2465 5859 2499
rect 6561 2465 6595 2499
rect 6837 2465 6871 2499
rect 7297 2465 7331 2499
rect 7849 2465 7883 2499
rect 8401 2465 8435 2499
rect 9597 2465 9631 2499
rect 9965 2465 9999 2499
rect 10425 2465 10459 2499
rect 10977 2465 11011 2499
rect 12541 2465 12575 2499
rect 13829 2465 13863 2499
rect 15209 2465 15243 2499
rect 15853 2465 15887 2499
rect 1409 2329 1443 2363
rect 6009 2329 6043 2363
rect 7481 2397 7515 2431
rect 8585 2397 8619 2431
rect 16589 2329 16623 2363
rect 6561 2261 6595 2295
<< metal1 >>
rect 2314 18028 2320 18080
rect 2372 18068 2378 18080
rect 8754 18068 8760 18080
rect 2372 18040 8760 18068
rect 2372 18028 2378 18040
rect 8754 18028 8760 18040
rect 8812 18028 8818 18080
rect 1104 17978 17296 18000
rect 1104 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 6571 17978
rect 6623 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 11904 17978
rect 11956 17926 11968 17978
rect 12020 17926 17296 17978
rect 1104 17904 17296 17926
rect 1486 17864 1492 17876
rect 1447 17836 1492 17864
rect 1486 17824 1492 17836
rect 1544 17824 1550 17876
rect 2133 17867 2191 17873
rect 2133 17864 2145 17867
rect 1596 17836 2145 17864
rect 1596 17805 1624 17836
rect 2133 17833 2145 17836
rect 2179 17833 2191 17867
rect 3418 17864 3424 17876
rect 2133 17827 2191 17833
rect 2332 17836 3424 17864
rect 1581 17799 1639 17805
rect 1581 17765 1593 17799
rect 1627 17765 1639 17799
rect 1581 17759 1639 17765
rect 2332 17737 2360 17836
rect 3418 17824 3424 17836
rect 3476 17824 3482 17876
rect 15654 17864 15660 17876
rect 7024 17836 15660 17864
rect 5994 17796 6000 17808
rect 3160 17768 6000 17796
rect 3160 17737 3188 17768
rect 5994 17756 6000 17768
rect 6052 17756 6058 17808
rect 2317 17731 2375 17737
rect 2317 17697 2329 17731
rect 2363 17697 2375 17731
rect 2317 17691 2375 17697
rect 3145 17731 3203 17737
rect 3145 17697 3157 17731
rect 3191 17697 3203 17731
rect 3145 17691 3203 17697
rect 4617 17731 4675 17737
rect 4617 17697 4629 17731
rect 4663 17697 4675 17731
rect 4617 17691 4675 17697
rect 5445 17731 5503 17737
rect 5445 17697 5457 17731
rect 5491 17697 5503 17731
rect 5445 17691 5503 17697
rect 1762 17620 1768 17672
rect 1820 17660 1826 17672
rect 4632 17660 4660 17691
rect 5350 17660 5356 17672
rect 1820 17632 5356 17660
rect 1820 17620 1826 17632
rect 5350 17620 5356 17632
rect 5408 17620 5414 17672
rect 5460 17660 5488 17691
rect 5534 17688 5540 17740
rect 5592 17728 5598 17740
rect 7024 17737 7052 17836
rect 15654 17824 15660 17836
rect 15712 17824 15718 17876
rect 14274 17796 14280 17808
rect 7668 17768 10548 17796
rect 7668 17740 7696 17768
rect 5629 17731 5687 17737
rect 5629 17728 5641 17731
rect 5592 17700 5641 17728
rect 5592 17688 5598 17700
rect 5629 17697 5641 17700
rect 5675 17697 5687 17731
rect 5629 17691 5687 17697
rect 7009 17731 7067 17737
rect 7009 17697 7021 17731
rect 7055 17697 7067 17731
rect 7650 17728 7656 17740
rect 7611 17700 7656 17728
rect 7009 17691 7067 17697
rect 7650 17688 7656 17700
rect 7708 17688 7714 17740
rect 8478 17728 8484 17740
rect 8439 17700 8484 17728
rect 8478 17688 8484 17700
rect 8536 17688 8542 17740
rect 9582 17728 9588 17740
rect 9543 17700 9588 17728
rect 9582 17688 9588 17700
rect 9640 17688 9646 17740
rect 9766 17728 9772 17740
rect 9727 17700 9772 17728
rect 9766 17688 9772 17700
rect 9824 17688 9830 17740
rect 10520 17737 10548 17768
rect 12360 17768 14280 17796
rect 12360 17737 12388 17768
rect 14274 17756 14280 17768
rect 14332 17756 14338 17808
rect 14918 17756 14924 17808
rect 14976 17796 14982 17808
rect 15013 17799 15071 17805
rect 15013 17796 15025 17799
rect 14976 17768 15025 17796
rect 14976 17756 14982 17768
rect 15013 17765 15025 17768
rect 15059 17765 15071 17799
rect 15013 17759 15071 17765
rect 16485 17799 16543 17805
rect 16485 17765 16497 17799
rect 16531 17796 16543 17799
rect 17034 17796 17040 17808
rect 16531 17768 17040 17796
rect 16531 17765 16543 17768
rect 16485 17759 16543 17765
rect 17034 17756 17040 17768
rect 17092 17756 17098 17808
rect 10505 17731 10563 17737
rect 10505 17697 10517 17731
rect 10551 17728 10563 17731
rect 11149 17731 11207 17737
rect 11149 17728 11161 17731
rect 10551 17700 11161 17728
rect 10551 17697 10563 17700
rect 10505 17691 10563 17697
rect 11149 17697 11161 17700
rect 11195 17697 11207 17731
rect 11149 17691 11207 17697
rect 12345 17731 12403 17737
rect 12345 17697 12357 17731
rect 12391 17697 12403 17731
rect 12345 17691 12403 17697
rect 12989 17731 13047 17737
rect 12989 17697 13001 17731
rect 13035 17728 13047 17731
rect 13817 17731 13875 17737
rect 13817 17728 13829 17731
rect 13035 17700 13829 17728
rect 13035 17697 13047 17700
rect 12989 17691 13047 17697
rect 13817 17697 13829 17700
rect 13863 17697 13875 17731
rect 14737 17731 14795 17737
rect 14737 17728 14749 17731
rect 13817 17691 13875 17697
rect 13924 17700 14749 17728
rect 5718 17660 5724 17672
rect 5460 17632 5724 17660
rect 5718 17620 5724 17632
rect 5776 17620 5782 17672
rect 11164 17660 11192 17691
rect 12434 17660 12440 17672
rect 11164 17632 12440 17660
rect 12434 17620 12440 17632
rect 12492 17660 12498 17672
rect 13004 17660 13032 17691
rect 12492 17632 13032 17660
rect 12492 17620 12498 17632
rect 13078 17620 13084 17672
rect 13136 17660 13142 17672
rect 13924 17660 13952 17700
rect 14737 17697 14749 17700
rect 14783 17697 14795 17731
rect 14737 17691 14795 17697
rect 14826 17688 14832 17740
rect 14884 17728 14890 17740
rect 15657 17731 15715 17737
rect 14884 17700 14929 17728
rect 14884 17688 14890 17700
rect 15657 17697 15669 17731
rect 15703 17728 15715 17731
rect 16022 17728 16028 17740
rect 15703 17700 16028 17728
rect 15703 17697 15715 17700
rect 15657 17691 15715 17697
rect 16022 17688 16028 17700
rect 16080 17688 16086 17740
rect 13136 17632 13952 17660
rect 14553 17663 14611 17669
rect 13136 17620 13142 17632
rect 14553 17629 14565 17663
rect 14599 17660 14611 17663
rect 15562 17660 15568 17672
rect 14599 17632 15568 17660
rect 14599 17629 14611 17632
rect 14553 17623 14611 17629
rect 15562 17620 15568 17632
rect 15620 17620 15626 17672
rect 3329 17595 3387 17601
rect 3329 17561 3341 17595
rect 3375 17592 3387 17595
rect 5626 17592 5632 17604
rect 3375 17564 5632 17592
rect 3375 17561 3387 17564
rect 3329 17555 3387 17561
rect 5626 17552 5632 17564
rect 5684 17552 5690 17604
rect 7193 17595 7251 17601
rect 7193 17561 7205 17595
rect 7239 17592 7251 17595
rect 10689 17595 10747 17601
rect 7239 17564 10640 17592
rect 7239 17561 7251 17564
rect 7193 17555 7251 17561
rect 4798 17524 4804 17536
rect 4759 17496 4804 17524
rect 4798 17484 4804 17496
rect 4856 17484 4862 17536
rect 5258 17524 5264 17536
rect 5219 17496 5264 17524
rect 5258 17484 5264 17496
rect 5316 17484 5322 17536
rect 7834 17524 7840 17536
rect 7795 17496 7840 17524
rect 7834 17484 7840 17496
rect 7892 17484 7898 17536
rect 8386 17524 8392 17536
rect 8347 17496 8392 17524
rect 8386 17484 8392 17496
rect 8444 17484 8450 17536
rect 9674 17524 9680 17536
rect 9635 17496 9680 17524
rect 9674 17484 9680 17496
rect 9732 17484 9738 17536
rect 10612 17524 10640 17564
rect 10689 17561 10701 17595
rect 10735 17592 10747 17595
rect 15102 17592 15108 17604
rect 10735 17564 15108 17592
rect 10735 17561 10747 17564
rect 10689 17555 10747 17561
rect 15102 17552 15108 17564
rect 15160 17552 15166 17604
rect 16114 17552 16120 17604
rect 16172 17592 16178 17604
rect 16301 17595 16359 17601
rect 16301 17592 16313 17595
rect 16172 17564 16313 17592
rect 16172 17552 16178 17564
rect 16301 17561 16313 17564
rect 16347 17561 16359 17595
rect 16301 17555 16359 17561
rect 11054 17524 11060 17536
rect 10612 17496 11060 17524
rect 11054 17484 11060 17496
rect 11112 17484 11118 17536
rect 11330 17524 11336 17536
rect 11291 17496 11336 17524
rect 11330 17484 11336 17496
rect 11388 17484 11394 17536
rect 12526 17524 12532 17536
rect 12487 17496 12532 17524
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 13170 17524 13176 17536
rect 13131 17496 13176 17524
rect 13170 17484 13176 17496
rect 13228 17484 13234 17536
rect 14001 17527 14059 17533
rect 14001 17493 14013 17527
rect 14047 17524 14059 17527
rect 14553 17527 14611 17533
rect 14553 17524 14565 17527
rect 14047 17496 14565 17524
rect 14047 17493 14059 17496
rect 14001 17487 14059 17493
rect 14553 17493 14565 17496
rect 14599 17493 14611 17527
rect 15010 17524 15016 17536
rect 14971 17496 15016 17524
rect 14553 17487 14611 17493
rect 15010 17484 15016 17496
rect 15068 17484 15074 17536
rect 15746 17524 15752 17536
rect 15707 17496 15752 17524
rect 15746 17484 15752 17496
rect 15804 17484 15810 17536
rect 1104 17434 17296 17456
rect 1104 17382 3680 17434
rect 3732 17382 3744 17434
rect 3796 17382 3808 17434
rect 3860 17382 3872 17434
rect 3924 17382 9078 17434
rect 9130 17382 9142 17434
rect 9194 17382 9206 17434
rect 9258 17382 9270 17434
rect 9322 17382 14475 17434
rect 14527 17382 14539 17434
rect 14591 17382 14603 17434
rect 14655 17382 14667 17434
rect 14719 17382 17296 17434
rect 1104 17360 17296 17382
rect 6914 17280 6920 17332
rect 6972 17320 6978 17332
rect 10410 17320 10416 17332
rect 6972 17292 10416 17320
rect 6972 17280 6978 17292
rect 10410 17280 10416 17292
rect 10468 17280 10474 17332
rect 12526 17280 12532 17332
rect 12584 17320 12590 17332
rect 14626 17323 14684 17329
rect 14626 17320 14638 17323
rect 12584 17292 14638 17320
rect 12584 17280 12590 17292
rect 14626 17289 14638 17292
rect 14672 17289 14684 17323
rect 14626 17283 14684 17289
rect 2869 17255 2927 17261
rect 2869 17221 2881 17255
rect 2915 17252 2927 17255
rect 2958 17252 2964 17264
rect 2915 17224 2964 17252
rect 2915 17221 2927 17224
rect 2869 17215 2927 17221
rect 2958 17212 2964 17224
rect 3016 17212 3022 17264
rect 5169 17255 5227 17261
rect 5169 17221 5181 17255
rect 5215 17252 5227 17255
rect 5718 17252 5724 17264
rect 5215 17224 5724 17252
rect 5215 17221 5227 17224
rect 5169 17215 5227 17221
rect 5718 17212 5724 17224
rect 5776 17212 5782 17264
rect 3326 17184 3332 17196
rect 2884 17156 3332 17184
rect 1762 17116 1768 17128
rect 1723 17088 1768 17116
rect 1762 17076 1768 17088
rect 1820 17076 1826 17128
rect 2593 17119 2651 17125
rect 2593 17085 2605 17119
rect 2639 17085 2651 17119
rect 2593 17079 2651 17085
rect 2731 17119 2789 17125
rect 2731 17085 2743 17119
rect 2777 17116 2789 17119
rect 2884 17116 2912 17156
rect 3326 17144 3332 17156
rect 3384 17144 3390 17196
rect 3697 17187 3755 17193
rect 3697 17153 3709 17187
rect 3743 17184 3755 17187
rect 5258 17184 5264 17196
rect 3743 17156 5264 17184
rect 3743 17153 3755 17156
rect 3697 17147 3755 17153
rect 5258 17144 5264 17156
rect 5316 17144 5322 17196
rect 8021 17187 8079 17193
rect 8021 17153 8033 17187
rect 8067 17184 8079 17187
rect 13633 17187 13691 17193
rect 8067 17156 10548 17184
rect 8067 17153 8079 17156
rect 8021 17147 8079 17153
rect 10520 17128 10548 17156
rect 13633 17153 13645 17187
rect 13679 17184 13691 17187
rect 15010 17184 15016 17196
rect 13679 17156 15016 17184
rect 13679 17153 13691 17156
rect 13633 17147 13691 17153
rect 15010 17144 15016 17156
rect 15068 17144 15074 17196
rect 2777 17088 2912 17116
rect 2961 17119 3019 17125
rect 2777 17085 2789 17088
rect 2731 17079 2789 17085
rect 2961 17085 2973 17119
rect 3007 17116 3019 17119
rect 3050 17116 3056 17128
rect 3007 17088 3056 17116
rect 3007 17085 3019 17088
rect 2961 17079 3019 17085
rect 1670 17008 1676 17060
rect 1728 17048 1734 17060
rect 2409 17051 2467 17057
rect 2409 17048 2421 17051
rect 1728 17020 2421 17048
rect 1728 17008 1734 17020
rect 2409 17017 2421 17020
rect 2455 17017 2467 17051
rect 2608 17048 2636 17079
rect 3050 17076 3056 17088
rect 3108 17076 3114 17128
rect 3418 17116 3424 17128
rect 3379 17088 3424 17116
rect 3418 17076 3424 17088
rect 3476 17076 3482 17128
rect 5350 17076 5356 17128
rect 5408 17116 5414 17128
rect 5813 17119 5871 17125
rect 5813 17116 5825 17119
rect 5408 17088 5825 17116
rect 5408 17076 5414 17088
rect 5813 17085 5825 17088
rect 5859 17116 5871 17119
rect 7285 17119 7343 17125
rect 7285 17116 7297 17119
rect 5859 17088 7297 17116
rect 5859 17085 5871 17088
rect 5813 17079 5871 17085
rect 7285 17085 7297 17088
rect 7331 17116 7343 17119
rect 7650 17116 7656 17128
rect 7331 17088 7656 17116
rect 7331 17085 7343 17088
rect 7285 17079 7343 17085
rect 7650 17076 7656 17088
rect 7708 17076 7714 17128
rect 7834 17076 7840 17128
rect 7892 17116 7898 17128
rect 9769 17119 9827 17125
rect 7892 17088 8418 17116
rect 7892 17076 7898 17088
rect 9769 17085 9781 17119
rect 9815 17085 9827 17119
rect 10410 17116 10416 17128
rect 10371 17088 10416 17116
rect 9769 17079 9827 17085
rect 2866 17048 2872 17060
rect 2608 17020 2872 17048
rect 2409 17011 2467 17017
rect 2866 17008 2872 17020
rect 2924 17008 2930 17060
rect 9493 17051 9551 17057
rect 4922 17020 5672 17048
rect 1946 16980 1952 16992
rect 1907 16952 1952 16980
rect 1946 16940 1952 16952
rect 2004 16940 2010 16992
rect 5644 16989 5672 17020
rect 9493 17017 9505 17051
rect 9539 17017 9551 17051
rect 9784 17048 9812 17079
rect 10410 17076 10416 17088
rect 10468 17076 10474 17128
rect 10502 17076 10508 17128
rect 10560 17116 10566 17128
rect 10781 17119 10839 17125
rect 10560 17088 10653 17116
rect 10560 17076 10566 17088
rect 10781 17085 10793 17119
rect 10827 17116 10839 17119
rect 10870 17116 10876 17128
rect 10827 17088 10876 17116
rect 10827 17085 10839 17088
rect 10781 17079 10839 17085
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 13909 17119 13967 17125
rect 13909 17085 13921 17119
rect 13955 17116 13967 17119
rect 14366 17116 14372 17128
rect 13955 17088 14372 17116
rect 13955 17085 13967 17088
rect 13909 17079 13967 17085
rect 14366 17076 14372 17088
rect 14424 17076 14430 17128
rect 9858 17048 9864 17060
rect 9784 17020 9864 17048
rect 9493 17011 9551 17017
rect 5629 16983 5687 16989
rect 5629 16949 5641 16983
rect 5675 16949 5687 16983
rect 5629 16943 5687 16949
rect 7469 16983 7527 16989
rect 7469 16949 7481 16983
rect 7515 16980 7527 16983
rect 7558 16980 7564 16992
rect 7515 16952 7564 16980
rect 7515 16949 7527 16952
rect 7469 16943 7527 16949
rect 7558 16940 7564 16952
rect 7616 16940 7622 16992
rect 9508 16980 9536 17011
rect 9858 17008 9864 17020
rect 9916 17008 9922 17060
rect 10597 17051 10655 17057
rect 10597 17017 10609 17051
rect 10643 17048 10655 17051
rect 11146 17048 11152 17060
rect 10643 17020 11152 17048
rect 10643 17017 10655 17020
rect 10597 17011 10655 17017
rect 11146 17008 11152 17020
rect 11204 17048 11210 17060
rect 11204 17020 12204 17048
rect 11204 17008 11210 17020
rect 12176 16989 12204 17020
rect 13170 17008 13176 17060
rect 13228 17008 13234 17060
rect 15102 17008 15108 17060
rect 15160 17008 15166 17060
rect 10229 16983 10287 16989
rect 10229 16980 10241 16983
rect 9508 16952 10241 16980
rect 10229 16949 10241 16952
rect 10275 16949 10287 16983
rect 10229 16943 10287 16949
rect 12161 16983 12219 16989
rect 12161 16949 12173 16983
rect 12207 16949 12219 16983
rect 12161 16943 12219 16949
rect 12250 16940 12256 16992
rect 12308 16980 12314 16992
rect 14826 16980 14832 16992
rect 12308 16952 14832 16980
rect 12308 16940 12314 16952
rect 14826 16940 14832 16952
rect 14884 16940 14890 16992
rect 15378 16940 15384 16992
rect 15436 16980 15442 16992
rect 16117 16983 16175 16989
rect 16117 16980 16129 16983
rect 15436 16952 16129 16980
rect 15436 16940 15442 16952
rect 16117 16949 16129 16952
rect 16163 16949 16175 16983
rect 16117 16943 16175 16949
rect 1104 16890 17296 16912
rect 1104 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 6571 16890
rect 6623 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 11904 16890
rect 11956 16838 11968 16890
rect 12020 16838 17296 16890
rect 1104 16816 17296 16838
rect 5813 16779 5871 16785
rect 5813 16745 5825 16779
rect 5859 16745 5871 16779
rect 9766 16776 9772 16788
rect 9727 16748 9772 16776
rect 5813 16739 5871 16745
rect 1670 16708 1676 16720
rect 1631 16680 1676 16708
rect 1670 16668 1676 16680
rect 1728 16668 1734 16720
rect 1946 16668 1952 16720
rect 2004 16708 2010 16720
rect 2004 16680 2162 16708
rect 2004 16668 2010 16680
rect 2958 16668 2964 16720
rect 3016 16708 3022 16720
rect 4709 16711 4767 16717
rect 4709 16708 4721 16711
rect 3016 16680 4721 16708
rect 3016 16668 3022 16680
rect 4709 16677 4721 16680
rect 4755 16677 4767 16711
rect 4709 16671 4767 16677
rect 5445 16711 5503 16717
rect 5445 16677 5457 16711
rect 5491 16708 5503 16711
rect 5718 16708 5724 16720
rect 5491 16680 5724 16708
rect 5491 16677 5503 16680
rect 5445 16671 5503 16677
rect 5718 16668 5724 16680
rect 5776 16668 5782 16720
rect 5828 16708 5856 16739
rect 9766 16736 9772 16748
rect 9824 16736 9830 16788
rect 12161 16779 12219 16785
rect 12161 16776 12173 16779
rect 11256 16748 12173 16776
rect 6549 16711 6607 16717
rect 6549 16708 6561 16711
rect 5828 16680 6561 16708
rect 6549 16677 6561 16680
rect 6595 16677 6607 16711
rect 6549 16671 6607 16677
rect 7558 16668 7564 16720
rect 7616 16668 7622 16720
rect 11146 16708 11152 16720
rect 11107 16680 11152 16708
rect 11146 16668 11152 16680
rect 11204 16668 11210 16720
rect 3326 16600 3332 16652
rect 3384 16640 3390 16652
rect 4617 16643 4675 16649
rect 4617 16640 4629 16643
rect 3384 16612 4629 16640
rect 3384 16600 3390 16612
rect 4617 16609 4629 16612
rect 4663 16609 4675 16643
rect 4617 16603 4675 16609
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16609 5319 16643
rect 5261 16603 5319 16609
rect 5537 16643 5595 16649
rect 5537 16609 5549 16643
rect 5583 16609 5595 16643
rect 5537 16603 5595 16609
rect 5629 16643 5687 16649
rect 5629 16609 5641 16643
rect 5675 16640 5687 16643
rect 9858 16640 9864 16652
rect 5675 16612 6224 16640
rect 5675 16609 5687 16612
rect 5629 16603 5687 16609
rect 1394 16572 1400 16584
rect 1355 16544 1400 16572
rect 1394 16532 1400 16544
rect 1452 16532 1458 16584
rect 5276 16504 5304 16603
rect 5552 16572 5580 16603
rect 6086 16572 6092 16584
rect 5552 16544 6092 16572
rect 6086 16532 6092 16544
rect 6144 16532 6150 16584
rect 5534 16504 5540 16516
rect 5276 16476 5540 16504
rect 5534 16464 5540 16476
rect 5592 16504 5598 16516
rect 5994 16504 6000 16516
rect 5592 16476 6000 16504
rect 5592 16464 5598 16476
rect 5994 16464 6000 16476
rect 6052 16464 6058 16516
rect 3050 16396 3056 16448
rect 3108 16436 3114 16448
rect 3145 16439 3203 16445
rect 3145 16436 3157 16439
rect 3108 16408 3157 16436
rect 3108 16396 3114 16408
rect 3145 16405 3157 16408
rect 3191 16405 3203 16439
rect 6196 16436 6224 16612
rect 9646 16612 9864 16640
rect 6273 16575 6331 16581
rect 6273 16541 6285 16575
rect 6319 16572 6331 16575
rect 9646 16572 9674 16612
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 10502 16600 10508 16652
rect 10560 16640 10566 16652
rect 10962 16640 10968 16652
rect 10560 16612 10968 16640
rect 10560 16600 10566 16612
rect 10962 16600 10968 16612
rect 11020 16640 11026 16652
rect 11057 16643 11115 16649
rect 11057 16640 11069 16643
rect 11020 16612 11069 16640
rect 11020 16600 11026 16612
rect 11057 16609 11069 16612
rect 11103 16609 11115 16643
rect 11057 16603 11115 16609
rect 9950 16572 9956 16584
rect 6319 16544 9674 16572
rect 9911 16544 9956 16572
rect 6319 16541 6331 16544
rect 6273 16535 6331 16541
rect 9950 16532 9956 16544
rect 10008 16532 10014 16584
rect 10045 16575 10103 16581
rect 10045 16541 10057 16575
rect 10091 16541 10103 16575
rect 10410 16572 10416 16584
rect 10371 16544 10416 16572
rect 10045 16535 10103 16541
rect 10060 16504 10088 16535
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 11164 16572 11192 16668
rect 11256 16652 11284 16748
rect 12161 16745 12173 16748
rect 12207 16776 12219 16779
rect 12250 16776 12256 16788
rect 12207 16748 12256 16776
rect 12207 16745 12219 16748
rect 12161 16739 12219 16745
rect 12250 16736 12256 16748
rect 12308 16736 12314 16788
rect 12805 16779 12863 16785
rect 12805 16745 12817 16779
rect 12851 16776 12863 16779
rect 13078 16776 13084 16788
rect 12851 16748 13084 16776
rect 12851 16745 12863 16748
rect 12805 16739 12863 16745
rect 13078 16736 13084 16748
rect 13136 16736 13142 16788
rect 11330 16668 11336 16720
rect 11388 16708 11394 16720
rect 11388 16680 15502 16708
rect 11388 16668 11394 16680
rect 11238 16600 11244 16652
rect 11296 16640 11302 16652
rect 11422 16640 11428 16652
rect 11296 16612 11341 16640
rect 11383 16612 11428 16640
rect 11296 16600 11302 16612
rect 11422 16600 11428 16612
rect 11480 16600 11486 16652
rect 12069 16643 12127 16649
rect 12069 16609 12081 16643
rect 12115 16609 12127 16643
rect 12710 16640 12716 16652
rect 12671 16612 12716 16640
rect 12069 16603 12127 16609
rect 12084 16572 12112 16603
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 12802 16600 12808 16652
rect 12860 16640 12866 16652
rect 12897 16643 12955 16649
rect 12897 16640 12909 16643
rect 12860 16612 12909 16640
rect 12860 16600 12866 16612
rect 12897 16609 12909 16612
rect 12943 16609 12955 16643
rect 13357 16643 13415 16649
rect 13357 16640 13369 16643
rect 12897 16603 12955 16609
rect 13004 16612 13369 16640
rect 12158 16572 12164 16584
rect 11164 16544 12164 16572
rect 12158 16532 12164 16544
rect 12216 16532 12222 16584
rect 13004 16572 13032 16612
rect 13357 16609 13369 16612
rect 13403 16609 13415 16643
rect 13357 16603 13415 16609
rect 12452 16544 13032 16572
rect 12452 16516 12480 16544
rect 14366 16532 14372 16584
rect 14424 16572 14430 16584
rect 14737 16575 14795 16581
rect 14737 16572 14749 16575
rect 14424 16544 14749 16572
rect 14424 16532 14430 16544
rect 14737 16541 14749 16544
rect 14783 16541 14795 16575
rect 14737 16535 14795 16541
rect 15013 16575 15071 16581
rect 15013 16541 15025 16575
rect 15059 16572 15071 16575
rect 15378 16572 15384 16584
rect 15059 16544 15384 16572
rect 15059 16541 15071 16544
rect 15013 16535 15071 16541
rect 15378 16532 15384 16544
rect 15436 16532 15442 16584
rect 10226 16504 10232 16516
rect 10060 16476 10232 16504
rect 10226 16464 10232 16476
rect 10284 16504 10290 16516
rect 10873 16507 10931 16513
rect 10873 16504 10885 16507
rect 10284 16476 10885 16504
rect 10284 16464 10290 16476
rect 10873 16473 10885 16476
rect 10919 16473 10931 16507
rect 10873 16467 10931 16473
rect 12342 16464 12348 16516
rect 12400 16504 12406 16516
rect 12434 16504 12440 16516
rect 12400 16476 12440 16504
rect 12400 16464 12406 16476
rect 12434 16464 12440 16476
rect 12492 16464 12498 16516
rect 6914 16436 6920 16448
rect 6196 16408 6920 16436
rect 3145 16399 3203 16405
rect 6914 16396 6920 16408
rect 6972 16396 6978 16448
rect 8018 16436 8024 16448
rect 7979 16408 8024 16436
rect 8018 16396 8024 16408
rect 8076 16396 8082 16448
rect 10134 16396 10140 16448
rect 10192 16436 10198 16448
rect 11514 16436 11520 16448
rect 10192 16408 11520 16436
rect 10192 16396 10198 16408
rect 11514 16396 11520 16408
rect 11572 16396 11578 16448
rect 13446 16396 13452 16448
rect 13504 16436 13510 16448
rect 13541 16439 13599 16445
rect 13541 16436 13553 16439
rect 13504 16408 13553 16436
rect 13504 16396 13510 16408
rect 13541 16405 13553 16408
rect 13587 16405 13599 16439
rect 16482 16436 16488 16448
rect 16443 16408 16488 16436
rect 13541 16399 13599 16405
rect 16482 16396 16488 16408
rect 16540 16396 16546 16448
rect 1104 16346 17296 16368
rect 1104 16294 3680 16346
rect 3732 16294 3744 16346
rect 3796 16294 3808 16346
rect 3860 16294 3872 16346
rect 3924 16294 9078 16346
rect 9130 16294 9142 16346
rect 9194 16294 9206 16346
rect 9258 16294 9270 16346
rect 9322 16294 14475 16346
rect 14527 16294 14539 16346
rect 14591 16294 14603 16346
rect 14655 16294 14667 16346
rect 14719 16294 17296 16346
rect 1104 16272 17296 16294
rect 2866 16232 2872 16244
rect 2827 16204 2872 16232
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 8294 16232 8300 16244
rect 2976 16204 8300 16232
rect 2976 16096 3004 16204
rect 8294 16192 8300 16204
rect 8352 16192 8358 16244
rect 9766 16192 9772 16244
rect 9824 16232 9830 16244
rect 11057 16235 11115 16241
rect 11057 16232 11069 16235
rect 9824 16204 10088 16232
rect 9824 16192 9830 16204
rect 9582 16164 9588 16176
rect 5552 16136 9588 16164
rect 2746 16068 3004 16096
rect 1489 16031 1547 16037
rect 1489 15997 1501 16031
rect 1535 16028 1547 16031
rect 1854 16028 1860 16040
rect 1535 16000 1860 16028
rect 1535 15997 1547 16000
rect 1489 15991 1547 15997
rect 1854 15988 1860 16000
rect 1912 15988 1918 16040
rect 2133 16031 2191 16037
rect 2133 15997 2145 16031
rect 2179 16028 2191 16031
rect 2746 16028 2774 16068
rect 3418 16056 3424 16108
rect 3476 16096 3482 16108
rect 3881 16099 3939 16105
rect 3881 16096 3893 16099
rect 3476 16068 3893 16096
rect 3476 16056 3482 16068
rect 3881 16065 3893 16068
rect 3927 16096 3939 16099
rect 4246 16096 4252 16108
rect 3927 16068 4252 16096
rect 3927 16065 3939 16068
rect 3881 16059 3939 16065
rect 4246 16056 4252 16068
rect 4304 16056 4310 16108
rect 2179 16000 2774 16028
rect 2961 16031 3019 16037
rect 2179 15997 2191 16000
rect 2133 15991 2191 15997
rect 2961 15997 2973 16031
rect 3007 16028 3019 16031
rect 3050 16028 3056 16040
rect 3007 16000 3056 16028
rect 3007 15997 3019 16000
rect 2961 15991 3019 15997
rect 3050 15988 3056 16000
rect 3108 15988 3114 16040
rect 474 15920 480 15972
rect 532 15960 538 15972
rect 1302 15960 1308 15972
rect 532 15932 1308 15960
rect 532 15920 538 15932
rect 1302 15920 1308 15932
rect 1360 15920 1366 15972
rect 4154 15960 4160 15972
rect 4115 15932 4160 15960
rect 4154 15920 4160 15932
rect 4212 15920 4218 15972
rect 4798 15920 4804 15972
rect 4856 15920 4862 15972
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 2317 15895 2375 15901
rect 2317 15861 2329 15895
rect 2363 15892 2375 15895
rect 5552 15892 5580 16136
rect 9582 16124 9588 16136
rect 9640 16164 9646 16176
rect 9640 16136 9812 16164
rect 9640 16124 9646 16136
rect 6086 16056 6092 16108
rect 6144 16096 6150 16108
rect 6270 16096 6276 16108
rect 6144 16068 6276 16096
rect 6144 16056 6150 16068
rect 6270 16056 6276 16068
rect 6328 16096 6334 16108
rect 7469 16099 7527 16105
rect 6328 16068 7420 16096
rect 6328 16056 6334 16068
rect 5718 15988 5724 16040
rect 5776 16028 5782 16040
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 5776 16000 6837 16028
rect 5776 15988 5782 16000
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 6825 15991 6883 15997
rect 7009 16031 7067 16037
rect 7009 15997 7021 16031
rect 7055 15997 7067 16031
rect 7282 16028 7288 16040
rect 7243 16000 7288 16028
rect 7009 15991 7067 15997
rect 6178 15960 6184 15972
rect 5644 15932 6184 15960
rect 5644 15901 5672 15932
rect 6178 15920 6184 15932
rect 6236 15960 6242 15972
rect 7024 15960 7052 15991
rect 7282 15988 7288 16000
rect 7340 15988 7346 16040
rect 7392 16028 7420 16068
rect 7469 16065 7481 16099
rect 7515 16096 7527 16099
rect 8662 16096 8668 16108
rect 7515 16068 8432 16096
rect 8623 16068 8668 16096
rect 7515 16065 7527 16068
rect 7469 16059 7527 16065
rect 7653 16031 7711 16037
rect 7653 16028 7665 16031
rect 7392 16000 7665 16028
rect 7653 15997 7665 16000
rect 7699 16028 7711 16031
rect 8018 16028 8024 16040
rect 7699 16000 8024 16028
rect 7699 15997 7711 16000
rect 7653 15991 7711 15997
rect 8018 15988 8024 16000
rect 8076 15988 8082 16040
rect 8404 16037 8432 16068
rect 8662 16056 8668 16068
rect 8720 16056 8726 16108
rect 8849 16099 8907 16105
rect 8849 16065 8861 16099
rect 8895 16096 8907 16099
rect 9674 16096 9680 16108
rect 8895 16068 9680 16096
rect 8895 16065 8907 16068
rect 8849 16059 8907 16065
rect 9674 16056 9680 16068
rect 9732 16056 9738 16108
rect 9784 16096 9812 16136
rect 10060 16105 10088 16204
rect 10152 16204 11069 16232
rect 10152 16105 10180 16204
rect 11057 16201 11069 16204
rect 11103 16232 11115 16235
rect 11422 16232 11428 16244
rect 11103 16204 11428 16232
rect 11103 16201 11115 16204
rect 11057 16195 11115 16201
rect 11422 16192 11428 16204
rect 11480 16192 11486 16244
rect 12710 16192 12716 16244
rect 12768 16232 12774 16244
rect 13170 16232 13176 16244
rect 12768 16204 13176 16232
rect 12768 16192 12774 16204
rect 13170 16192 13176 16204
rect 13228 16232 13234 16244
rect 14185 16235 14243 16241
rect 14185 16232 14197 16235
rect 13228 16204 14197 16232
rect 13228 16192 13234 16204
rect 14185 16201 14197 16204
rect 14231 16201 14243 16235
rect 14185 16195 14243 16201
rect 11238 16164 11244 16176
rect 10336 16136 11244 16164
rect 10045 16099 10103 16105
rect 9784 16068 9996 16096
rect 8389 16031 8447 16037
rect 8389 15997 8401 16031
rect 8435 15997 8447 16031
rect 8389 15991 8447 15997
rect 8478 15988 8484 16040
rect 8536 16028 8542 16040
rect 9766 16028 9772 16040
rect 8536 16000 8629 16028
rect 9727 16000 9772 16028
rect 8536 15988 8542 16000
rect 9766 15988 9772 16000
rect 9824 15988 9830 16040
rect 9968 16037 9996 16068
rect 10045 16065 10057 16099
rect 10091 16065 10103 16099
rect 10045 16059 10103 16065
rect 10137 16099 10195 16105
rect 10137 16065 10149 16099
rect 10183 16065 10195 16099
rect 10137 16059 10195 16065
rect 10336 16037 10364 16136
rect 11238 16124 11244 16136
rect 11296 16124 11302 16176
rect 16482 16164 16488 16176
rect 15304 16136 16488 16164
rect 13906 16096 13912 16108
rect 10612 16068 13912 16096
rect 9953 16031 10011 16037
rect 9953 15997 9965 16031
rect 9999 15997 10011 16031
rect 9953 15991 10011 15997
rect 10321 16031 10379 16037
rect 10321 15997 10333 16031
rect 10367 15997 10379 16031
rect 10321 15991 10379 15997
rect 6236 15932 7052 15960
rect 8205 15963 8263 15969
rect 6236 15920 6242 15932
rect 8205 15929 8217 15963
rect 8251 15929 8263 15963
rect 8205 15923 8263 15929
rect 2363 15864 5580 15892
rect 5629 15895 5687 15901
rect 2363 15861 2375 15864
rect 2317 15855 2375 15861
rect 5629 15861 5641 15895
rect 5675 15861 5687 15895
rect 5629 15855 5687 15861
rect 6086 15852 6092 15904
rect 6144 15892 6150 15904
rect 8220 15892 8248 15923
rect 6144 15864 8248 15892
rect 8496 15892 8524 15988
rect 8757 15963 8815 15969
rect 8757 15929 8769 15963
rect 8803 15960 8815 15963
rect 10612 15960 10640 16068
rect 13906 16056 13912 16068
rect 13964 16056 13970 16108
rect 10962 16028 10968 16040
rect 10923 16000 10968 16028
rect 10962 15988 10968 16000
rect 11020 15988 11026 16040
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 15997 12035 16031
rect 11977 15991 12035 15997
rect 12437 16031 12495 16037
rect 12437 15997 12449 16031
rect 12483 15997 12495 16031
rect 12437 15991 12495 15997
rect 8803 15932 10640 15960
rect 8803 15929 8815 15932
rect 8757 15923 8815 15929
rect 10686 15920 10692 15972
rect 10744 15960 10750 15972
rect 11992 15960 12020 15991
rect 10744 15932 12020 15960
rect 10744 15920 10750 15932
rect 10505 15895 10563 15901
rect 10505 15892 10517 15895
rect 8496 15864 10517 15892
rect 6144 15852 6150 15864
rect 10505 15861 10517 15864
rect 10551 15861 10563 15895
rect 10505 15855 10563 15861
rect 11238 15852 11244 15904
rect 11296 15892 11302 15904
rect 11793 15895 11851 15901
rect 11793 15892 11805 15895
rect 11296 15864 11805 15892
rect 11296 15852 11302 15864
rect 11793 15861 11805 15864
rect 11839 15861 11851 15895
rect 12452 15892 12480 15991
rect 15194 15988 15200 16040
rect 15252 16028 15258 16040
rect 15304 16028 15332 16136
rect 16316 16105 16344 16136
rect 16482 16124 16488 16136
rect 16540 16124 16546 16176
rect 16301 16099 16359 16105
rect 16301 16065 16313 16099
rect 16347 16065 16359 16099
rect 16301 16059 16359 16065
rect 15473 16031 15531 16037
rect 15473 16028 15485 16031
rect 15252 16000 15485 16028
rect 15252 15988 15258 16000
rect 15473 15997 15485 16000
rect 15519 15997 15531 16031
rect 15473 15991 15531 15997
rect 15657 16031 15715 16037
rect 15657 15997 15669 16031
rect 15703 15997 15715 16031
rect 15657 15991 15715 15997
rect 16209 16031 16267 16037
rect 16209 15997 16221 16031
rect 16255 16028 16267 16031
rect 16574 16028 16580 16040
rect 16255 16000 16580 16028
rect 16255 15997 16267 16000
rect 16209 15991 16267 15997
rect 12710 15960 12716 15972
rect 12671 15932 12716 15960
rect 12710 15920 12716 15932
rect 12768 15920 12774 15972
rect 13446 15920 13452 15972
rect 13504 15920 13510 15972
rect 15010 15920 15016 15972
rect 15068 15960 15074 15972
rect 15105 15963 15163 15969
rect 15105 15960 15117 15963
rect 15068 15932 15117 15960
rect 15068 15920 15074 15932
rect 15105 15929 15117 15932
rect 15151 15929 15163 15963
rect 15672 15960 15700 15991
rect 16224 15960 16252 15991
rect 16574 15988 16580 16000
rect 16632 15988 16638 16040
rect 15672 15932 16252 15960
rect 15105 15923 15163 15929
rect 14366 15892 14372 15904
rect 12452 15864 14372 15892
rect 11793 15855 11851 15861
rect 14366 15852 14372 15864
rect 14424 15852 14430 15904
rect 1104 15802 17296 15824
rect 1104 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 6571 15802
rect 6623 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 11904 15802
rect 11956 15750 11968 15802
rect 12020 15750 17296 15802
rect 1104 15728 17296 15750
rect 1670 15648 1676 15700
rect 1728 15688 1734 15700
rect 1728 15660 4108 15688
rect 1728 15648 1734 15660
rect 2777 15623 2835 15629
rect 2777 15589 2789 15623
rect 2823 15589 2835 15623
rect 4080 15620 4108 15660
rect 4154 15648 4160 15700
rect 4212 15688 4218 15700
rect 5813 15691 5871 15697
rect 5813 15688 5825 15691
rect 4212 15660 5825 15688
rect 4212 15648 4218 15660
rect 5813 15657 5825 15660
rect 5859 15657 5871 15691
rect 5813 15651 5871 15657
rect 5920 15660 7788 15688
rect 5718 15620 5724 15632
rect 4080 15592 5724 15620
rect 2777 15583 2835 15589
rect 1762 15512 1768 15564
rect 1820 15552 1826 15564
rect 1857 15555 1915 15561
rect 1857 15552 1869 15555
rect 1820 15524 1869 15552
rect 1820 15512 1826 15524
rect 1857 15521 1869 15524
rect 1903 15521 1915 15555
rect 1857 15515 1915 15521
rect 2685 15555 2743 15561
rect 2685 15521 2697 15555
rect 2731 15521 2743 15555
rect 2685 15515 2743 15521
rect 2700 15416 2728 15515
rect 2792 15496 2820 15583
rect 5718 15580 5724 15592
rect 5776 15580 5782 15632
rect 5920 15620 5948 15660
rect 6178 15620 6184 15632
rect 5828 15592 5948 15620
rect 6139 15592 6184 15620
rect 2866 15512 2872 15564
rect 2924 15552 2930 15564
rect 3007 15555 3065 15561
rect 2924 15524 2969 15552
rect 2924 15512 2930 15524
rect 3007 15521 3019 15555
rect 3053 15552 3065 15555
rect 3970 15552 3976 15564
rect 3053 15524 3976 15552
rect 3053 15521 3065 15524
rect 3007 15515 3065 15521
rect 3970 15512 3976 15524
rect 4028 15552 4034 15564
rect 4249 15555 4307 15561
rect 4249 15552 4261 15555
rect 4028 15524 4261 15552
rect 4028 15512 4034 15524
rect 4249 15521 4261 15524
rect 4295 15521 4307 15555
rect 4249 15515 4307 15521
rect 5353 15555 5411 15561
rect 5353 15521 5365 15555
rect 5399 15552 5411 15555
rect 5828 15552 5856 15592
rect 6178 15580 6184 15592
rect 6236 15580 6242 15632
rect 5994 15552 6000 15564
rect 5399 15524 5856 15552
rect 5955 15524 6000 15552
rect 5399 15521 5411 15524
rect 5353 15515 5411 15521
rect 5994 15512 6000 15524
rect 6052 15512 6058 15564
rect 6093 15555 6151 15561
rect 6093 15521 6105 15555
rect 6139 15521 6151 15555
rect 6093 15515 6151 15521
rect 6365 15555 6423 15561
rect 6365 15521 6377 15555
rect 6411 15552 6423 15555
rect 6914 15552 6920 15564
rect 6411 15524 6920 15552
rect 6411 15521 6423 15524
rect 6365 15515 6423 15521
rect 2774 15444 2780 15496
rect 2832 15444 2838 15496
rect 3145 15487 3203 15493
rect 3145 15453 3157 15487
rect 3191 15484 3203 15487
rect 3326 15484 3332 15496
rect 3191 15456 3332 15484
rect 3191 15453 3203 15456
rect 3145 15447 3203 15453
rect 3326 15444 3332 15456
rect 3384 15444 3390 15496
rect 6104 15484 6132 15515
rect 6914 15512 6920 15524
rect 6972 15512 6978 15564
rect 7009 15555 7067 15561
rect 7009 15521 7021 15555
rect 7055 15521 7067 15555
rect 7190 15552 7196 15564
rect 7151 15524 7196 15552
rect 7009 15515 7067 15521
rect 6270 15484 6276 15496
rect 6104 15456 6276 15484
rect 6270 15444 6276 15456
rect 6328 15444 6334 15496
rect 7024 15484 7052 15515
rect 7190 15512 7196 15524
rect 7248 15512 7254 15564
rect 7561 15555 7619 15561
rect 7561 15521 7573 15555
rect 7607 15521 7619 15555
rect 7561 15515 7619 15521
rect 7374 15484 7380 15496
rect 6656 15456 7380 15484
rect 2958 15416 2964 15428
rect 2700 15388 2964 15416
rect 2958 15376 2964 15388
rect 3016 15376 3022 15428
rect 6656 15416 6684 15456
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 6196 15388 6684 15416
rect 2041 15351 2099 15357
rect 2041 15317 2053 15351
rect 2087 15348 2099 15351
rect 2130 15348 2136 15360
rect 2087 15320 2136 15348
rect 2087 15317 2099 15320
rect 2041 15311 2099 15317
rect 2130 15308 2136 15320
rect 2188 15308 2194 15360
rect 2222 15308 2228 15360
rect 2280 15348 2286 15360
rect 2501 15351 2559 15357
rect 2501 15348 2513 15351
rect 2280 15320 2513 15348
rect 2280 15308 2286 15320
rect 2501 15317 2513 15320
rect 2547 15317 2559 15351
rect 4338 15348 4344 15360
rect 4299 15320 4344 15348
rect 2501 15311 2559 15317
rect 4338 15308 4344 15320
rect 4396 15308 4402 15360
rect 5261 15351 5319 15357
rect 5261 15317 5273 15351
rect 5307 15348 5319 15351
rect 6196 15348 6224 15388
rect 6730 15376 6736 15428
rect 6788 15416 6794 15428
rect 7576 15416 7604 15515
rect 7760 15493 7788 15660
rect 9766 15648 9772 15700
rect 9824 15688 9830 15700
rect 10410 15688 10416 15700
rect 9824 15660 10416 15688
rect 9824 15648 9830 15660
rect 10410 15648 10416 15660
rect 10468 15648 10474 15700
rect 10594 15648 10600 15700
rect 10652 15688 10658 15700
rect 10870 15688 10876 15700
rect 10652 15660 10876 15688
rect 10652 15648 10658 15660
rect 10870 15648 10876 15660
rect 10928 15688 10934 15700
rect 12710 15688 12716 15700
rect 10928 15660 12020 15688
rect 12671 15660 12716 15688
rect 10928 15648 10934 15660
rect 9950 15580 9956 15632
rect 10008 15620 10014 15632
rect 10045 15623 10103 15629
rect 10045 15620 10057 15623
rect 10008 15592 10057 15620
rect 10008 15580 10014 15592
rect 10045 15589 10057 15592
rect 10091 15589 10103 15623
rect 10226 15620 10232 15632
rect 10187 15592 10232 15620
rect 10045 15583 10103 15589
rect 10226 15580 10232 15592
rect 10284 15580 10290 15632
rect 11606 15620 11612 15632
rect 10336 15592 11612 15620
rect 7929 15555 7987 15561
rect 7929 15521 7941 15555
rect 7975 15552 7987 15555
rect 7975 15524 8248 15552
rect 7975 15521 7987 15524
rect 7929 15515 7987 15521
rect 7745 15487 7803 15493
rect 7745 15453 7757 15487
rect 7791 15453 7803 15487
rect 7745 15447 7803 15453
rect 8021 15487 8079 15493
rect 8021 15453 8033 15487
rect 8067 15484 8079 15487
rect 8110 15484 8116 15496
rect 8067 15456 8116 15484
rect 8067 15453 8079 15456
rect 8021 15447 8079 15453
rect 6788 15388 7604 15416
rect 7760 15416 7788 15447
rect 8110 15444 8116 15456
rect 8168 15444 8174 15496
rect 8220 15484 8248 15524
rect 8294 15512 8300 15564
rect 8352 15552 8358 15564
rect 10336 15552 10364 15592
rect 11606 15580 11612 15592
rect 11664 15580 11670 15632
rect 11992 15561 12020 15660
rect 12710 15648 12716 15660
rect 12768 15648 12774 15700
rect 16574 15688 16580 15700
rect 16535 15660 16580 15688
rect 16574 15648 16580 15660
rect 16632 15648 16638 15700
rect 13078 15620 13084 15632
rect 12268 15592 13084 15620
rect 8352 15524 10364 15552
rect 11149 15555 11207 15561
rect 8352 15512 8358 15524
rect 11149 15521 11161 15555
rect 11195 15521 11207 15555
rect 11149 15515 11207 15521
rect 11977 15555 12035 15561
rect 11977 15521 11989 15555
rect 12023 15521 12035 15555
rect 12158 15552 12164 15564
rect 12119 15524 12164 15552
rect 11977 15515 12035 15521
rect 8662 15484 8668 15496
rect 8220 15456 8668 15484
rect 8662 15444 8668 15456
rect 8720 15484 8726 15496
rect 10873 15487 10931 15493
rect 10873 15484 10885 15487
rect 8720 15456 10885 15484
rect 8720 15444 8726 15456
rect 10873 15453 10885 15456
rect 10919 15453 10931 15487
rect 10873 15447 10931 15453
rect 8754 15416 8760 15428
rect 7760 15388 8760 15416
rect 6788 15376 6794 15388
rect 8754 15376 8760 15388
rect 8812 15376 8818 15428
rect 9674 15376 9680 15428
rect 9732 15416 9738 15428
rect 10965 15419 11023 15425
rect 10965 15416 10977 15419
rect 9732 15388 10977 15416
rect 9732 15376 9738 15388
rect 10965 15385 10977 15388
rect 11011 15385 11023 15419
rect 11164 15416 11192 15515
rect 12158 15512 12164 15524
rect 12216 15512 12222 15564
rect 12268 15561 12296 15592
rect 13078 15580 13084 15592
rect 13136 15580 13142 15632
rect 15105 15623 15163 15629
rect 15105 15589 15117 15623
rect 15151 15620 15163 15623
rect 15194 15620 15200 15632
rect 15151 15592 15200 15620
rect 15151 15589 15163 15592
rect 15105 15583 15163 15589
rect 15194 15580 15200 15592
rect 15252 15580 15258 15632
rect 15562 15580 15568 15632
rect 15620 15580 15626 15632
rect 12253 15555 12311 15561
rect 12253 15521 12265 15555
rect 12299 15521 12311 15555
rect 12253 15515 12311 15521
rect 12345 15555 12403 15561
rect 12345 15521 12357 15555
rect 12391 15552 12403 15555
rect 12434 15552 12440 15564
rect 12391 15524 12440 15552
rect 12391 15521 12403 15524
rect 12345 15515 12403 15521
rect 12434 15512 12440 15524
rect 12492 15512 12498 15564
rect 12529 15555 12587 15561
rect 12529 15521 12541 15555
rect 12575 15552 12587 15555
rect 13170 15552 13176 15564
rect 12575 15524 13176 15552
rect 12575 15521 12587 15524
rect 12529 15515 12587 15521
rect 13170 15512 13176 15524
rect 13228 15512 13234 15564
rect 13262 15512 13268 15564
rect 13320 15552 13326 15564
rect 13814 15552 13820 15564
rect 13320 15524 13820 15552
rect 13320 15512 13326 15524
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 12176 15484 12204 15512
rect 13078 15484 13084 15496
rect 12176 15456 13084 15484
rect 13078 15444 13084 15456
rect 13136 15444 13142 15496
rect 14366 15444 14372 15496
rect 14424 15484 14430 15496
rect 14829 15487 14887 15493
rect 14829 15484 14841 15487
rect 14424 15456 14841 15484
rect 14424 15444 14430 15456
rect 14829 15453 14841 15456
rect 14875 15453 14887 15487
rect 14829 15447 14887 15453
rect 13725 15419 13783 15425
rect 13725 15416 13737 15419
rect 11164 15388 13737 15416
rect 10965 15379 11023 15385
rect 13725 15385 13737 15388
rect 13771 15385 13783 15419
rect 13725 15379 13783 15385
rect 5307 15320 6224 15348
rect 5307 15317 5319 15320
rect 5261 15311 5319 15317
rect 6270 15308 6276 15360
rect 6328 15348 6334 15360
rect 10686 15348 10692 15360
rect 6328 15320 10692 15348
rect 6328 15308 6334 15320
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 11057 15351 11115 15357
rect 11057 15317 11069 15351
rect 11103 15348 11115 15351
rect 13630 15348 13636 15360
rect 11103 15320 13636 15348
rect 11103 15317 11115 15320
rect 11057 15311 11115 15317
rect 13630 15308 13636 15320
rect 13688 15308 13694 15360
rect 1104 15258 17296 15280
rect 1104 15206 3680 15258
rect 3732 15206 3744 15258
rect 3796 15206 3808 15258
rect 3860 15206 3872 15258
rect 3924 15206 9078 15258
rect 9130 15206 9142 15258
rect 9194 15206 9206 15258
rect 9258 15206 9270 15258
rect 9322 15206 14475 15258
rect 14527 15206 14539 15258
rect 14591 15206 14603 15258
rect 14655 15206 14667 15258
rect 14719 15206 17296 15258
rect 1104 15184 17296 15206
rect 4065 15147 4123 15153
rect 4065 15113 4077 15147
rect 4111 15144 4123 15147
rect 5813 15147 5871 15153
rect 4111 15116 4844 15144
rect 4111 15113 4123 15116
rect 4065 15107 4123 15113
rect 2774 15036 2780 15088
rect 2832 15076 2838 15088
rect 2832 15048 4660 15076
rect 2832 15036 2838 15048
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 2222 15008 2228 15020
rect 1719 14980 2228 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 2222 14968 2228 14980
rect 2280 14968 2286 15020
rect 3145 15011 3203 15017
rect 3145 14977 3157 15011
rect 3191 15008 3203 15011
rect 3970 15008 3976 15020
rect 3191 14980 3976 15008
rect 3191 14977 3203 14980
rect 3145 14971 3203 14977
rect 1394 14940 1400 14952
rect 1355 14912 1400 14940
rect 1394 14900 1400 14912
rect 1452 14900 1458 14952
rect 3804 14949 3832 14980
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 4632 15017 4660 15048
rect 4816 15017 4844 15116
rect 5813 15113 5825 15147
rect 5859 15144 5871 15147
rect 7190 15144 7196 15156
rect 5859 15116 7196 15144
rect 5859 15113 5871 15116
rect 5813 15107 5871 15113
rect 7190 15104 7196 15116
rect 7248 15104 7254 15156
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 10137 15147 10195 15153
rect 10137 15144 10149 15147
rect 10008 15116 10149 15144
rect 10008 15104 10014 15116
rect 10137 15113 10149 15116
rect 10183 15113 10195 15147
rect 10137 15107 10195 15113
rect 13081 15147 13139 15153
rect 13081 15113 13093 15147
rect 13127 15144 13139 15147
rect 13262 15144 13268 15156
rect 13127 15116 13268 15144
rect 13127 15113 13139 15116
rect 13081 15107 13139 15113
rect 13262 15104 13268 15116
rect 13320 15104 13326 15156
rect 14918 15144 14924 15156
rect 13464 15116 14924 15144
rect 7282 15036 7288 15088
rect 7340 15076 7346 15088
rect 10962 15076 10968 15088
rect 7340 15048 10968 15076
rect 7340 15036 7346 15048
rect 4617 15011 4675 15017
rect 4617 14977 4629 15011
rect 4663 14977 4675 15011
rect 4617 14971 4675 14977
rect 4801 15011 4859 15017
rect 4801 14977 4813 15011
rect 4847 15008 4859 15011
rect 5166 15008 5172 15020
rect 4847 14980 5172 15008
rect 4847 14977 4859 14980
rect 4801 14971 4859 14977
rect 5166 14968 5172 14980
rect 5224 14968 5230 15020
rect 7392 15017 7420 15048
rect 10962 15036 10968 15048
rect 11020 15036 11026 15088
rect 11054 15036 11060 15088
rect 11112 15076 11118 15088
rect 13464 15076 13492 15116
rect 14918 15104 14924 15116
rect 14976 15104 14982 15156
rect 11112 15048 13032 15076
rect 11112 15036 11118 15048
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 14977 7435 15011
rect 9766 15008 9772 15020
rect 7377 14971 7435 14977
rect 8588 14980 9772 15008
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14909 3847 14943
rect 3789 14903 3847 14909
rect 3881 14943 3939 14949
rect 3881 14909 3893 14943
rect 3927 14909 3939 14943
rect 3881 14903 3939 14909
rect 4157 14943 4215 14949
rect 4157 14909 4169 14943
rect 4203 14940 4215 14943
rect 4338 14940 4344 14952
rect 4203 14912 4344 14940
rect 4203 14909 4215 14912
rect 4157 14903 4215 14909
rect 2130 14832 2136 14884
rect 2188 14832 2194 14884
rect 3896 14872 3924 14903
rect 4338 14900 4344 14912
rect 4396 14900 4402 14952
rect 4893 14943 4951 14949
rect 4893 14909 4905 14943
rect 4939 14909 4951 14943
rect 4893 14903 4951 14909
rect 4356 14872 4384 14900
rect 4908 14872 4936 14903
rect 5626 14900 5632 14952
rect 5684 14940 5690 14952
rect 5721 14943 5779 14949
rect 5721 14940 5733 14943
rect 5684 14912 5733 14940
rect 5684 14900 5690 14912
rect 5721 14909 5733 14912
rect 5767 14940 5779 14943
rect 6730 14940 6736 14952
rect 5767 14912 6736 14940
rect 5767 14909 5779 14912
rect 5721 14903 5779 14909
rect 6730 14900 6736 14912
rect 6788 14900 6794 14952
rect 6914 14940 6920 14952
rect 6875 14912 6920 14940
rect 6914 14900 6920 14912
rect 6972 14900 6978 14952
rect 8386 14940 8392 14952
rect 8347 14912 8392 14940
rect 8386 14900 8392 14912
rect 8444 14900 8450 14952
rect 8588 14949 8616 14980
rect 9766 14968 9772 14980
rect 9824 14968 9830 15020
rect 9950 14968 9956 15020
rect 10008 15008 10014 15020
rect 10781 15011 10839 15017
rect 10781 15008 10793 15011
rect 10008 14980 10793 15008
rect 10008 14968 10014 14980
rect 10781 14977 10793 14980
rect 10827 15008 10839 15011
rect 12161 15011 12219 15017
rect 12161 15008 12173 15011
rect 10827 14980 12173 15008
rect 10827 14977 10839 14980
rect 10781 14971 10839 14977
rect 12161 14977 12173 14980
rect 12207 14977 12219 15011
rect 12161 14971 12219 14977
rect 8573 14943 8631 14949
rect 8573 14909 8585 14943
rect 8619 14909 8631 14943
rect 8754 14940 8760 14952
rect 8715 14912 8760 14940
rect 8573 14903 8631 14909
rect 8754 14900 8760 14912
rect 8812 14900 8818 14952
rect 8941 14943 8999 14949
rect 8941 14909 8953 14943
rect 8987 14909 8999 14943
rect 8941 14903 8999 14909
rect 9309 14943 9367 14949
rect 9309 14909 9321 14943
rect 9355 14940 9367 14943
rect 9674 14940 9680 14952
rect 9355 14912 9680 14940
rect 9355 14909 9367 14912
rect 9309 14903 9367 14909
rect 7926 14872 7932 14884
rect 3896 14844 4200 14872
rect 4356 14844 4936 14872
rect 7887 14844 7932 14872
rect 4172 14816 4200 14844
rect 7926 14832 7932 14844
rect 7984 14832 7990 14884
rect 8018 14832 8024 14884
rect 8076 14872 8082 14884
rect 8956 14872 8984 14903
rect 9674 14900 9680 14912
rect 9732 14900 9738 14952
rect 10318 14940 10324 14952
rect 10279 14912 10324 14940
rect 10318 14900 10324 14912
rect 10376 14900 10382 14952
rect 10686 14940 10692 14952
rect 10647 14912 10692 14940
rect 10686 14900 10692 14912
rect 10744 14900 10750 14952
rect 12069 14943 12127 14949
rect 12069 14909 12081 14943
rect 12115 14909 12127 14943
rect 12069 14903 12127 14909
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 12618 14940 12624 14952
rect 12299 14912 12624 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12084 14872 12112 14903
rect 12618 14900 12624 14912
rect 12676 14940 12682 14952
rect 13004 14949 13032 15048
rect 13372 15048 13492 15076
rect 13372 15008 13400 15048
rect 13814 15036 13820 15088
rect 13872 15076 13878 15088
rect 13872 15048 15332 15076
rect 13872 15036 13878 15048
rect 13630 15008 13636 15020
rect 13188 14980 13400 15008
rect 13591 14980 13636 15008
rect 13188 14949 13216 14980
rect 13630 14968 13636 14980
rect 13688 15008 13694 15020
rect 14553 15011 14611 15017
rect 14553 15008 14565 15011
rect 13688 14980 14565 15008
rect 13688 14968 13694 14980
rect 14553 14977 14565 14980
rect 14599 14977 14611 15011
rect 14553 14971 14611 14977
rect 14660 14980 15056 15008
rect 12989 14943 13047 14949
rect 12676 14912 12848 14940
rect 12676 14900 12682 14912
rect 12434 14872 12440 14884
rect 8076 14844 8984 14872
rect 10336 14844 12440 14872
rect 8076 14832 8082 14844
rect 3326 14764 3332 14816
rect 3384 14804 3390 14816
rect 3605 14807 3663 14813
rect 3605 14804 3617 14807
rect 3384 14776 3617 14804
rect 3384 14764 3390 14776
rect 3605 14773 3617 14776
rect 3651 14773 3663 14807
rect 3605 14767 3663 14773
rect 4154 14764 4160 14816
rect 4212 14764 4218 14816
rect 4617 14807 4675 14813
rect 4617 14773 4629 14807
rect 4663 14804 4675 14807
rect 5074 14804 5080 14816
rect 4663 14776 5080 14804
rect 4663 14773 4675 14776
rect 4617 14767 4675 14773
rect 5074 14764 5080 14776
rect 5132 14764 5138 14816
rect 10226 14764 10232 14816
rect 10284 14804 10290 14816
rect 10336 14813 10364 14844
rect 12434 14832 12440 14844
rect 12492 14832 12498 14884
rect 10321 14807 10379 14813
rect 10321 14804 10333 14807
rect 10284 14776 10333 14804
rect 10284 14764 10290 14776
rect 10321 14773 10333 14776
rect 10367 14773 10379 14807
rect 12820 14804 12848 14912
rect 12989 14909 13001 14943
rect 13035 14909 13047 14943
rect 12989 14903 13047 14909
rect 13173 14943 13231 14949
rect 13173 14909 13185 14943
rect 13219 14909 13231 14943
rect 13173 14903 13231 14909
rect 13817 14943 13875 14949
rect 13817 14909 13829 14943
rect 13863 14940 13875 14943
rect 13906 14940 13912 14952
rect 13863 14912 13912 14940
rect 13863 14909 13875 14912
rect 13817 14903 13875 14909
rect 13004 14872 13032 14903
rect 13906 14900 13912 14912
rect 13964 14900 13970 14952
rect 14093 14943 14151 14949
rect 14093 14909 14105 14943
rect 14139 14940 14151 14943
rect 14660 14940 14688 14980
rect 14139 14912 14688 14940
rect 14737 14943 14795 14949
rect 14139 14909 14151 14912
rect 14093 14903 14151 14909
rect 14737 14909 14749 14943
rect 14783 14909 14795 14943
rect 14918 14940 14924 14952
rect 14879 14912 14924 14940
rect 14737 14903 14795 14909
rect 14752 14872 14780 14903
rect 14918 14900 14924 14912
rect 14976 14900 14982 14952
rect 15028 14949 15056 14980
rect 15013 14943 15071 14949
rect 15013 14909 15025 14943
rect 15059 14909 15071 14943
rect 15013 14903 15071 14909
rect 13004 14844 14780 14872
rect 15028 14872 15056 14903
rect 15102 14900 15108 14952
rect 15160 14940 15166 14952
rect 15304 14949 15332 15048
rect 15289 14943 15347 14949
rect 15160 14912 15205 14940
rect 15160 14900 15166 14912
rect 15289 14909 15301 14943
rect 15335 14909 15347 14943
rect 15289 14903 15347 14909
rect 15749 14943 15807 14949
rect 15749 14909 15761 14943
rect 15795 14940 15807 14943
rect 15930 14940 15936 14952
rect 15795 14912 15936 14940
rect 15795 14909 15807 14912
rect 15749 14903 15807 14909
rect 15930 14900 15936 14912
rect 15988 14900 15994 14952
rect 16206 14872 16212 14884
rect 15028 14844 16212 14872
rect 16206 14832 16212 14844
rect 16264 14832 16270 14884
rect 13170 14804 13176 14816
rect 12820 14776 13176 14804
rect 10321 14767 10379 14773
rect 13170 14764 13176 14776
rect 13228 14764 13234 14816
rect 14001 14807 14059 14813
rect 14001 14773 14013 14807
rect 14047 14804 14059 14807
rect 15102 14804 15108 14816
rect 14047 14776 15108 14804
rect 14047 14773 14059 14776
rect 14001 14767 14059 14773
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 15838 14804 15844 14816
rect 15799 14776 15844 14804
rect 15838 14764 15844 14776
rect 15896 14764 15902 14816
rect 1104 14714 17296 14736
rect 1104 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 6571 14714
rect 6623 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 11904 14714
rect 11956 14662 11968 14714
rect 12020 14662 17296 14714
rect 1104 14640 17296 14662
rect 2501 14603 2559 14609
rect 2501 14569 2513 14603
rect 2547 14600 2559 14603
rect 2774 14600 2780 14612
rect 2547 14572 2780 14600
rect 2547 14569 2559 14572
rect 2501 14563 2559 14569
rect 2774 14560 2780 14572
rect 2832 14560 2838 14612
rect 2958 14600 2964 14612
rect 2919 14572 2964 14600
rect 2958 14560 2964 14572
rect 3016 14560 3022 14612
rect 7745 14603 7803 14609
rect 3896 14572 6592 14600
rect 3326 14532 3332 14544
rect 2332 14504 3332 14532
rect 1673 14467 1731 14473
rect 1673 14433 1685 14467
rect 1719 14464 1731 14467
rect 1762 14464 1768 14476
rect 1719 14436 1768 14464
rect 1719 14433 1731 14436
rect 1673 14427 1731 14433
rect 1762 14424 1768 14436
rect 1820 14424 1826 14476
rect 2332 14473 2360 14504
rect 3326 14492 3332 14504
rect 3384 14492 3390 14544
rect 2317 14467 2375 14473
rect 2317 14433 2329 14467
rect 2363 14433 2375 14467
rect 2317 14427 2375 14433
rect 2501 14467 2559 14473
rect 2501 14433 2513 14467
rect 2547 14464 2559 14467
rect 3050 14464 3056 14476
rect 2547 14436 3056 14464
rect 2547 14433 2559 14436
rect 2501 14427 2559 14433
rect 3050 14424 3056 14436
rect 3108 14464 3114 14476
rect 3145 14467 3203 14473
rect 3145 14464 3157 14467
rect 3108 14436 3157 14464
rect 3108 14424 3114 14436
rect 3145 14433 3157 14436
rect 3191 14433 3203 14467
rect 3145 14427 3203 14433
rect 1946 14356 1952 14408
rect 2004 14396 2010 14408
rect 3896 14396 3924 14572
rect 6564 14532 6592 14572
rect 7745 14569 7757 14603
rect 7791 14600 7803 14603
rect 8018 14600 8024 14612
rect 7791 14572 8024 14600
rect 7791 14569 7803 14572
rect 7745 14563 7803 14569
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 8573 14603 8631 14609
rect 8573 14569 8585 14603
rect 8619 14600 8631 14603
rect 8754 14600 8760 14612
rect 8619 14572 8760 14600
rect 8619 14569 8631 14572
rect 8573 14563 8631 14569
rect 8754 14560 8760 14572
rect 8812 14560 8818 14612
rect 10137 14603 10195 14609
rect 10137 14569 10149 14603
rect 10183 14600 10195 14603
rect 10318 14600 10324 14612
rect 10183 14572 10324 14600
rect 10183 14569 10195 14572
rect 10137 14563 10195 14569
rect 10318 14560 10324 14572
rect 10376 14600 10382 14612
rect 10376 14572 12296 14600
rect 10376 14560 10382 14572
rect 8386 14532 8392 14544
rect 2004 14368 3924 14396
rect 3988 14504 5290 14532
rect 6564 14504 8392 14532
rect 2004 14356 2010 14368
rect 1857 14331 1915 14337
rect 1857 14297 1869 14331
rect 1903 14328 1915 14331
rect 3988 14328 4016 14504
rect 8386 14492 8392 14504
rect 8444 14492 8450 14544
rect 10962 14532 10968 14544
rect 10923 14504 10968 14532
rect 10962 14492 10968 14504
rect 11020 14492 11026 14544
rect 7377 14467 7435 14473
rect 7377 14433 7389 14467
rect 7423 14464 7435 14467
rect 8018 14464 8024 14476
rect 7423 14436 8024 14464
rect 7423 14433 7435 14436
rect 7377 14427 7435 14433
rect 8018 14424 8024 14436
rect 8076 14424 8082 14476
rect 8202 14464 8208 14476
rect 8163 14436 8208 14464
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 9950 14464 9956 14476
rect 9911 14436 9956 14464
rect 9950 14424 9956 14436
rect 10008 14424 10014 14476
rect 10226 14464 10232 14476
rect 10187 14436 10232 14464
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 12268 14464 12296 14572
rect 12434 14560 12440 14612
rect 12492 14600 12498 14612
rect 12492 14572 12537 14600
rect 12492 14560 12498 14572
rect 13170 14560 13176 14612
rect 13228 14600 13234 14612
rect 13228 14572 13308 14600
rect 13228 14560 13234 14572
rect 12526 14492 12532 14544
rect 12584 14532 12590 14544
rect 13280 14541 13308 14572
rect 15930 14560 15936 14612
rect 15988 14560 15994 14612
rect 16206 14560 16212 14612
rect 16264 14600 16270 14612
rect 16393 14603 16451 14609
rect 16393 14600 16405 14603
rect 16264 14572 16405 14600
rect 16264 14560 16270 14572
rect 16393 14569 16405 14572
rect 16439 14569 16451 14603
rect 16393 14563 16451 14569
rect 13265 14535 13323 14541
rect 12584 14504 13216 14532
rect 12584 14492 12590 14504
rect 13188 14476 13216 14504
rect 13265 14501 13277 14535
rect 13311 14501 13323 14535
rect 14826 14532 14832 14544
rect 13265 14495 13323 14501
rect 13464 14504 14832 14532
rect 12434 14464 12440 14476
rect 4246 14356 4252 14408
rect 4304 14396 4310 14408
rect 4525 14399 4583 14405
rect 4525 14396 4537 14399
rect 4304 14368 4537 14396
rect 4304 14356 4310 14368
rect 4525 14365 4537 14368
rect 4571 14365 4583 14399
rect 4525 14359 4583 14365
rect 4801 14399 4859 14405
rect 4801 14365 4813 14399
rect 4847 14396 4859 14399
rect 5258 14396 5264 14408
rect 4847 14368 5264 14396
rect 4847 14365 4859 14368
rect 4801 14359 4859 14365
rect 1903 14300 4016 14328
rect 1903 14297 1915 14300
rect 1857 14291 1915 14297
rect 4540 14260 4568 14359
rect 5258 14356 5264 14368
rect 5316 14356 5322 14408
rect 7190 14356 7196 14408
rect 7248 14396 7254 14408
rect 7469 14399 7527 14405
rect 7469 14396 7481 14399
rect 7248 14368 7481 14396
rect 7248 14356 7254 14368
rect 7469 14365 7481 14368
rect 7515 14365 7527 14399
rect 7469 14359 7527 14365
rect 8478 14356 8484 14408
rect 8536 14396 8542 14408
rect 9858 14396 9864 14408
rect 8536 14368 9864 14396
rect 8536 14356 8542 14368
rect 9858 14356 9864 14368
rect 9916 14396 9922 14408
rect 10689 14399 10747 14405
rect 10689 14396 10701 14399
rect 9916 14368 10701 14396
rect 9916 14356 9922 14368
rect 10689 14365 10701 14368
rect 10735 14396 10747 14399
rect 11330 14396 11336 14408
rect 10735 14368 11336 14396
rect 10735 14365 10747 14368
rect 10689 14359 10747 14365
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 12084 14396 12112 14450
rect 12268 14436 12440 14464
rect 12434 14424 12440 14436
rect 12492 14464 12498 14476
rect 12618 14464 12624 14476
rect 12492 14436 12624 14464
rect 12492 14424 12498 14436
rect 12618 14424 12624 14436
rect 12676 14424 12682 14476
rect 13078 14464 13084 14476
rect 13039 14436 13084 14464
rect 13078 14424 13084 14436
rect 13136 14424 13142 14476
rect 13170 14424 13176 14476
rect 13228 14464 13234 14476
rect 13464 14473 13492 14504
rect 14826 14492 14832 14504
rect 14884 14492 14890 14544
rect 15197 14535 15255 14541
rect 15197 14501 15209 14535
rect 15243 14532 15255 14535
rect 15948 14532 15976 14560
rect 15243 14504 15976 14532
rect 15243 14501 15255 14504
rect 15197 14495 15255 14501
rect 13449 14467 13507 14473
rect 13228 14436 13273 14464
rect 13228 14424 13234 14436
rect 13449 14433 13461 14467
rect 13495 14433 13507 14467
rect 13449 14427 13507 14433
rect 13541 14467 13599 14473
rect 13541 14433 13553 14467
rect 13587 14433 13599 14467
rect 13541 14427 13599 14433
rect 12342 14396 12348 14408
rect 12084 14368 12348 14396
rect 12342 14356 12348 14368
rect 12400 14356 12406 14408
rect 8496 14328 8524 14356
rect 13556 14328 13584 14427
rect 14274 14424 14280 14476
rect 14332 14464 14338 14476
rect 15010 14464 15016 14476
rect 14332 14436 15016 14464
rect 14332 14424 14338 14436
rect 15010 14424 15016 14436
rect 15068 14464 15074 14476
rect 15105 14467 15163 14473
rect 15105 14464 15117 14467
rect 15068 14436 15117 14464
rect 15068 14424 15074 14436
rect 15105 14433 15117 14436
rect 15151 14433 15163 14467
rect 15105 14427 15163 14433
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 15473 14467 15531 14473
rect 15473 14433 15485 14467
rect 15519 14464 15531 14467
rect 15654 14464 15660 14476
rect 15519 14436 15660 14464
rect 15519 14433 15531 14436
rect 15473 14427 15531 14433
rect 14090 14356 14096 14408
rect 14148 14396 14154 14408
rect 15304 14396 15332 14427
rect 14148 14368 15332 14396
rect 14148 14356 14154 14368
rect 14734 14328 14740 14340
rect 5828 14300 8524 14328
rect 12406 14300 14740 14328
rect 4982 14260 4988 14272
rect 4540 14232 4988 14260
rect 4982 14220 4988 14232
rect 5040 14260 5046 14272
rect 5828 14260 5856 14300
rect 5040 14232 5856 14260
rect 5040 14220 5046 14232
rect 6086 14220 6092 14272
rect 6144 14260 6150 14272
rect 6273 14263 6331 14269
rect 6273 14260 6285 14263
rect 6144 14232 6285 14260
rect 6144 14220 6150 14232
rect 6273 14229 6285 14232
rect 6319 14229 6331 14263
rect 7374 14260 7380 14272
rect 7335 14232 7380 14260
rect 6273 14223 6331 14229
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 9766 14260 9772 14272
rect 9727 14232 9772 14260
rect 9766 14220 9772 14232
rect 9824 14220 9830 14272
rect 11146 14220 11152 14272
rect 11204 14260 11210 14272
rect 12406 14260 12434 14300
rect 14734 14288 14740 14300
rect 14792 14328 14798 14340
rect 15488 14328 15516 14427
rect 15654 14424 15660 14436
rect 15712 14424 15718 14476
rect 15838 14424 15844 14476
rect 15896 14464 15902 14476
rect 15933 14467 15991 14473
rect 15933 14464 15945 14467
rect 15896 14436 15945 14464
rect 15896 14424 15902 14436
rect 15933 14433 15945 14436
rect 15979 14433 15991 14467
rect 15933 14427 15991 14433
rect 16025 14467 16083 14473
rect 16025 14433 16037 14467
rect 16071 14464 16083 14467
rect 16209 14467 16267 14473
rect 16071 14436 16160 14464
rect 16071 14433 16083 14436
rect 16025 14427 16083 14433
rect 16132 14396 16160 14436
rect 16209 14433 16221 14467
rect 16255 14464 16267 14467
rect 16298 14464 16304 14476
rect 16255 14436 16304 14464
rect 16255 14433 16267 14436
rect 16209 14427 16267 14433
rect 16298 14424 16304 14436
rect 16356 14424 16362 14476
rect 16482 14396 16488 14408
rect 16132 14368 16488 14396
rect 16482 14356 16488 14368
rect 16540 14356 16546 14408
rect 14792 14300 15516 14328
rect 14792 14288 14798 14300
rect 11204 14232 12434 14260
rect 11204 14220 11210 14232
rect 12618 14220 12624 14272
rect 12676 14260 12682 14272
rect 12897 14263 12955 14269
rect 12897 14260 12909 14263
rect 12676 14232 12909 14260
rect 12676 14220 12682 14232
rect 12897 14229 12909 14232
rect 12943 14229 12955 14263
rect 14918 14260 14924 14272
rect 14879 14232 14924 14260
rect 12897 14223 12955 14229
rect 14918 14220 14924 14232
rect 14976 14220 14982 14272
rect 1104 14170 17296 14192
rect 1104 14118 3680 14170
rect 3732 14118 3744 14170
rect 3796 14118 3808 14170
rect 3860 14118 3872 14170
rect 3924 14118 9078 14170
rect 9130 14118 9142 14170
rect 9194 14118 9206 14170
rect 9258 14118 9270 14170
rect 9322 14118 14475 14170
rect 14527 14118 14539 14170
rect 14591 14118 14603 14170
rect 14655 14118 14667 14170
rect 14719 14118 17296 14170
rect 1104 14096 17296 14118
rect 3234 14056 3240 14068
rect 1872 14028 3240 14056
rect 1872 13861 1900 14028
rect 3234 14016 3240 14028
rect 3292 14016 3298 14068
rect 5074 14056 5080 14068
rect 3344 14028 5080 14056
rect 2041 13991 2099 13997
rect 2041 13957 2053 13991
rect 2087 13988 2099 13991
rect 2590 13988 2596 14000
rect 2087 13960 2596 13988
rect 2087 13957 2099 13960
rect 2041 13951 2099 13957
rect 2590 13948 2596 13960
rect 2648 13948 2654 14000
rect 1857 13855 1915 13861
rect 1857 13821 1869 13855
rect 1903 13821 1915 13855
rect 1857 13815 1915 13821
rect 2685 13855 2743 13861
rect 2685 13821 2697 13855
rect 2731 13852 2743 13855
rect 3344 13852 3372 14028
rect 5074 14016 5080 14028
rect 5132 14016 5138 14068
rect 5258 14056 5264 14068
rect 5219 14028 5264 14056
rect 5258 14016 5264 14028
rect 5316 14016 5322 14068
rect 6730 14016 6736 14068
rect 6788 14056 6794 14068
rect 6917 14059 6975 14065
rect 6917 14056 6929 14059
rect 6788 14028 6929 14056
rect 6788 14016 6794 14028
rect 6917 14025 6929 14028
rect 6963 14056 6975 14059
rect 7926 14056 7932 14068
rect 6963 14028 7932 14056
rect 6963 14025 6975 14028
rect 6917 14019 6975 14025
rect 7926 14016 7932 14028
rect 7984 14016 7990 14068
rect 8110 14056 8116 14068
rect 8071 14028 8116 14056
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 9953 14059 10011 14065
rect 9953 14056 9965 14059
rect 9824 14028 9965 14056
rect 9824 14016 9830 14028
rect 9953 14025 9965 14028
rect 9999 14025 10011 14059
rect 9953 14019 10011 14025
rect 10962 14016 10968 14068
rect 11020 14056 11026 14068
rect 11149 14059 11207 14065
rect 11149 14056 11161 14059
rect 11020 14028 11161 14056
rect 11020 14016 11026 14028
rect 11149 14025 11161 14028
rect 11195 14025 11207 14059
rect 14090 14056 14096 14068
rect 14051 14028 14096 14056
rect 11149 14019 11207 14025
rect 14090 14016 14096 14028
rect 14148 14016 14154 14068
rect 15930 14016 15936 14068
rect 15988 14056 15994 14068
rect 16393 14059 16451 14065
rect 16393 14056 16405 14059
rect 15988 14028 16405 14056
rect 15988 14016 15994 14028
rect 16393 14025 16405 14028
rect 16439 14025 16451 14059
rect 16393 14019 16451 14025
rect 3789 13991 3847 13997
rect 3789 13957 3801 13991
rect 3835 13988 3847 13991
rect 4338 13988 4344 14000
rect 3835 13960 4344 13988
rect 3835 13957 3847 13960
rect 3789 13951 3847 13957
rect 4338 13948 4344 13960
rect 4396 13948 4402 14000
rect 5169 13991 5227 13997
rect 5169 13957 5181 13991
rect 5215 13988 5227 13991
rect 5902 13988 5908 14000
rect 5215 13960 5908 13988
rect 5215 13957 5227 13960
rect 5169 13951 5227 13957
rect 5902 13948 5908 13960
rect 5960 13948 5966 14000
rect 8202 13948 8208 14000
rect 8260 13988 8266 14000
rect 9401 13991 9459 13997
rect 9401 13988 9413 13991
rect 8260 13960 9413 13988
rect 8260 13948 8266 13960
rect 3970 13880 3976 13932
rect 4028 13920 4034 13932
rect 7101 13923 7159 13929
rect 7101 13920 7113 13923
rect 4028 13892 5488 13920
rect 4028 13880 4034 13892
rect 3510 13852 3516 13864
rect 2731 13824 3372 13852
rect 3471 13824 3516 13852
rect 2731 13821 2743 13824
rect 2685 13815 2743 13821
rect 3510 13812 3516 13824
rect 3568 13812 3574 13864
rect 3605 13855 3663 13861
rect 3605 13821 3617 13855
rect 3651 13852 3663 13855
rect 3881 13855 3939 13861
rect 3651 13824 3832 13852
rect 3651 13821 3663 13824
rect 3605 13815 3663 13821
rect 2869 13787 2927 13793
rect 2869 13753 2881 13787
rect 2915 13753 2927 13787
rect 2869 13747 2927 13753
rect 2501 13719 2559 13725
rect 2501 13685 2513 13719
rect 2547 13716 2559 13719
rect 2774 13716 2780 13728
rect 2547 13688 2780 13716
rect 2547 13685 2559 13688
rect 2501 13679 2559 13685
rect 2774 13676 2780 13688
rect 2832 13676 2838 13728
rect 2884 13716 2912 13747
rect 2958 13744 2964 13796
rect 3016 13784 3022 13796
rect 3804 13784 3832 13824
rect 3881 13821 3893 13855
rect 3927 13852 3939 13855
rect 4062 13852 4068 13864
rect 3927 13824 4068 13852
rect 3927 13821 3939 13824
rect 3881 13815 3939 13821
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 4338 13852 4344 13864
rect 4299 13824 4344 13852
rect 4338 13812 4344 13824
rect 4396 13812 4402 13864
rect 5460 13861 5488 13892
rect 6748 13892 7113 13920
rect 5169 13855 5227 13861
rect 5169 13852 5181 13855
rect 4632 13824 5181 13852
rect 4154 13784 4160 13796
rect 3016 13756 3464 13784
rect 3804 13756 4160 13784
rect 3016 13744 3022 13756
rect 3326 13716 3332 13728
rect 2884 13688 3332 13716
rect 3326 13676 3332 13688
rect 3384 13676 3390 13728
rect 3436 13716 3464 13756
rect 4154 13744 4160 13756
rect 4212 13784 4218 13796
rect 4433 13787 4491 13793
rect 4433 13784 4445 13787
rect 4212 13756 4445 13784
rect 4212 13744 4218 13756
rect 4433 13753 4445 13756
rect 4479 13784 4491 13787
rect 4632 13784 4660 13824
rect 5169 13821 5181 13824
rect 5215 13821 5227 13855
rect 5169 13815 5227 13821
rect 5445 13855 5503 13861
rect 5445 13821 5457 13855
rect 5491 13821 5503 13855
rect 5445 13815 5503 13821
rect 5905 13855 5963 13861
rect 5905 13821 5917 13855
rect 5951 13852 5963 13855
rect 5994 13852 6000 13864
rect 5951 13824 6000 13852
rect 5951 13821 5963 13824
rect 5905 13815 5963 13821
rect 5994 13812 6000 13824
rect 6052 13812 6058 13864
rect 4479 13756 4660 13784
rect 5537 13787 5595 13793
rect 4479 13753 4491 13756
rect 4433 13747 4491 13753
rect 5537 13753 5549 13787
rect 5583 13753 5595 13787
rect 5537 13747 5595 13753
rect 4614 13716 4620 13728
rect 3436 13688 4620 13716
rect 4614 13676 4620 13688
rect 4672 13676 4678 13728
rect 5552 13716 5580 13747
rect 5626 13744 5632 13796
rect 5684 13784 5690 13796
rect 5767 13787 5825 13793
rect 5684 13756 5729 13784
rect 5684 13744 5690 13756
rect 5767 13753 5779 13787
rect 5813 13784 5825 13787
rect 6086 13784 6092 13796
rect 5813 13756 6092 13784
rect 5813 13753 5825 13756
rect 5767 13747 5825 13753
rect 6086 13744 6092 13756
rect 6144 13744 6150 13796
rect 6748 13716 6776 13892
rect 7101 13889 7113 13892
rect 7147 13920 7159 13923
rect 7190 13920 7196 13932
rect 7147 13892 7196 13920
rect 7147 13889 7159 13892
rect 7101 13883 7159 13889
rect 7190 13880 7196 13892
rect 7248 13880 7254 13932
rect 8312 13929 8340 13960
rect 9401 13957 9413 13960
rect 9447 13957 9459 13991
rect 9401 13951 9459 13957
rect 10505 13991 10563 13997
rect 10505 13957 10517 13991
rect 10551 13988 10563 13991
rect 11054 13988 11060 14000
rect 10551 13960 11060 13988
rect 10551 13957 10563 13960
rect 10505 13951 10563 13957
rect 11054 13948 11060 13960
rect 11112 13948 11118 14000
rect 11330 13948 11336 14000
rect 11388 13988 11394 14000
rect 11388 13960 12388 13988
rect 11388 13948 11394 13960
rect 8297 13923 8355 13929
rect 8297 13889 8309 13923
rect 8343 13889 8355 13923
rect 8297 13883 8355 13889
rect 8386 13880 8392 13932
rect 8444 13920 8450 13932
rect 8754 13920 8760 13932
rect 8444 13892 8489 13920
rect 8715 13892 8760 13920
rect 8444 13880 8450 13892
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 10045 13923 10103 13929
rect 10045 13889 10057 13923
rect 10091 13920 10103 13923
rect 10686 13920 10692 13932
rect 10091 13892 10692 13920
rect 10091 13889 10103 13892
rect 10045 13883 10103 13889
rect 6825 13855 6883 13861
rect 6825 13821 6837 13855
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 9582 13855 9640 13861
rect 9582 13821 9594 13855
rect 9628 13852 9640 13855
rect 10060 13852 10088 13883
rect 10686 13880 10692 13892
rect 10744 13880 10750 13932
rect 12360 13929 12388 13960
rect 12345 13923 12403 13929
rect 10796 13892 12296 13920
rect 10796 13861 10824 13892
rect 9628 13824 10088 13852
rect 10505 13855 10563 13861
rect 9628 13821 9640 13824
rect 9582 13815 9640 13821
rect 10505 13821 10517 13855
rect 10551 13852 10563 13855
rect 10597 13855 10655 13861
rect 10597 13852 10609 13855
rect 10551 13824 10609 13852
rect 10551 13821 10563 13824
rect 10505 13815 10563 13821
rect 10597 13821 10609 13824
rect 10643 13821 10655 13855
rect 10597 13815 10655 13821
rect 10781 13855 10839 13861
rect 10781 13821 10793 13855
rect 10827 13821 10839 13855
rect 10962 13852 10968 13864
rect 10923 13824 10968 13852
rect 10781 13815 10839 13821
rect 6840 13784 6868 13815
rect 10962 13812 10968 13824
rect 11020 13812 11026 13864
rect 7006 13784 7012 13796
rect 6840 13756 7012 13784
rect 7006 13744 7012 13756
rect 7064 13744 7070 13796
rect 10226 13744 10232 13796
rect 10284 13784 10290 13796
rect 10873 13787 10931 13793
rect 10873 13784 10885 13787
rect 10284 13756 10885 13784
rect 10284 13744 10290 13756
rect 10873 13753 10885 13756
rect 10919 13753 10931 13787
rect 12268 13784 12296 13892
rect 12345 13889 12357 13923
rect 12391 13889 12403 13923
rect 12618 13920 12624 13932
rect 12579 13892 12624 13920
rect 12345 13883 12403 13889
rect 12618 13880 12624 13892
rect 12676 13880 12682 13932
rect 14918 13920 14924 13932
rect 14879 13892 14924 13920
rect 14918 13880 14924 13892
rect 14976 13880 14982 13932
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 14645 13855 14703 13861
rect 14645 13852 14657 13855
rect 14424 13824 14657 13852
rect 14424 13812 14430 13824
rect 14645 13821 14657 13824
rect 14691 13821 14703 13855
rect 14645 13815 14703 13821
rect 12268 13756 12434 13784
rect 10873 13747 10931 13753
rect 12406 13728 12434 13756
rect 12526 13744 12532 13796
rect 12584 13784 12590 13796
rect 16206 13784 16212 13796
rect 12584 13756 13110 13784
rect 16146 13756 16212 13784
rect 12584 13744 12590 13756
rect 16206 13744 16212 13756
rect 16264 13744 16270 13796
rect 5552 13688 6776 13716
rect 7101 13719 7159 13725
rect 7101 13685 7113 13719
rect 7147 13716 7159 13719
rect 7650 13716 7656 13728
rect 7147 13688 7656 13716
rect 7147 13685 7159 13688
rect 7101 13679 7159 13685
rect 7650 13676 7656 13688
rect 7708 13676 7714 13728
rect 9585 13719 9643 13725
rect 9585 13685 9597 13719
rect 9631 13716 9643 13719
rect 9766 13716 9772 13728
rect 9631 13688 9772 13716
rect 9631 13685 9643 13688
rect 9585 13679 9643 13685
rect 9766 13676 9772 13688
rect 9824 13676 9830 13728
rect 12406 13688 12440 13728
rect 12434 13676 12440 13688
rect 12492 13676 12498 13728
rect 1104 13626 17296 13648
rect 1104 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 6571 13626
rect 6623 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 11904 13626
rect 11956 13574 11968 13626
rect 12020 13574 17296 13626
rect 1104 13552 17296 13574
rect 2866 13512 2872 13524
rect 1412 13484 2872 13512
rect 1412 13385 1440 13484
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 4246 13512 4252 13524
rect 2976 13484 4252 13512
rect 2976 13453 3004 13484
rect 4246 13472 4252 13484
rect 4304 13472 4310 13524
rect 7190 13512 7196 13524
rect 7151 13484 7196 13512
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 7926 13512 7932 13524
rect 7887 13484 7932 13512
rect 7926 13472 7932 13484
rect 7984 13472 7990 13524
rect 10686 13512 10692 13524
rect 10647 13484 10692 13512
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 10870 13512 10876 13524
rect 10831 13484 10876 13512
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 10962 13472 10968 13524
rect 11020 13512 11026 13524
rect 12897 13515 12955 13521
rect 11020 13484 12756 13512
rect 11020 13472 11026 13484
rect 2961 13447 3019 13453
rect 2961 13413 2973 13447
rect 3007 13413 3019 13447
rect 2961 13407 3019 13413
rect 3191 13447 3249 13453
rect 3191 13413 3203 13447
rect 3237 13444 3249 13447
rect 3510 13444 3516 13456
rect 3237 13416 3516 13444
rect 3237 13413 3249 13416
rect 3191 13407 3249 13413
rect 3510 13404 3516 13416
rect 3568 13404 3574 13456
rect 4433 13447 4491 13453
rect 4433 13413 4445 13447
rect 4479 13444 4491 13447
rect 4798 13444 4804 13456
rect 4479 13416 4804 13444
rect 4479 13413 4491 13416
rect 4433 13407 4491 13413
rect 4798 13404 4804 13416
rect 4856 13444 4862 13456
rect 5169 13447 5227 13453
rect 5169 13444 5181 13447
rect 4856 13416 5181 13444
rect 4856 13404 4862 13416
rect 5169 13413 5181 13416
rect 5215 13413 5227 13447
rect 5169 13407 5227 13413
rect 6181 13447 6239 13453
rect 6181 13413 6193 13447
rect 6227 13444 6239 13447
rect 7098 13444 7104 13456
rect 6227 13416 7104 13444
rect 6227 13413 6239 13416
rect 6181 13407 6239 13413
rect 7098 13404 7104 13416
rect 7156 13404 7162 13456
rect 7650 13404 7656 13456
rect 7708 13444 7714 13456
rect 7708 13416 9536 13444
rect 7708 13404 7714 13416
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13345 1455 13379
rect 1397 13339 1455 13345
rect 1762 13336 1768 13388
rect 1820 13376 1826 13388
rect 2041 13379 2099 13385
rect 2041 13376 2053 13379
rect 1820 13348 2053 13376
rect 1820 13336 1826 13348
rect 2041 13345 2053 13348
rect 2087 13345 2099 13379
rect 2041 13339 2099 13345
rect 2056 13308 2084 13339
rect 2774 13336 2780 13388
rect 2832 13376 2838 13388
rect 2869 13379 2927 13385
rect 2869 13376 2881 13379
rect 2832 13348 2881 13376
rect 2832 13336 2838 13348
rect 2869 13345 2881 13348
rect 2915 13345 2927 13379
rect 2869 13339 2927 13345
rect 3050 13336 3056 13388
rect 3108 13376 3114 13388
rect 4614 13376 4620 13388
rect 3108 13348 3832 13376
rect 4575 13348 4620 13376
rect 3108 13336 3114 13348
rect 3329 13311 3387 13317
rect 2056 13280 3004 13308
rect 2976 13252 3004 13280
rect 3329 13277 3341 13311
rect 3375 13308 3387 13311
rect 3602 13308 3608 13320
rect 3375 13280 3608 13308
rect 3375 13277 3387 13280
rect 3329 13271 3387 13277
rect 3602 13268 3608 13280
rect 3660 13268 3666 13320
rect 3804 13308 3832 13348
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 5074 13376 5080 13388
rect 5035 13348 5080 13376
rect 5074 13336 5080 13348
rect 5132 13336 5138 13388
rect 5902 13336 5908 13388
rect 5960 13385 5966 13388
rect 5960 13379 6009 13385
rect 5960 13345 5963 13379
rect 5997 13345 6009 13379
rect 6086 13376 6092 13388
rect 6047 13348 6092 13376
rect 5960 13339 6009 13345
rect 5960 13336 5966 13339
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 6365 13379 6423 13385
rect 6365 13345 6377 13379
rect 6411 13376 6423 13379
rect 6730 13376 6736 13388
rect 6411 13348 6736 13376
rect 6411 13345 6423 13348
rect 6365 13339 6423 13345
rect 6730 13336 6736 13348
rect 6788 13336 6794 13388
rect 6825 13379 6883 13385
rect 6825 13345 6837 13379
rect 6871 13345 6883 13379
rect 7006 13376 7012 13388
rect 6967 13348 7012 13376
rect 6825 13339 6883 13345
rect 5626 13308 5632 13320
rect 3804 13280 5632 13308
rect 5626 13268 5632 13280
rect 5684 13268 5690 13320
rect 6840 13308 6868 13339
rect 7006 13336 7012 13348
rect 7064 13336 7070 13388
rect 8202 13376 8208 13388
rect 8163 13348 8208 13376
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 9508 13385 9536 13416
rect 12434 13404 12440 13456
rect 12492 13444 12498 13456
rect 12621 13447 12679 13453
rect 12621 13444 12633 13447
rect 12492 13416 12633 13444
rect 12492 13404 12498 13416
rect 12621 13413 12633 13416
rect 12667 13413 12679 13447
rect 12621 13407 12679 13413
rect 9493 13379 9551 13385
rect 9493 13345 9505 13379
rect 9539 13345 9551 13379
rect 9493 13339 9551 13345
rect 10870 13379 10928 13385
rect 10870 13345 10882 13379
rect 10916 13376 10928 13379
rect 11606 13376 11612 13388
rect 10916 13348 11612 13376
rect 10916 13345 10928 13348
rect 10870 13339 10928 13345
rect 11606 13336 11612 13348
rect 11664 13336 11670 13388
rect 11977 13379 12035 13385
rect 11977 13345 11989 13379
rect 12023 13376 12035 13379
rect 12158 13376 12164 13388
rect 12023 13348 12164 13376
rect 12023 13345 12035 13348
rect 11977 13339 12035 13345
rect 12158 13336 12164 13348
rect 12216 13376 12222 13388
rect 12342 13376 12348 13388
rect 12216 13348 12348 13376
rect 12216 13336 12222 13348
rect 12342 13336 12348 13348
rect 12400 13336 12406 13388
rect 12728 13376 12756 13484
rect 12897 13481 12909 13515
rect 12943 13512 12955 13515
rect 13078 13512 13084 13524
rect 12943 13484 13084 13512
rect 12943 13481 12955 13484
rect 12897 13475 12955 13481
rect 13078 13472 13084 13484
rect 13136 13472 13142 13524
rect 15010 13512 15016 13524
rect 14971 13484 15016 13512
rect 15010 13472 15016 13484
rect 15068 13472 15074 13524
rect 16025 13515 16083 13521
rect 16025 13481 16037 13515
rect 16071 13512 16083 13515
rect 16298 13512 16304 13524
rect 16071 13484 16304 13512
rect 16071 13481 16083 13484
rect 16025 13475 16083 13481
rect 12805 13447 12863 13453
rect 12805 13413 12817 13447
rect 12851 13444 12863 13447
rect 13170 13444 13176 13456
rect 12851 13416 13176 13444
rect 12851 13413 12863 13416
rect 12805 13407 12863 13413
rect 13170 13404 13176 13416
rect 13228 13444 13234 13456
rect 13725 13447 13783 13453
rect 13725 13444 13737 13447
rect 13228 13416 13737 13444
rect 13228 13404 13234 13416
rect 13725 13413 13737 13416
rect 13771 13413 13783 13447
rect 15197 13447 15255 13453
rect 15197 13444 15209 13447
rect 13725 13407 13783 13413
rect 14936 13416 15209 13444
rect 12989 13379 13047 13385
rect 12989 13376 13001 13379
rect 12728 13348 13001 13376
rect 12820 13320 12848 13348
rect 12989 13345 13001 13348
rect 13035 13345 13047 13379
rect 12989 13339 13047 13345
rect 13262 13336 13268 13388
rect 13320 13376 13326 13388
rect 14936 13385 14964 13416
rect 15197 13413 15209 13416
rect 15243 13444 15255 13447
rect 15746 13444 15752 13456
rect 15243 13416 15752 13444
rect 15243 13413 15255 13416
rect 15197 13407 15255 13413
rect 15746 13404 15752 13416
rect 15804 13404 15810 13456
rect 16040 13444 16068 13475
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 15948 13416 16068 13444
rect 13633 13379 13691 13385
rect 13633 13376 13645 13379
rect 13320 13348 13645 13376
rect 13320 13336 13326 13348
rect 13633 13345 13645 13348
rect 13679 13345 13691 13379
rect 13633 13339 13691 13345
rect 14737 13379 14795 13385
rect 14737 13345 14749 13379
rect 14783 13345 14795 13379
rect 14737 13339 14795 13345
rect 14921 13379 14979 13385
rect 14921 13345 14933 13379
rect 14967 13345 14979 13379
rect 14921 13339 14979 13345
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13345 15347 13379
rect 15838 13376 15844 13388
rect 15799 13348 15844 13376
rect 15289 13339 15347 13345
rect 5828 13280 6868 13308
rect 1581 13243 1639 13249
rect 1581 13209 1593 13243
rect 1627 13240 1639 13243
rect 1627 13212 2912 13240
rect 1627 13209 1639 13212
rect 1581 13203 1639 13209
rect 2222 13172 2228 13184
rect 2183 13144 2228 13172
rect 2222 13132 2228 13144
rect 2280 13132 2286 13184
rect 2682 13172 2688 13184
rect 2643 13144 2688 13172
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 2884 13172 2912 13212
rect 2958 13200 2964 13252
rect 3016 13200 3022 13252
rect 4338 13240 4344 13252
rect 3068 13212 4344 13240
rect 3068 13172 3096 13212
rect 4338 13200 4344 13212
rect 4396 13200 4402 13252
rect 5828 13184 5856 13280
rect 7834 13268 7840 13320
rect 7892 13308 7898 13320
rect 7929 13311 7987 13317
rect 7929 13308 7941 13311
rect 7892 13280 7941 13308
rect 7892 13268 7898 13280
rect 7929 13277 7941 13280
rect 7975 13277 7987 13311
rect 8110 13308 8116 13320
rect 8071 13280 8116 13308
rect 7929 13271 7987 13277
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 11330 13308 11336 13320
rect 11291 13280 11336 13308
rect 11330 13268 11336 13280
rect 11388 13268 11394 13320
rect 12802 13268 12808 13320
rect 12860 13268 12866 13320
rect 14752 13308 14780 13339
rect 15304 13308 15332 13339
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 15562 13308 15568 13320
rect 14752 13280 15568 13308
rect 15562 13268 15568 13280
rect 15620 13308 15626 13320
rect 15948 13308 15976 13416
rect 16117 13379 16175 13385
rect 16117 13345 16129 13379
rect 16163 13376 16175 13379
rect 16482 13376 16488 13388
rect 16163 13348 16488 13376
rect 16163 13345 16175 13348
rect 16117 13339 16175 13345
rect 15620 13280 15976 13308
rect 15620 13268 15626 13280
rect 5902 13200 5908 13252
rect 5960 13240 5966 13252
rect 6178 13240 6184 13252
rect 5960 13212 6184 13240
rect 5960 13200 5966 13212
rect 6178 13200 6184 13212
rect 6236 13200 6242 13252
rect 7374 13200 7380 13252
rect 7432 13240 7438 13252
rect 9585 13243 9643 13249
rect 9585 13240 9597 13243
rect 7432 13212 9597 13240
rect 7432 13200 7438 13212
rect 9585 13209 9597 13212
rect 9631 13209 9643 13243
rect 9585 13203 9643 13209
rect 14826 13200 14832 13252
rect 14884 13240 14890 13252
rect 16132 13240 16160 13339
rect 16482 13336 16488 13348
rect 16540 13336 16546 13388
rect 14884 13212 16160 13240
rect 14884 13200 14890 13212
rect 5810 13172 5816 13184
rect 2884 13144 3096 13172
rect 5771 13144 5816 13172
rect 5810 13132 5816 13144
rect 5868 13132 5874 13184
rect 6730 13132 6736 13184
rect 6788 13172 6794 13184
rect 7190 13172 7196 13184
rect 6788 13144 7196 13172
rect 6788 13132 6794 13144
rect 7190 13132 7196 13144
rect 7248 13132 7254 13184
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 11241 13175 11299 13181
rect 11241 13172 11253 13175
rect 11112 13144 11253 13172
rect 11112 13132 11118 13144
rect 11241 13141 11253 13144
rect 11287 13141 11299 13175
rect 11790 13172 11796 13184
rect 11751 13144 11796 13172
rect 11241 13135 11299 13141
rect 11790 13132 11796 13144
rect 11848 13132 11854 13184
rect 13170 13172 13176 13184
rect 13131 13144 13176 13172
rect 13170 13132 13176 13144
rect 13228 13132 13234 13184
rect 1104 13082 17296 13104
rect 1104 13030 3680 13082
rect 3732 13030 3744 13082
rect 3796 13030 3808 13082
rect 3860 13030 3872 13082
rect 3924 13030 9078 13082
rect 9130 13030 9142 13082
rect 9194 13030 9206 13082
rect 9258 13030 9270 13082
rect 9322 13030 14475 13082
rect 14527 13030 14539 13082
rect 14591 13030 14603 13082
rect 14655 13030 14667 13082
rect 14719 13030 17296 13082
rect 1104 13008 17296 13030
rect 1394 12968 1400 12980
rect 1307 12940 1400 12968
rect 1394 12928 1400 12940
rect 1452 12968 1458 12980
rect 3145 12971 3203 12977
rect 1452 12940 2728 12968
rect 1452 12928 1458 12940
rect 1412 12841 1440 12928
rect 2700 12900 2728 12940
rect 3145 12937 3157 12971
rect 3191 12968 3203 12971
rect 3234 12968 3240 12980
rect 3191 12940 3240 12968
rect 3191 12937 3203 12940
rect 3145 12931 3203 12937
rect 3234 12928 3240 12940
rect 3292 12968 3298 12980
rect 3510 12968 3516 12980
rect 3292 12940 3516 12968
rect 3292 12928 3298 12940
rect 3510 12928 3516 12940
rect 3568 12928 3574 12980
rect 4341 12971 4399 12977
rect 4341 12937 4353 12971
rect 4387 12968 4399 12971
rect 4433 12971 4491 12977
rect 4433 12968 4445 12971
rect 4387 12940 4445 12968
rect 4387 12937 4399 12940
rect 4341 12931 4399 12937
rect 4433 12937 4445 12940
rect 4479 12968 4491 12971
rect 7006 12968 7012 12980
rect 4479 12940 7012 12968
rect 4479 12937 4491 12940
rect 4433 12931 4491 12937
rect 7006 12928 7012 12940
rect 7064 12928 7070 12980
rect 7834 12968 7840 12980
rect 7795 12940 7840 12968
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 11054 12968 11060 12980
rect 11015 12940 11060 12968
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 11330 12928 11336 12980
rect 11388 12968 11394 12980
rect 12069 12971 12127 12977
rect 12069 12968 12081 12971
rect 11388 12940 12081 12968
rect 11388 12928 11394 12940
rect 12069 12937 12081 12940
rect 12115 12937 12127 12971
rect 12069 12931 12127 12937
rect 12897 12971 12955 12977
rect 12897 12937 12909 12971
rect 12943 12968 12955 12971
rect 13814 12968 13820 12980
rect 12943 12940 13820 12968
rect 12943 12937 12955 12940
rect 12897 12931 12955 12937
rect 13814 12928 13820 12940
rect 13872 12968 13878 12980
rect 14645 12971 14703 12977
rect 14645 12968 14657 12971
rect 13872 12940 14657 12968
rect 13872 12928 13878 12940
rect 14645 12937 14657 12940
rect 14691 12968 14703 12971
rect 14826 12968 14832 12980
rect 14691 12940 14832 12968
rect 14691 12937 14703 12940
rect 14645 12931 14703 12937
rect 14826 12928 14832 12940
rect 14884 12928 14890 12980
rect 16206 12968 16212 12980
rect 16167 12940 16212 12968
rect 16206 12928 16212 12940
rect 16264 12928 16270 12980
rect 4982 12900 4988 12912
rect 2700 12872 4988 12900
rect 4982 12860 4988 12872
rect 5040 12860 5046 12912
rect 5626 12860 5632 12912
rect 5684 12900 5690 12912
rect 8110 12900 8116 12912
rect 5684 12872 8116 12900
rect 5684 12860 5690 12872
rect 8110 12860 8116 12872
rect 8168 12860 8174 12912
rect 15197 12903 15255 12909
rect 15197 12900 15209 12903
rect 10796 12872 15209 12900
rect 1397 12835 1455 12841
rect 1397 12801 1409 12835
rect 1443 12801 1455 12835
rect 1397 12795 1455 12801
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 2682 12832 2688 12844
rect 1719 12804 2688 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 2682 12792 2688 12804
rect 2740 12792 2746 12844
rect 3142 12792 3148 12844
rect 3200 12832 3206 12844
rect 3510 12832 3516 12844
rect 3200 12804 3516 12832
rect 3200 12792 3206 12804
rect 3510 12792 3516 12804
rect 3568 12792 3574 12844
rect 4798 12832 4804 12844
rect 4759 12804 4804 12832
rect 4798 12792 4804 12804
rect 4856 12792 4862 12844
rect 4893 12835 4951 12841
rect 4893 12801 4905 12835
rect 4939 12832 4951 12835
rect 5994 12832 6000 12844
rect 4939 12804 6000 12832
rect 4939 12801 4951 12804
rect 4893 12795 4951 12801
rect 5994 12792 6000 12804
rect 6052 12792 6058 12844
rect 7926 12792 7932 12844
rect 7984 12832 7990 12844
rect 8573 12835 8631 12841
rect 8573 12832 8585 12835
rect 7984 12804 8585 12832
rect 7984 12792 7990 12804
rect 8573 12801 8585 12804
rect 8619 12801 8631 12835
rect 8573 12795 8631 12801
rect 10796 12776 10824 12872
rect 15197 12869 15209 12872
rect 15243 12869 15255 12903
rect 15197 12863 15255 12869
rect 10870 12792 10876 12844
rect 10928 12832 10934 12844
rect 12713 12835 12771 12841
rect 10928 12804 12112 12832
rect 10928 12792 10934 12804
rect 12084 12776 12112 12804
rect 12713 12801 12725 12835
rect 12759 12832 12771 12835
rect 13630 12832 13636 12844
rect 12759 12804 13636 12832
rect 12759 12801 12771 12804
rect 12713 12795 12771 12801
rect 13630 12792 13636 12804
rect 13688 12792 13694 12844
rect 3326 12724 3332 12776
rect 3384 12764 3390 12776
rect 3697 12767 3755 12773
rect 3697 12764 3709 12767
rect 3384 12736 3709 12764
rect 3384 12724 3390 12736
rect 3697 12733 3709 12736
rect 3743 12733 3755 12767
rect 3697 12727 3755 12733
rect 3789 12767 3847 12773
rect 3789 12733 3801 12767
rect 3835 12764 3847 12767
rect 4614 12764 4620 12776
rect 3835 12736 4620 12764
rect 3835 12733 3847 12736
rect 3789 12727 3847 12733
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 4706 12724 4712 12776
rect 4764 12764 4770 12776
rect 5074 12764 5080 12776
rect 4764 12736 4809 12764
rect 5035 12736 5080 12764
rect 4764 12724 4770 12736
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 5905 12767 5963 12773
rect 5905 12733 5917 12767
rect 5951 12733 5963 12767
rect 5905 12727 5963 12733
rect 2222 12656 2228 12708
rect 2280 12656 2286 12708
rect 5920 12696 5948 12727
rect 6730 12724 6736 12776
rect 6788 12764 6794 12776
rect 7374 12773 7380 12776
rect 7193 12767 7251 12773
rect 7193 12764 7205 12767
rect 6788 12736 7205 12764
rect 6788 12724 6794 12736
rect 7193 12733 7205 12736
rect 7239 12733 7251 12767
rect 7193 12727 7251 12733
rect 7341 12767 7380 12773
rect 7341 12733 7353 12767
rect 7341 12727 7380 12733
rect 7374 12724 7380 12727
rect 7432 12724 7438 12776
rect 7650 12724 7656 12776
rect 7708 12773 7714 12776
rect 7708 12764 7716 12773
rect 8297 12767 8355 12773
rect 7708 12736 7753 12764
rect 7708 12727 7716 12736
rect 8297 12733 8309 12767
rect 8343 12733 8355 12767
rect 10778 12764 10784 12776
rect 10691 12736 10784 12764
rect 8297 12727 8355 12733
rect 7708 12724 7714 12727
rect 7466 12696 7472 12708
rect 5920 12668 7472 12696
rect 7466 12656 7472 12668
rect 7524 12656 7530 12708
rect 7561 12699 7619 12705
rect 7561 12665 7573 12699
rect 7607 12665 7619 12699
rect 8312 12696 8340 12727
rect 10778 12724 10784 12736
rect 10836 12764 10842 12776
rect 10965 12767 11023 12773
rect 10965 12764 10977 12767
rect 10836 12736 10977 12764
rect 10836 12724 10842 12736
rect 10965 12733 10977 12736
rect 11011 12733 11023 12767
rect 12066 12764 12072 12776
rect 11979 12736 12072 12764
rect 10965 12727 11023 12733
rect 12066 12724 12072 12736
rect 12124 12724 12130 12776
rect 12250 12764 12256 12776
rect 12211 12736 12256 12764
rect 12250 12724 12256 12736
rect 12308 12724 12314 12776
rect 12986 12724 12992 12776
rect 13044 12764 13050 12776
rect 13044 12736 13089 12764
rect 13044 12724 13050 12736
rect 13170 12724 13176 12776
rect 13228 12764 13234 12776
rect 13909 12767 13967 12773
rect 13909 12764 13921 12767
rect 13228 12736 13921 12764
rect 13228 12724 13234 12736
rect 13909 12733 13921 12736
rect 13955 12733 13967 12767
rect 13909 12727 13967 12733
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 14553 12767 14611 12773
rect 14553 12764 14565 12767
rect 14148 12736 14565 12764
rect 14148 12724 14154 12736
rect 14553 12733 14565 12736
rect 14599 12733 14611 12767
rect 15378 12764 15384 12776
rect 15339 12736 15384 12764
rect 14553 12727 14611 12733
rect 15378 12724 15384 12736
rect 15436 12724 15442 12776
rect 15562 12764 15568 12776
rect 15523 12736 15568 12764
rect 15562 12724 15568 12736
rect 15620 12724 15626 12776
rect 15746 12764 15752 12776
rect 15707 12736 15752 12764
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 16298 12724 16304 12776
rect 16356 12764 16362 12776
rect 16393 12767 16451 12773
rect 16393 12764 16405 12767
rect 16356 12736 16405 12764
rect 16356 12724 16362 12736
rect 16393 12733 16405 12736
rect 16439 12733 16451 12767
rect 16393 12727 16451 12733
rect 8478 12696 8484 12708
rect 8312 12668 8484 12696
rect 7561 12659 7619 12665
rect 3326 12588 3332 12640
rect 3384 12628 3390 12640
rect 4341 12631 4399 12637
rect 4341 12628 4353 12631
rect 3384 12600 4353 12628
rect 3384 12588 3390 12600
rect 4341 12597 4353 12600
rect 4387 12597 4399 12631
rect 4341 12591 4399 12597
rect 5813 12631 5871 12637
rect 5813 12597 5825 12631
rect 5859 12628 5871 12631
rect 7576 12628 7604 12659
rect 8478 12656 8484 12668
rect 8536 12656 8542 12708
rect 11790 12696 11796 12708
rect 9798 12668 11796 12696
rect 11790 12656 11796 12668
rect 11848 12656 11854 12708
rect 13722 12696 13728 12708
rect 13683 12668 13728 12696
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 15470 12696 15476 12708
rect 15431 12668 15476 12696
rect 15470 12656 15476 12668
rect 15528 12656 15534 12708
rect 5859 12600 7604 12628
rect 5859 12597 5871 12600
rect 5813 12591 5871 12597
rect 7834 12588 7840 12640
rect 7892 12628 7898 12640
rect 9490 12628 9496 12640
rect 7892 12600 9496 12628
rect 7892 12588 7898 12600
rect 9490 12588 9496 12600
rect 9548 12628 9554 12640
rect 10045 12631 10103 12637
rect 10045 12628 10057 12631
rect 9548 12600 10057 12628
rect 9548 12588 9554 12600
rect 10045 12597 10057 12600
rect 10091 12597 10103 12631
rect 12710 12628 12716 12640
rect 12671 12600 12716 12628
rect 10045 12591 10103 12597
rect 12710 12588 12716 12600
rect 12768 12588 12774 12640
rect 14090 12628 14096 12640
rect 14051 12600 14096 12628
rect 14090 12588 14096 12600
rect 14148 12588 14154 12640
rect 1104 12538 17296 12560
rect 1104 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 6571 12538
rect 6623 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 11904 12538
rect 11956 12486 11968 12538
rect 12020 12486 17296 12538
rect 1104 12464 17296 12486
rect 3329 12427 3387 12433
rect 3329 12393 3341 12427
rect 3375 12424 3387 12427
rect 3970 12424 3976 12436
rect 3375 12396 3976 12424
rect 3375 12393 3387 12396
rect 3329 12387 3387 12393
rect 3970 12384 3976 12396
rect 4028 12384 4034 12436
rect 4246 12384 4252 12436
rect 4304 12384 4310 12436
rect 7282 12424 7288 12436
rect 5920 12396 7288 12424
rect 2314 12356 2320 12368
rect 1872 12328 2320 12356
rect 1872 12297 1900 12328
rect 2314 12316 2320 12328
rect 2372 12316 2378 12368
rect 1857 12291 1915 12297
rect 1857 12257 1869 12291
rect 1903 12257 1915 12291
rect 1857 12251 1915 12257
rect 2038 12248 2044 12300
rect 2096 12288 2102 12300
rect 2501 12291 2559 12297
rect 2501 12288 2513 12291
rect 2096 12260 2513 12288
rect 2096 12248 2102 12260
rect 2501 12257 2513 12260
rect 2547 12257 2559 12291
rect 3142 12288 3148 12300
rect 3103 12260 3148 12288
rect 2501 12251 2559 12257
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 3326 12288 3332 12300
rect 3287 12260 3332 12288
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 4264 12229 4292 12384
rect 4525 12291 4583 12297
rect 4525 12288 4537 12291
rect 4356 12260 4537 12288
rect 4249 12223 4307 12229
rect 4249 12189 4261 12223
rect 4295 12189 4307 12223
rect 4249 12183 4307 12189
rect 4062 12112 4068 12164
rect 4120 12152 4126 12164
rect 4356 12152 4384 12260
rect 4525 12257 4537 12260
rect 4571 12257 4583 12291
rect 4525 12251 4583 12257
rect 4706 12248 4712 12300
rect 4764 12288 4770 12300
rect 5169 12291 5227 12297
rect 5169 12288 5181 12291
rect 4764 12260 5181 12288
rect 4764 12248 4770 12260
rect 5169 12257 5181 12260
rect 5215 12288 5227 12291
rect 5350 12288 5356 12300
rect 5215 12260 5356 12288
rect 5215 12257 5227 12260
rect 5169 12251 5227 12257
rect 5350 12248 5356 12260
rect 5408 12248 5414 12300
rect 5920 12297 5948 12396
rect 7282 12384 7288 12396
rect 7340 12384 7346 12436
rect 7466 12424 7472 12436
rect 7427 12396 7472 12424
rect 7466 12384 7472 12396
rect 7524 12384 7530 12436
rect 8662 12384 8668 12436
rect 8720 12424 8726 12436
rect 10689 12427 10747 12433
rect 10689 12424 10701 12427
rect 8720 12396 10701 12424
rect 8720 12384 8726 12396
rect 10689 12393 10701 12396
rect 10735 12393 10747 12427
rect 12250 12424 12256 12436
rect 10689 12387 10747 12393
rect 11992 12396 12256 12424
rect 6086 12316 6092 12368
rect 6144 12356 6150 12368
rect 6638 12356 6644 12368
rect 6144 12328 6644 12356
rect 6144 12316 6150 12328
rect 6638 12316 6644 12328
rect 6696 12316 6702 12368
rect 7834 12356 7840 12368
rect 6932 12328 7840 12356
rect 5905 12291 5963 12297
rect 5905 12257 5917 12291
rect 5951 12257 5963 12291
rect 5905 12251 5963 12257
rect 6546 12248 6552 12300
rect 6604 12288 6610 12300
rect 6604 12260 6649 12288
rect 6604 12248 6610 12260
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12220 4491 12223
rect 5074 12220 5080 12232
rect 4479 12192 5080 12220
rect 4479 12189 4491 12192
rect 4433 12183 4491 12189
rect 5074 12180 5080 12192
rect 5132 12180 5138 12232
rect 6733 12223 6791 12229
rect 6733 12220 6745 12223
rect 6564 12192 6745 12220
rect 6564 12164 6592 12192
rect 6733 12189 6745 12192
rect 6779 12189 6791 12223
rect 6733 12183 6791 12189
rect 6842 12223 6900 12229
rect 6842 12189 6854 12223
rect 6888 12220 6900 12223
rect 6932 12220 6960 12328
rect 7834 12316 7840 12328
rect 7892 12316 7898 12368
rect 11330 12316 11336 12368
rect 11388 12356 11394 12368
rect 11793 12359 11851 12365
rect 11793 12356 11805 12359
rect 11388 12328 11805 12356
rect 11388 12316 11394 12328
rect 11793 12325 11805 12328
rect 11839 12325 11851 12359
rect 11793 12319 11851 12325
rect 7009 12291 7067 12297
rect 7009 12257 7021 12291
rect 7055 12288 7067 12291
rect 7190 12288 7196 12300
rect 7055 12260 7196 12288
rect 7055 12257 7067 12260
rect 7009 12251 7067 12257
rect 7190 12248 7196 12260
rect 7248 12248 7254 12300
rect 7650 12288 7656 12300
rect 7611 12260 7656 12288
rect 7650 12248 7656 12260
rect 7708 12248 7714 12300
rect 7745 12291 7803 12297
rect 7745 12257 7757 12291
rect 7791 12257 7803 12291
rect 7745 12251 7803 12257
rect 8021 12291 8079 12297
rect 8021 12257 8033 12291
rect 8067 12288 8079 12291
rect 8202 12288 8208 12300
rect 8067 12260 8208 12288
rect 8067 12257 8079 12260
rect 8021 12251 8079 12257
rect 6888 12192 6960 12220
rect 7208 12220 7236 12248
rect 7374 12220 7380 12232
rect 7208 12192 7380 12220
rect 6888 12189 6900 12192
rect 6842 12183 6900 12189
rect 7374 12180 7380 12192
rect 7432 12220 7438 12232
rect 7760 12220 7788 12251
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 9490 12288 9496 12300
rect 9451 12260 9496 12288
rect 9490 12248 9496 12260
rect 9548 12248 9554 12300
rect 10778 12248 10784 12300
rect 10836 12288 10842 12300
rect 10873 12291 10931 12297
rect 10873 12288 10885 12291
rect 10836 12260 10885 12288
rect 10836 12248 10842 12260
rect 10873 12257 10885 12260
rect 10919 12257 10931 12291
rect 10873 12251 10931 12257
rect 10965 12291 11023 12297
rect 10965 12257 10977 12291
rect 11011 12288 11023 12291
rect 11241 12291 11299 12297
rect 11241 12288 11253 12291
rect 11011 12260 11253 12288
rect 11011 12257 11023 12260
rect 10965 12251 11023 12257
rect 11241 12257 11253 12260
rect 11287 12288 11299 12291
rect 11287 12260 11468 12288
rect 11287 12257 11299 12260
rect 11241 12251 11299 12257
rect 7432 12192 7788 12220
rect 8220 12220 8248 12248
rect 9585 12223 9643 12229
rect 9585 12220 9597 12223
rect 8220 12192 9597 12220
rect 7432 12180 7438 12192
rect 9585 12189 9597 12192
rect 9631 12189 9643 12223
rect 10888 12220 10916 12251
rect 11333 12223 11391 12229
rect 11333 12220 11345 12223
rect 10888 12192 11345 12220
rect 9585 12183 9643 12189
rect 11333 12189 11345 12192
rect 11379 12189 11391 12223
rect 11333 12183 11391 12189
rect 4120 12124 4384 12152
rect 4120 12112 4126 12124
rect 5626 12112 5632 12164
rect 5684 12152 5690 12164
rect 6362 12152 6368 12164
rect 5684 12124 6368 12152
rect 5684 12112 5690 12124
rect 6362 12112 6368 12124
rect 6420 12112 6426 12164
rect 6546 12112 6552 12164
rect 6604 12112 6610 12164
rect 6641 12155 6699 12161
rect 6641 12121 6653 12155
rect 6687 12152 6699 12155
rect 7466 12152 7472 12164
rect 6687 12124 7472 12152
rect 6687 12121 6699 12124
rect 6641 12115 6699 12121
rect 7466 12112 7472 12124
rect 7524 12112 7530 12164
rect 11440 12152 11468 12260
rect 11606 12248 11612 12300
rect 11664 12288 11670 12300
rect 11992 12297 12020 12396
rect 12250 12384 12256 12396
rect 12308 12424 12314 12436
rect 12308 12396 13676 12424
rect 12308 12384 12314 12396
rect 13262 12356 13268 12368
rect 12912 12328 13268 12356
rect 11977 12291 12035 12297
rect 11977 12288 11989 12291
rect 11664 12260 11989 12288
rect 11664 12248 11670 12260
rect 11977 12257 11989 12260
rect 12023 12257 12035 12291
rect 11977 12251 12035 12257
rect 12066 12248 12072 12300
rect 12124 12288 12130 12300
rect 12124 12260 12169 12288
rect 12124 12248 12130 12260
rect 12710 12248 12716 12300
rect 12768 12288 12774 12300
rect 12912 12297 12940 12328
rect 13262 12316 13268 12328
rect 13320 12316 13326 12368
rect 12805 12291 12863 12297
rect 12805 12288 12817 12291
rect 12768 12260 12817 12288
rect 12768 12248 12774 12260
rect 12805 12257 12817 12260
rect 12851 12257 12863 12291
rect 12805 12251 12863 12257
rect 12897 12291 12955 12297
rect 12897 12257 12909 12291
rect 12943 12257 12955 12291
rect 12897 12251 12955 12257
rect 13081 12291 13139 12297
rect 13081 12257 13093 12291
rect 13127 12288 13139 12291
rect 13170 12288 13176 12300
rect 13127 12260 13176 12288
rect 13127 12257 13139 12260
rect 13081 12251 13139 12257
rect 13170 12248 13176 12260
rect 13228 12248 13234 12300
rect 13648 12297 13676 12396
rect 15102 12384 15108 12436
rect 15160 12424 15166 12436
rect 16393 12427 16451 12433
rect 16393 12424 16405 12427
rect 15160 12396 16405 12424
rect 15160 12384 15166 12396
rect 16393 12393 16405 12396
rect 16439 12393 16451 12427
rect 16393 12387 16451 12393
rect 15378 12356 15384 12368
rect 15291 12328 15384 12356
rect 15378 12316 15384 12328
rect 15436 12356 15442 12368
rect 15930 12356 15936 12368
rect 15436 12328 15936 12356
rect 15436 12316 15442 12328
rect 15930 12316 15936 12328
rect 15988 12316 15994 12368
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12257 13691 12291
rect 13633 12251 13691 12257
rect 14274 12248 14280 12300
rect 14332 12288 14338 12300
rect 15289 12291 15347 12297
rect 15289 12288 15301 12291
rect 14332 12260 15301 12288
rect 14332 12248 14338 12260
rect 15289 12257 15301 12260
rect 15335 12257 15347 12291
rect 15470 12288 15476 12300
rect 15431 12260 15476 12288
rect 15289 12251 15347 12257
rect 15470 12248 15476 12260
rect 15528 12248 15534 12300
rect 15654 12288 15660 12300
rect 15615 12260 15660 12288
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 16574 12288 16580 12300
rect 16535 12260 16580 12288
rect 16574 12248 16580 12260
rect 16632 12248 16638 12300
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 11793 12155 11851 12161
rect 11793 12152 11805 12155
rect 11440 12124 11805 12152
rect 11793 12121 11805 12124
rect 11839 12121 11851 12155
rect 11793 12115 11851 12121
rect 12802 12112 12808 12164
rect 12860 12152 12866 12164
rect 13004 12152 13032 12183
rect 14274 12152 14280 12164
rect 12860 12124 14280 12152
rect 12860 12112 12866 12124
rect 14274 12112 14280 12124
rect 14332 12112 14338 12164
rect 2041 12087 2099 12093
rect 2041 12053 2053 12087
rect 2087 12084 2099 12087
rect 2222 12084 2228 12096
rect 2087 12056 2228 12084
rect 2087 12053 2099 12056
rect 2041 12047 2099 12053
rect 2222 12044 2228 12056
rect 2280 12044 2286 12096
rect 2685 12087 2743 12093
rect 2685 12053 2697 12087
rect 2731 12084 2743 12087
rect 2774 12084 2780 12096
rect 2731 12056 2780 12084
rect 2731 12053 2743 12056
rect 2685 12047 2743 12053
rect 2774 12044 2780 12056
rect 2832 12044 2838 12096
rect 4246 12044 4252 12096
rect 4304 12084 4310 12096
rect 4341 12087 4399 12093
rect 4341 12084 4353 12087
rect 4304 12056 4353 12084
rect 4304 12044 4310 12056
rect 4341 12053 4353 12056
rect 4387 12053 4399 12087
rect 4341 12047 4399 12053
rect 4614 12044 4620 12096
rect 4672 12084 4678 12096
rect 5077 12087 5135 12093
rect 5077 12084 5089 12087
rect 4672 12056 5089 12084
rect 4672 12044 4678 12056
rect 5077 12053 5089 12056
rect 5123 12053 5135 12087
rect 5810 12084 5816 12096
rect 5771 12056 5816 12084
rect 5077 12047 5135 12053
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 6178 12044 6184 12096
rect 6236 12084 6242 12096
rect 7742 12084 7748 12096
rect 6236 12056 7748 12084
rect 6236 12044 6242 12056
rect 7742 12044 7748 12056
rect 7800 12084 7806 12096
rect 7929 12087 7987 12093
rect 7929 12084 7941 12087
rect 7800 12056 7941 12084
rect 7800 12044 7806 12056
rect 7929 12053 7941 12056
rect 7975 12053 7987 12087
rect 12618 12084 12624 12096
rect 12579 12056 12624 12084
rect 7929 12047 7987 12053
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 13078 12044 13084 12096
rect 13136 12084 13142 12096
rect 13630 12084 13636 12096
rect 13136 12056 13636 12084
rect 13136 12044 13142 12056
rect 13630 12044 13636 12056
rect 13688 12084 13694 12096
rect 13725 12087 13783 12093
rect 13725 12084 13737 12087
rect 13688 12056 13737 12084
rect 13688 12044 13694 12056
rect 13725 12053 13737 12056
rect 13771 12053 13783 12087
rect 15102 12084 15108 12096
rect 15063 12056 15108 12084
rect 13725 12047 13783 12053
rect 15102 12044 15108 12056
rect 15160 12044 15166 12096
rect 1104 11994 17296 12016
rect 1104 11942 3680 11994
rect 3732 11942 3744 11994
rect 3796 11942 3808 11994
rect 3860 11942 3872 11994
rect 3924 11942 9078 11994
rect 9130 11942 9142 11994
rect 9194 11942 9206 11994
rect 9258 11942 9270 11994
rect 9322 11942 14475 11994
rect 14527 11942 14539 11994
rect 14591 11942 14603 11994
rect 14655 11942 14667 11994
rect 14719 11942 17296 11994
rect 1104 11920 17296 11942
rect 4154 11840 4160 11892
rect 4212 11880 4218 11892
rect 4212 11852 4476 11880
rect 4212 11840 4218 11852
rect 4448 11812 4476 11852
rect 4522 11840 4528 11892
rect 4580 11880 4586 11892
rect 4890 11880 4896 11892
rect 4580 11852 4896 11880
rect 4580 11840 4586 11852
rect 4890 11840 4896 11852
rect 4948 11840 4954 11892
rect 5350 11880 5356 11892
rect 5311 11852 5356 11880
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 5813 11883 5871 11889
rect 5813 11849 5825 11883
rect 5859 11880 5871 11883
rect 6178 11880 6184 11892
rect 5859 11852 6184 11880
rect 5859 11849 5871 11852
rect 5813 11843 5871 11849
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 12253 11883 12311 11889
rect 12253 11849 12265 11883
rect 12299 11880 12311 11883
rect 12526 11880 12532 11892
rect 12299 11852 12532 11880
rect 12299 11849 12311 11852
rect 12253 11843 12311 11849
rect 12526 11840 12532 11852
rect 12584 11840 12590 11892
rect 13081 11883 13139 11889
rect 13081 11849 13093 11883
rect 13127 11880 13139 11883
rect 13541 11883 13599 11889
rect 13127 11852 13492 11880
rect 13127 11849 13139 11852
rect 13081 11843 13139 11849
rect 12713 11815 12771 11821
rect 4448 11784 4757 11812
rect 2314 11704 2320 11756
rect 2372 11744 2378 11756
rect 2593 11747 2651 11753
rect 2593 11744 2605 11747
rect 2372 11716 2605 11744
rect 2372 11704 2378 11716
rect 2593 11713 2605 11716
rect 2639 11713 2651 11747
rect 4522 11744 4528 11756
rect 2593 11707 2651 11713
rect 4264 11716 4528 11744
rect 3789 11679 3847 11685
rect 3789 11645 3801 11679
rect 3835 11676 3847 11679
rect 4154 11676 4160 11688
rect 3835 11648 4160 11676
rect 3835 11645 3847 11648
rect 3789 11639 3847 11645
rect 4154 11636 4160 11648
rect 4212 11636 4218 11688
rect 4264 11685 4292 11716
rect 4522 11704 4528 11716
rect 4580 11704 4586 11756
rect 4249 11679 4307 11685
rect 4249 11645 4261 11679
rect 4295 11645 4307 11679
rect 4249 11639 4307 11645
rect 4342 11679 4400 11685
rect 4342 11645 4354 11679
rect 4388 11645 4400 11679
rect 4614 11676 4620 11688
rect 4575 11648 4620 11676
rect 4342 11639 4400 11645
rect 2041 11611 2099 11617
rect 2041 11577 2053 11611
rect 2087 11608 2099 11611
rect 2498 11608 2504 11620
rect 2087 11580 2504 11608
rect 2087 11577 2099 11580
rect 2041 11571 2099 11577
rect 2498 11568 2504 11580
rect 2556 11568 2562 11620
rect 2590 11568 2596 11620
rect 2648 11608 2654 11620
rect 2777 11611 2835 11617
rect 2777 11608 2789 11611
rect 2648 11580 2789 11608
rect 2648 11568 2654 11580
rect 2777 11577 2789 11580
rect 2823 11577 2835 11611
rect 2777 11571 2835 11577
rect 3697 11611 3755 11617
rect 3697 11577 3709 11611
rect 3743 11608 3755 11611
rect 4356 11608 4384 11639
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 4729 11685 4757 11784
rect 12713 11781 12725 11815
rect 12759 11812 12771 11815
rect 13262 11812 13268 11824
rect 12759 11784 13268 11812
rect 12759 11781 12771 11784
rect 12713 11775 12771 11781
rect 13262 11772 13268 11784
rect 13320 11772 13326 11824
rect 13464 11812 13492 11852
rect 13541 11849 13553 11883
rect 13587 11880 13599 11883
rect 13722 11880 13728 11892
rect 13587 11852 13728 11880
rect 13587 11849 13599 11852
rect 13541 11843 13599 11849
rect 13722 11840 13728 11852
rect 13780 11840 13786 11892
rect 15381 11883 15439 11889
rect 15381 11849 15393 11883
rect 15427 11880 15439 11883
rect 15746 11880 15752 11892
rect 15427 11852 15752 11880
rect 15427 11849 15439 11852
rect 15381 11843 15439 11849
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 15838 11840 15844 11892
rect 15896 11880 15902 11892
rect 16114 11880 16120 11892
rect 15896 11852 16120 11880
rect 15896 11840 15902 11852
rect 16114 11840 16120 11852
rect 16172 11840 16178 11892
rect 13814 11812 13820 11824
rect 13464 11784 13820 11812
rect 13814 11772 13820 11784
rect 13872 11772 13878 11824
rect 5074 11704 5080 11756
rect 5132 11744 5138 11756
rect 7374 11744 7380 11756
rect 5132 11716 7380 11744
rect 5132 11704 5138 11716
rect 5644 11685 5672 11716
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 12986 11744 12992 11756
rect 12947 11716 12992 11744
rect 12986 11704 12992 11716
rect 13044 11744 13050 11756
rect 13998 11744 14004 11756
rect 13044 11716 13768 11744
rect 13959 11716 14004 11744
rect 13044 11704 13050 11716
rect 4714 11679 4772 11685
rect 4714 11645 4726 11679
rect 4760 11645 4772 11679
rect 4714 11639 4772 11645
rect 5537 11679 5595 11685
rect 5537 11645 5549 11679
rect 5583 11645 5595 11679
rect 5537 11639 5595 11645
rect 5629 11679 5687 11685
rect 5629 11645 5641 11679
rect 5675 11645 5687 11679
rect 5902 11676 5908 11688
rect 5863 11648 5908 11676
rect 5629 11639 5687 11645
rect 3743 11580 4384 11608
rect 4525 11611 4583 11617
rect 3743 11577 3755 11580
rect 3697 11571 3755 11577
rect 4525 11577 4537 11611
rect 4571 11608 4583 11611
rect 5350 11608 5356 11620
rect 4571 11580 5356 11608
rect 4571 11577 4583 11580
rect 4525 11571 4583 11577
rect 5350 11568 5356 11580
rect 5408 11568 5414 11620
rect 5552 11608 5580 11639
rect 5902 11636 5908 11648
rect 5960 11636 5966 11688
rect 6730 11636 6736 11688
rect 6788 11676 6794 11688
rect 7006 11685 7012 11688
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6788 11648 6837 11676
rect 6788 11636 6794 11648
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 6973 11679 7012 11685
rect 6973 11645 6985 11679
rect 6973 11639 7012 11645
rect 7006 11636 7012 11639
rect 7064 11636 7070 11688
rect 7282 11636 7288 11688
rect 7340 11685 7346 11688
rect 7340 11676 7348 11685
rect 8478 11676 8484 11688
rect 7340 11648 7385 11676
rect 8439 11648 8484 11676
rect 7340 11639 7348 11648
rect 7340 11636 7346 11639
rect 8478 11636 8484 11648
rect 8536 11636 8542 11688
rect 10965 11679 11023 11685
rect 10965 11645 10977 11679
rect 11011 11676 11023 11679
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 11011 11648 12081 11676
rect 11011 11645 11023 11648
rect 10965 11639 11023 11645
rect 12069 11645 12081 11648
rect 12115 11676 12127 11679
rect 12158 11676 12164 11688
rect 12115 11648 12164 11676
rect 12115 11645 12127 11648
rect 12069 11639 12127 11645
rect 12158 11636 12164 11648
rect 12216 11636 12222 11688
rect 13078 11636 13084 11688
rect 13136 11676 13142 11688
rect 13740 11685 13768 11716
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 14108 11716 14964 11744
rect 13725 11679 13783 11685
rect 13136 11648 13181 11676
rect 13136 11636 13142 11648
rect 13725 11645 13737 11679
rect 13771 11645 13783 11679
rect 13725 11639 13783 11645
rect 5810 11608 5816 11620
rect 5552 11580 5816 11608
rect 5810 11568 5816 11580
rect 5868 11568 5874 11620
rect 6362 11568 6368 11620
rect 6420 11608 6426 11620
rect 7101 11611 7159 11617
rect 7101 11608 7113 11611
rect 6420 11580 7113 11608
rect 6420 11568 6426 11580
rect 7101 11577 7113 11580
rect 7147 11577 7159 11611
rect 7101 11571 7159 11577
rect 7193 11611 7251 11617
rect 7193 11577 7205 11611
rect 7239 11577 7251 11611
rect 8754 11608 8760 11620
rect 8715 11580 8760 11608
rect 7193 11571 7251 11577
rect 2133 11543 2191 11549
rect 2133 11509 2145 11543
rect 2179 11540 2191 11543
rect 2406 11540 2412 11552
rect 2179 11512 2412 11540
rect 2179 11509 2191 11512
rect 2133 11503 2191 11509
rect 2406 11500 2412 11512
rect 2464 11500 2470 11552
rect 4890 11540 4896 11552
rect 4851 11512 4896 11540
rect 4890 11500 4896 11512
rect 4948 11500 4954 11552
rect 6178 11500 6184 11552
rect 6236 11540 6242 11552
rect 7208 11540 7236 11571
rect 8754 11568 8760 11580
rect 8812 11568 8818 11620
rect 13740 11608 13768 11639
rect 13814 11636 13820 11688
rect 13872 11676 13878 11688
rect 14108 11685 14136 11716
rect 13909 11679 13967 11685
rect 13909 11676 13921 11679
rect 13872 11648 13921 11676
rect 13872 11636 13878 11648
rect 13909 11645 13921 11648
rect 13955 11645 13967 11679
rect 13909 11639 13967 11645
rect 14093 11679 14151 11685
rect 14093 11645 14105 11679
rect 14139 11645 14151 11679
rect 14274 11676 14280 11688
rect 14235 11648 14280 11676
rect 14093 11639 14151 11645
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 14936 11685 14964 11716
rect 15470 11704 15476 11756
rect 15528 11744 15534 11756
rect 15528 11716 16068 11744
rect 15528 11704 15534 11716
rect 15580 11685 15608 11716
rect 16040 11688 16068 11716
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11676 14979 11679
rect 15562 11679 15620 11685
rect 15562 11676 15574 11679
rect 14967 11648 15574 11676
rect 14967 11645 14979 11648
rect 14921 11639 14979 11645
rect 15562 11645 15574 11648
rect 15608 11645 15620 11679
rect 15930 11676 15936 11688
rect 15891 11648 15936 11676
rect 15562 11639 15620 11645
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 16022 11636 16028 11688
rect 16080 11676 16086 11688
rect 16080 11648 16125 11676
rect 16080 11636 16086 11648
rect 14829 11611 14887 11617
rect 14829 11608 14841 11611
rect 9982 11580 10824 11608
rect 13740 11580 14841 11608
rect 6236 11512 7236 11540
rect 7469 11543 7527 11549
rect 6236 11500 6242 11512
rect 7469 11509 7481 11543
rect 7515 11540 7527 11543
rect 8018 11540 8024 11552
rect 7515 11512 8024 11540
rect 7515 11509 7527 11512
rect 7469 11503 7527 11509
rect 8018 11500 8024 11512
rect 8076 11500 8082 11552
rect 10226 11540 10232 11552
rect 10187 11512 10232 11540
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 10796 11549 10824 11580
rect 14829 11577 14841 11580
rect 14875 11577 14887 11611
rect 14829 11571 14887 11577
rect 10781 11543 10839 11549
rect 10781 11509 10793 11543
rect 10827 11509 10839 11543
rect 10781 11503 10839 11509
rect 15565 11543 15623 11549
rect 15565 11509 15577 11543
rect 15611 11540 15623 11543
rect 15930 11540 15936 11552
rect 15611 11512 15936 11540
rect 15611 11509 15623 11512
rect 15565 11503 15623 11509
rect 15930 11500 15936 11512
rect 15988 11500 15994 11552
rect 1104 11450 17296 11472
rect 1104 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 6571 11450
rect 6623 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 11904 11450
rect 11956 11398 11968 11450
rect 12020 11398 17296 11450
rect 1104 11376 17296 11398
rect 2501 11339 2559 11345
rect 2501 11336 2513 11339
rect 1964 11308 2513 11336
rect 1964 11277 1992 11308
rect 2501 11305 2513 11308
rect 2547 11336 2559 11339
rect 2590 11336 2596 11348
rect 2547 11308 2596 11336
rect 2547 11305 2559 11308
rect 2501 11299 2559 11305
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 7466 11336 7472 11348
rect 7248 11308 7472 11336
rect 7248 11296 7254 11308
rect 7466 11296 7472 11308
rect 7524 11336 7530 11348
rect 8021 11339 8079 11345
rect 7524 11308 7972 11336
rect 7524 11296 7530 11308
rect 1949 11271 2007 11277
rect 1949 11237 1961 11271
rect 1995 11237 2007 11271
rect 1949 11231 2007 11237
rect 4154 11228 4160 11280
rect 4212 11268 4218 11280
rect 7742 11268 7748 11280
rect 4212 11240 5014 11268
rect 7484 11240 7748 11268
rect 4212 11228 4218 11240
rect 1489 11203 1547 11209
rect 1489 11169 1501 11203
rect 1535 11169 1547 11203
rect 2038 11200 2044 11212
rect 1999 11172 2044 11200
rect 1489 11163 1547 11169
rect 1504 11132 1532 11163
rect 2038 11160 2044 11172
rect 2096 11160 2102 11212
rect 2498 11200 2504 11212
rect 2459 11172 2504 11200
rect 2498 11160 2504 11172
rect 2556 11160 2562 11212
rect 7190 11200 7196 11212
rect 7151 11172 7196 11200
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11200 7343 11203
rect 7374 11200 7380 11212
rect 7331 11172 7380 11200
rect 7331 11169 7343 11172
rect 7285 11163 7343 11169
rect 7374 11160 7380 11172
rect 7432 11160 7438 11212
rect 2130 11132 2136 11144
rect 1504 11104 2136 11132
rect 2130 11092 2136 11104
rect 2188 11132 2194 11144
rect 2869 11135 2927 11141
rect 2869 11132 2881 11135
rect 2188 11104 2881 11132
rect 2188 11092 2194 11104
rect 2869 11101 2881 11104
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 4249 11135 4307 11141
rect 4249 11101 4261 11135
rect 4295 11101 4307 11135
rect 4522 11132 4528 11144
rect 4483 11104 4528 11132
rect 4249 11095 4307 11101
rect 4264 10996 4292 11095
rect 4522 11092 4528 11104
rect 4580 11092 4586 11144
rect 7484 11141 7512 11240
rect 7742 11228 7748 11240
rect 7800 11228 7806 11280
rect 7944 11268 7972 11308
rect 8021 11305 8033 11339
rect 8067 11336 8079 11339
rect 8754 11336 8760 11348
rect 8067 11308 8760 11336
rect 8067 11305 8079 11308
rect 8021 11299 8079 11305
rect 8754 11296 8760 11308
rect 8812 11296 8818 11348
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 11333 11339 11391 11345
rect 11333 11336 11345 11339
rect 10928 11308 11345 11336
rect 10928 11296 10934 11308
rect 11333 11305 11345 11308
rect 11379 11305 11391 11339
rect 11333 11299 11391 11305
rect 11606 11296 11612 11348
rect 11664 11336 11670 11348
rect 11664 11308 13400 11336
rect 11664 11296 11670 11308
rect 7944 11240 8340 11268
rect 7561 11203 7619 11209
rect 7561 11169 7573 11203
rect 7607 11169 7619 11203
rect 7561 11163 7619 11169
rect 7469 11135 7527 11141
rect 7469 11101 7481 11135
rect 7515 11101 7527 11135
rect 7576 11132 7604 11163
rect 8110 11160 8116 11212
rect 8168 11200 8174 11212
rect 8312 11209 8340 11240
rect 8478 11228 8484 11280
rect 8536 11268 8542 11280
rect 9950 11268 9956 11280
rect 8536 11240 9956 11268
rect 8536 11228 8542 11240
rect 9600 11209 9628 11240
rect 9950 11228 9956 11240
rect 10008 11228 10014 11280
rect 12066 11268 12072 11280
rect 11086 11240 12072 11268
rect 12066 11228 12072 11240
rect 12124 11228 12130 11280
rect 12802 11228 12808 11280
rect 12860 11228 12866 11280
rect 13372 11268 13400 11308
rect 15930 11296 15936 11348
rect 15988 11336 15994 11348
rect 16577 11339 16635 11345
rect 16577 11336 16589 11339
rect 15988 11308 16589 11336
rect 15988 11296 15994 11308
rect 16577 11305 16589 11308
rect 16623 11305 16635 11339
rect 16577 11299 16635 11305
rect 13817 11271 13875 11277
rect 13817 11268 13829 11271
rect 13372 11240 13829 11268
rect 13817 11237 13829 11240
rect 13863 11237 13875 11271
rect 15102 11268 15108 11280
rect 15063 11240 15108 11268
rect 13817 11231 13875 11237
rect 15102 11228 15108 11240
rect 15160 11228 15166 11280
rect 8205 11203 8263 11209
rect 8205 11200 8217 11203
rect 8168 11172 8217 11200
rect 8168 11160 8174 11172
rect 8205 11169 8217 11172
rect 8251 11169 8263 11203
rect 8205 11163 8263 11169
rect 8297 11203 8355 11209
rect 8297 11169 8309 11203
rect 8343 11169 8355 11203
rect 8297 11163 8355 11169
rect 9585 11203 9643 11209
rect 9585 11169 9597 11203
rect 9631 11169 9643 11203
rect 9585 11163 9643 11169
rect 14366 11160 14372 11212
rect 14424 11200 14430 11212
rect 14829 11203 14887 11209
rect 14829 11200 14841 11203
rect 14424 11172 14841 11200
rect 14424 11160 14430 11172
rect 14829 11169 14841 11172
rect 14875 11169 14887 11203
rect 14829 11163 14887 11169
rect 16206 11160 16212 11212
rect 16264 11160 16270 11212
rect 8018 11132 8024 11144
rect 7576 11104 7696 11132
rect 7979 11104 8024 11132
rect 7469 11095 7527 11101
rect 7009 11067 7067 11073
rect 7009 11033 7021 11067
rect 7055 11064 7067 11067
rect 7282 11064 7288 11076
rect 7055 11036 7288 11064
rect 7055 11033 7067 11036
rect 7009 11027 7067 11033
rect 7282 11024 7288 11036
rect 7340 11024 7346 11076
rect 4338 10996 4344 11008
rect 4251 10968 4344 10996
rect 4338 10956 4344 10968
rect 4396 10996 4402 11008
rect 4982 10996 4988 11008
rect 4396 10968 4988 10996
rect 4396 10956 4402 10968
rect 4982 10956 4988 10968
rect 5040 10956 5046 11008
rect 5810 10956 5816 11008
rect 5868 10996 5874 11008
rect 5997 10999 6055 11005
rect 5997 10996 6009 10999
rect 5868 10968 6009 10996
rect 5868 10956 5874 10968
rect 5997 10965 6009 10968
rect 6043 10965 6055 10999
rect 5997 10959 6055 10965
rect 6822 10956 6828 11008
rect 6880 10996 6886 11008
rect 7668 10996 7696 11104
rect 8018 11092 8024 11104
rect 8076 11092 8082 11144
rect 9858 11132 9864 11144
rect 9819 11104 9864 11132
rect 9858 11092 9864 11104
rect 9916 11092 9922 11144
rect 9950 11092 9956 11144
rect 10008 11132 10014 11144
rect 11793 11135 11851 11141
rect 11793 11132 11805 11135
rect 10008 11104 11805 11132
rect 10008 11092 10014 11104
rect 11793 11101 11805 11104
rect 11839 11101 11851 11135
rect 11793 11095 11851 11101
rect 12069 11135 12127 11141
rect 12069 11101 12081 11135
rect 12115 11132 12127 11135
rect 12618 11132 12624 11144
rect 12115 11104 12624 11132
rect 12115 11101 12127 11104
rect 12069 11095 12127 11101
rect 11808 11064 11836 11095
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 14366 11064 14372 11076
rect 11808 11036 11928 11064
rect 6880 10968 7696 10996
rect 11900 10996 11928 11036
rect 13096 11036 14372 11064
rect 13096 10996 13124 11036
rect 14366 11024 14372 11036
rect 14424 11024 14430 11076
rect 11900 10968 13124 10996
rect 6880 10956 6886 10968
rect 1104 10906 17296 10928
rect 1104 10854 3680 10906
rect 3732 10854 3744 10906
rect 3796 10854 3808 10906
rect 3860 10854 3872 10906
rect 3924 10854 9078 10906
rect 9130 10854 9142 10906
rect 9194 10854 9206 10906
rect 9258 10854 9270 10906
rect 9322 10854 14475 10906
rect 14527 10854 14539 10906
rect 14591 10854 14603 10906
rect 14655 10854 14667 10906
rect 14719 10854 17296 10906
rect 1104 10832 17296 10854
rect 2130 10792 2136 10804
rect 2091 10764 2136 10792
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 3789 10795 3847 10801
rect 3789 10761 3801 10795
rect 3835 10792 3847 10795
rect 4154 10792 4160 10804
rect 3835 10764 4160 10792
rect 3835 10761 3847 10764
rect 3789 10755 3847 10761
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 4433 10795 4491 10801
rect 4433 10761 4445 10795
rect 4479 10792 4491 10795
rect 4522 10792 4528 10804
rect 4479 10764 4528 10792
rect 4479 10761 4491 10764
rect 4433 10755 4491 10761
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 6178 10792 6184 10804
rect 5215 10764 6184 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 6178 10752 6184 10764
rect 6236 10752 6242 10804
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 7193 10795 7251 10801
rect 7193 10792 7205 10795
rect 7156 10764 7205 10792
rect 7156 10752 7162 10764
rect 7193 10761 7205 10764
rect 7239 10761 7251 10795
rect 7193 10755 7251 10761
rect 9858 10752 9864 10804
rect 9916 10792 9922 10804
rect 10597 10795 10655 10801
rect 10597 10792 10609 10795
rect 9916 10764 10609 10792
rect 9916 10752 9922 10764
rect 10597 10761 10609 10764
rect 10643 10761 10655 10795
rect 12066 10792 12072 10804
rect 12027 10764 12072 10792
rect 10597 10755 10655 10761
rect 12066 10752 12072 10764
rect 12124 10752 12130 10804
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 12897 10795 12955 10801
rect 12897 10792 12909 10795
rect 12860 10764 12909 10792
rect 12860 10752 12866 10764
rect 12897 10761 12909 10764
rect 12943 10761 12955 10795
rect 12897 10755 12955 10761
rect 2774 10684 2780 10736
rect 2832 10724 2838 10736
rect 8205 10727 8263 10733
rect 8205 10724 8217 10727
rect 2832 10696 2877 10724
rect 3160 10696 8217 10724
rect 2832 10684 2838 10696
rect 3160 10668 3188 10696
rect 8205 10693 8217 10696
rect 8251 10693 8263 10727
rect 8205 10687 8263 10693
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10656 1639 10659
rect 1946 10656 1952 10668
rect 1627 10628 1952 10656
rect 1627 10625 1639 10628
rect 1581 10619 1639 10625
rect 1946 10616 1952 10628
rect 2004 10616 2010 10668
rect 3142 10656 3148 10668
rect 3055 10628 3148 10656
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 4341 10659 4399 10665
rect 4341 10656 4353 10659
rect 3528 10628 4353 10656
rect 3050 10548 3056 10600
rect 3108 10588 3114 10600
rect 3528 10588 3556 10628
rect 4341 10625 4353 10628
rect 4387 10625 4399 10659
rect 4341 10619 4399 10625
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10656 4583 10659
rect 4890 10656 4896 10668
rect 4571 10628 4896 10656
rect 4571 10625 4583 10628
rect 4525 10619 4583 10625
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 6270 10656 6276 10668
rect 5592 10628 6276 10656
rect 5592 10616 5598 10628
rect 6270 10616 6276 10628
rect 6328 10616 6334 10668
rect 8662 10656 8668 10668
rect 8623 10628 8668 10656
rect 8662 10616 8668 10628
rect 8720 10616 8726 10668
rect 8754 10616 8760 10668
rect 8812 10656 8818 10668
rect 10962 10656 10968 10668
rect 8812 10628 8857 10656
rect 10796 10628 10968 10656
rect 8812 10616 8818 10628
rect 3108 10560 3556 10588
rect 3605 10591 3663 10597
rect 3108 10548 3114 10560
rect 3605 10557 3617 10591
rect 3651 10588 3663 10591
rect 3970 10588 3976 10600
rect 3651 10560 3976 10588
rect 3651 10557 3663 10560
rect 3605 10551 3663 10557
rect 1673 10523 1731 10529
rect 1673 10489 1685 10523
rect 1719 10520 1731 10523
rect 1719 10492 2912 10520
rect 1719 10489 1731 10492
rect 1673 10483 1731 10489
rect 1762 10412 1768 10464
rect 1820 10452 1826 10464
rect 1820 10424 1865 10452
rect 1820 10412 1826 10424
rect 2406 10412 2412 10464
rect 2464 10452 2470 10464
rect 2777 10455 2835 10461
rect 2777 10452 2789 10455
rect 2464 10424 2789 10452
rect 2464 10412 2470 10424
rect 2777 10421 2789 10424
rect 2823 10421 2835 10455
rect 2884 10452 2912 10492
rect 2958 10480 2964 10532
rect 3016 10520 3022 10532
rect 3620 10520 3648 10551
rect 3970 10548 3976 10560
rect 4028 10548 4034 10600
rect 4249 10591 4307 10597
rect 4249 10557 4261 10591
rect 4295 10557 4307 10591
rect 4249 10551 4307 10557
rect 5261 10591 5319 10597
rect 5261 10557 5273 10591
rect 5307 10588 5319 10591
rect 5626 10588 5632 10600
rect 5307 10560 5632 10588
rect 5307 10557 5319 10560
rect 5261 10551 5319 10557
rect 3016 10492 3648 10520
rect 4264 10520 4292 10551
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10588 5779 10591
rect 5810 10588 5816 10600
rect 5767 10560 5816 10588
rect 5767 10557 5779 10560
rect 5721 10551 5779 10557
rect 5810 10548 5816 10560
rect 5868 10548 5874 10600
rect 6730 10548 6736 10600
rect 6788 10588 6794 10600
rect 7101 10591 7159 10597
rect 7101 10588 7113 10591
rect 6788 10560 7113 10588
rect 6788 10548 6794 10560
rect 7101 10557 7113 10560
rect 7147 10557 7159 10591
rect 7101 10551 7159 10557
rect 9953 10591 10011 10597
rect 9953 10557 9965 10591
rect 9999 10588 10011 10591
rect 10226 10588 10232 10600
rect 9999 10560 10232 10588
rect 9999 10557 10011 10560
rect 9953 10551 10011 10557
rect 10226 10548 10232 10560
rect 10284 10588 10290 10600
rect 10796 10597 10824 10628
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 14090 10656 14096 10668
rect 14051 10628 14096 10656
rect 14090 10616 14096 10628
rect 14148 10616 14154 10668
rect 15841 10659 15899 10665
rect 15841 10625 15853 10659
rect 15887 10656 15899 10659
rect 16022 10656 16028 10668
rect 15887 10628 16028 10656
rect 15887 10625 15899 10628
rect 15841 10619 15899 10625
rect 16022 10616 16028 10628
rect 16080 10616 16086 10668
rect 10781 10591 10839 10597
rect 10284 10560 10732 10588
rect 10284 10548 10290 10560
rect 10594 10520 10600 10532
rect 4264 10492 5856 10520
rect 3016 10480 3022 10492
rect 5534 10452 5540 10464
rect 2884 10424 5540 10452
rect 2777 10415 2835 10421
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 5828 10461 5856 10492
rect 10060 10492 10600 10520
rect 5813 10455 5871 10461
rect 5813 10421 5825 10455
rect 5859 10452 5871 10455
rect 5902 10452 5908 10464
rect 5859 10424 5908 10452
rect 5859 10421 5871 10424
rect 5813 10415 5871 10421
rect 5902 10412 5908 10424
rect 5960 10452 5966 10464
rect 6178 10452 6184 10464
rect 5960 10424 6184 10452
rect 5960 10412 5966 10424
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 8570 10452 8576 10464
rect 8531 10424 8576 10452
rect 8570 10412 8576 10424
rect 8628 10412 8634 10464
rect 9674 10412 9680 10464
rect 9732 10452 9738 10464
rect 10060 10461 10088 10492
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 10045 10455 10103 10461
rect 10045 10452 10057 10455
rect 9732 10424 10057 10452
rect 9732 10412 9738 10424
rect 10045 10421 10057 10424
rect 10091 10421 10103 10455
rect 10704 10452 10732 10560
rect 10781 10557 10793 10591
rect 10827 10557 10839 10591
rect 10781 10551 10839 10557
rect 10870 10548 10876 10600
rect 10928 10588 10934 10600
rect 11146 10588 11152 10600
rect 10928 10560 10973 10588
rect 11107 10560 11152 10588
rect 10928 10548 10934 10560
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 12158 10548 12164 10600
rect 12216 10588 12222 10600
rect 12253 10591 12311 10597
rect 12253 10588 12265 10591
rect 12216 10560 12265 10588
rect 12216 10548 12222 10560
rect 12253 10557 12265 10560
rect 12299 10588 12311 10591
rect 13081 10591 13139 10597
rect 13081 10588 13093 10591
rect 12299 10560 13093 10588
rect 12299 10557 12311 10560
rect 12253 10551 12311 10557
rect 13081 10557 13093 10560
rect 13127 10588 13139 10591
rect 13354 10588 13360 10600
rect 13127 10560 13360 10588
rect 13127 10557 13139 10560
rect 13081 10551 13139 10557
rect 13354 10548 13360 10560
rect 13412 10548 13418 10600
rect 13817 10591 13875 10597
rect 13817 10557 13829 10591
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 10965 10523 11023 10529
rect 10965 10489 10977 10523
rect 11011 10520 11023 10523
rect 11606 10520 11612 10532
rect 11011 10492 11612 10520
rect 11011 10489 11023 10492
rect 10965 10483 11023 10489
rect 11606 10480 11612 10492
rect 11664 10480 11670 10532
rect 13832 10520 13860 10551
rect 14366 10520 14372 10532
rect 13832 10492 14372 10520
rect 14366 10480 14372 10492
rect 14424 10480 14430 10532
rect 14826 10480 14832 10532
rect 14884 10480 14890 10532
rect 12434 10452 12440 10464
rect 10704 10424 12440 10452
rect 10045 10415 10103 10421
rect 12434 10412 12440 10424
rect 12492 10412 12498 10464
rect 1104 10362 17296 10384
rect 1104 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 6571 10362
rect 6623 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 11904 10362
rect 11956 10310 11968 10362
rect 12020 10310 17296 10362
rect 1104 10288 17296 10310
rect 1486 10248 1492 10260
rect 1447 10220 1492 10248
rect 1486 10208 1492 10220
rect 1544 10208 1550 10260
rect 1762 10208 1768 10260
rect 1820 10248 1826 10260
rect 6089 10251 6147 10257
rect 6089 10248 6101 10251
rect 1820 10220 6101 10248
rect 1820 10208 1826 10220
rect 6089 10217 6101 10220
rect 6135 10217 6147 10251
rect 6089 10211 6147 10217
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 7834 10248 7840 10260
rect 7432 10220 7840 10248
rect 7432 10208 7438 10220
rect 7834 10208 7840 10220
rect 7892 10208 7898 10260
rect 8570 10208 8576 10260
rect 8628 10248 8634 10260
rect 9493 10251 9551 10257
rect 9493 10248 9505 10251
rect 8628 10220 9505 10248
rect 8628 10208 8634 10220
rect 9493 10217 9505 10220
rect 9539 10217 9551 10251
rect 9493 10211 9551 10217
rect 9858 10208 9864 10260
rect 9916 10248 9922 10260
rect 9916 10220 10916 10248
rect 9916 10208 9922 10220
rect 2406 10140 2412 10192
rect 2464 10180 2470 10192
rect 2685 10183 2743 10189
rect 2685 10180 2697 10183
rect 2464 10152 2697 10180
rect 2464 10140 2470 10152
rect 2685 10149 2697 10152
rect 2731 10149 2743 10183
rect 2685 10143 2743 10149
rect 4062 10140 4068 10192
rect 4120 10180 4126 10192
rect 4525 10183 4583 10189
rect 4525 10180 4537 10183
rect 4120 10152 4537 10180
rect 4120 10140 4126 10152
rect 4525 10149 4537 10152
rect 4571 10149 4583 10183
rect 4525 10143 4583 10149
rect 4893 10183 4951 10189
rect 4893 10149 4905 10183
rect 4939 10180 4951 10183
rect 9398 10180 9404 10192
rect 4939 10152 8064 10180
rect 4939 10149 4951 10152
rect 4893 10143 4951 10149
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10081 1639 10115
rect 1581 10075 1639 10081
rect 1596 10044 1624 10075
rect 2038 10072 2044 10124
rect 2096 10112 2102 10124
rect 2590 10112 2596 10124
rect 2096 10084 2596 10112
rect 2096 10072 2102 10084
rect 2590 10072 2596 10084
rect 2648 10072 2654 10124
rect 3142 10112 3148 10124
rect 3103 10084 3148 10112
rect 3142 10072 3148 10084
rect 3200 10072 3206 10124
rect 4709 10115 4767 10121
rect 4709 10081 4721 10115
rect 4755 10081 4767 10115
rect 4709 10075 4767 10081
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10112 5687 10115
rect 6273 10115 6331 10121
rect 6273 10112 6285 10115
rect 5675 10084 6285 10112
rect 5675 10081 5687 10084
rect 5629 10075 5687 10081
rect 6273 10081 6285 10084
rect 6319 10112 6331 10115
rect 7190 10112 7196 10124
rect 6319 10084 7196 10112
rect 6319 10081 6331 10084
rect 6273 10075 6331 10081
rect 2958 10044 2964 10056
rect 1596 10016 2964 10044
rect 2958 10004 2964 10016
rect 3016 10004 3022 10056
rect 4724 10044 4752 10075
rect 7190 10072 7196 10084
rect 7248 10072 7254 10124
rect 7374 10112 7380 10124
rect 7335 10084 7380 10112
rect 7374 10072 7380 10084
rect 7432 10072 7438 10124
rect 7466 10072 7472 10124
rect 7524 10112 7530 10124
rect 8036 10121 8064 10152
rect 8312 10152 9404 10180
rect 8312 10124 8340 10152
rect 9398 10140 9404 10152
rect 9456 10180 9462 10192
rect 9456 10152 10272 10180
rect 9456 10140 9462 10152
rect 8021 10115 8079 10121
rect 7524 10084 7569 10112
rect 7524 10072 7530 10084
rect 8021 10081 8033 10115
rect 8067 10081 8079 10115
rect 8021 10075 8079 10081
rect 8205 10115 8263 10121
rect 8205 10081 8217 10115
rect 8251 10112 8263 10115
rect 8294 10112 8300 10124
rect 8251 10084 8300 10112
rect 8251 10081 8263 10084
rect 8205 10075 8263 10081
rect 6178 10044 6184 10056
rect 4724 10016 6184 10044
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 6365 10047 6423 10053
rect 6365 10013 6377 10047
rect 6411 10013 6423 10047
rect 6365 10007 6423 10013
rect 6457 10047 6515 10053
rect 6457 10013 6469 10047
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 6822 10044 6828 10056
rect 6595 10016 6828 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 5626 9936 5632 9988
rect 5684 9976 5690 9988
rect 6380 9976 6408 10007
rect 5684 9948 6408 9976
rect 6472 9976 6500 10007
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 7650 10044 7656 10056
rect 6932 10016 7656 10044
rect 6932 9988 6960 10016
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 8036 10044 8064 10075
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 9769 10115 9827 10121
rect 9769 10081 9781 10115
rect 9815 10112 9827 10115
rect 9950 10112 9956 10124
rect 9815 10084 9956 10112
rect 9815 10081 9827 10084
rect 9769 10075 9827 10081
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 10244 10121 10272 10152
rect 10594 10140 10600 10192
rect 10652 10180 10658 10192
rect 10888 10189 10916 10220
rect 14826 10208 14832 10260
rect 14884 10248 14890 10260
rect 14921 10251 14979 10257
rect 14921 10248 14933 10251
rect 14884 10220 14933 10248
rect 14884 10208 14890 10220
rect 14921 10217 14933 10220
rect 14967 10217 14979 10251
rect 14921 10211 14979 10217
rect 15838 10208 15844 10260
rect 15896 10248 15902 10260
rect 15933 10251 15991 10257
rect 15933 10248 15945 10251
rect 15896 10220 15945 10248
rect 15896 10208 15902 10220
rect 15933 10217 15945 10220
rect 15979 10217 15991 10251
rect 15933 10211 15991 10217
rect 16206 10208 16212 10260
rect 16264 10248 16270 10260
rect 16393 10251 16451 10257
rect 16393 10248 16405 10251
rect 16264 10220 16405 10248
rect 16264 10208 16270 10220
rect 16393 10217 16405 10220
rect 16439 10217 16451 10251
rect 16393 10211 16451 10217
rect 10873 10183 10931 10189
rect 10652 10152 10824 10180
rect 10652 10140 10658 10152
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10081 10287 10115
rect 10229 10075 10287 10081
rect 10689 10115 10747 10121
rect 10689 10081 10701 10115
rect 10735 10081 10747 10115
rect 10796 10112 10824 10152
rect 10873 10149 10885 10183
rect 10919 10149 10931 10183
rect 11054 10180 11060 10192
rect 10967 10152 11060 10180
rect 10873 10143 10931 10149
rect 11054 10140 11060 10152
rect 11112 10180 11118 10192
rect 12253 10183 12311 10189
rect 12253 10180 12265 10183
rect 11112 10152 12265 10180
rect 11112 10140 11118 10152
rect 12253 10149 12265 10152
rect 12299 10149 12311 10183
rect 12253 10143 12311 10149
rect 11517 10115 11575 10121
rect 11517 10112 11529 10115
rect 10796 10084 11529 10112
rect 10689 10075 10747 10081
rect 11517 10081 11529 10084
rect 11563 10081 11575 10115
rect 11517 10075 11575 10081
rect 11701 10115 11759 10121
rect 11701 10081 11713 10115
rect 11747 10081 11759 10115
rect 12434 10112 12440 10124
rect 12395 10084 12440 10112
rect 11701 10075 11759 10081
rect 8938 10044 8944 10056
rect 8036 10016 8944 10044
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9861 10047 9919 10053
rect 9861 10013 9873 10047
rect 9907 10044 9919 10047
rect 10318 10044 10324 10056
rect 9907 10016 10324 10044
rect 9907 10013 9919 10016
rect 9861 10007 9919 10013
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 6914 9976 6920 9988
rect 6472 9948 6920 9976
rect 5684 9936 5690 9948
rect 5537 9911 5595 9917
rect 5537 9877 5549 9911
rect 5583 9908 5595 9911
rect 5810 9908 5816 9920
rect 5583 9880 5816 9908
rect 5583 9877 5595 9880
rect 5537 9871 5595 9877
rect 5810 9868 5816 9880
rect 5868 9908 5874 9920
rect 5994 9908 6000 9920
rect 5868 9880 6000 9908
rect 5868 9868 5874 9880
rect 5994 9868 6000 9880
rect 6052 9868 6058 9920
rect 6380 9908 6408 9948
rect 6914 9936 6920 9948
rect 6972 9936 6978 9988
rect 7285 9979 7343 9985
rect 7285 9945 7297 9979
rect 7331 9976 7343 9979
rect 8294 9976 8300 9988
rect 7331 9948 8300 9976
rect 7331 9945 7343 9948
rect 7285 9939 7343 9945
rect 8294 9936 8300 9948
rect 8352 9936 8358 9988
rect 9674 9936 9680 9988
rect 9732 9976 9738 9988
rect 9953 9979 10011 9985
rect 9953 9976 9965 9979
rect 9732 9948 9965 9976
rect 9732 9936 9738 9948
rect 9953 9945 9965 9948
rect 9999 9945 10011 9979
rect 9953 9939 10011 9945
rect 10134 9936 10140 9988
rect 10192 9976 10198 9988
rect 10704 9976 10732 10075
rect 10778 10004 10784 10056
rect 10836 10044 10842 10056
rect 11716 10044 11744 10075
rect 12434 10072 12440 10084
rect 12492 10072 12498 10124
rect 12894 10072 12900 10124
rect 12952 10112 12958 10124
rect 13265 10115 13323 10121
rect 13265 10112 13277 10115
rect 12952 10084 13277 10112
rect 12952 10072 12958 10084
rect 13265 10081 13277 10084
rect 13311 10081 13323 10115
rect 13265 10075 13323 10081
rect 13354 10072 13360 10124
rect 13412 10112 13418 10124
rect 14737 10115 14795 10121
rect 14737 10112 14749 10115
rect 13412 10084 14749 10112
rect 13412 10072 13418 10084
rect 14737 10081 14749 10084
rect 14783 10112 14795 10115
rect 16298 10112 16304 10124
rect 14783 10084 16304 10112
rect 14783 10081 14795 10084
rect 14737 10075 14795 10081
rect 16298 10072 16304 10084
rect 16356 10112 16362 10124
rect 16577 10115 16635 10121
rect 16577 10112 16589 10115
rect 16356 10084 16589 10112
rect 16356 10072 16362 10084
rect 16577 10081 16589 10084
rect 16623 10081 16635 10115
rect 16577 10075 16635 10081
rect 15562 10044 15568 10056
rect 10836 10016 11744 10044
rect 15523 10016 15568 10044
rect 10836 10004 10842 10016
rect 15562 10004 15568 10016
rect 15620 10004 15626 10056
rect 15930 9976 15936 9988
rect 10192 9948 10732 9976
rect 15891 9948 15936 9976
rect 10192 9936 10198 9948
rect 15930 9936 15936 9948
rect 15988 9936 15994 9988
rect 6730 9908 6736 9920
rect 6380 9880 6736 9908
rect 6730 9868 6736 9880
rect 6788 9868 6794 9920
rect 7098 9868 7104 9920
rect 7156 9908 7162 9920
rect 8021 9911 8079 9917
rect 8021 9908 8033 9911
rect 7156 9880 8033 9908
rect 7156 9868 7162 9880
rect 8021 9877 8033 9880
rect 8067 9908 8079 9911
rect 8110 9908 8116 9920
rect 8067 9880 8116 9908
rect 8067 9877 8079 9880
rect 8021 9871 8079 9877
rect 8110 9868 8116 9880
rect 8168 9868 8174 9920
rect 8389 9911 8447 9917
rect 8389 9877 8401 9911
rect 8435 9908 8447 9911
rect 9766 9908 9772 9920
rect 8435 9880 9772 9908
rect 8435 9877 8447 9880
rect 8389 9871 8447 9877
rect 9766 9868 9772 9880
rect 9824 9868 9830 9920
rect 10042 9908 10048 9920
rect 10003 9880 10048 9908
rect 10042 9868 10048 9880
rect 10100 9868 10106 9920
rect 11330 9868 11336 9920
rect 11388 9908 11394 9920
rect 11609 9911 11667 9917
rect 11609 9908 11621 9911
rect 11388 9880 11621 9908
rect 11388 9868 11394 9880
rect 11609 9877 11621 9880
rect 11655 9877 11667 9911
rect 12618 9908 12624 9920
rect 12579 9880 12624 9908
rect 11609 9871 11667 9877
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 13078 9908 13084 9920
rect 13039 9880 13084 9908
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 1104 9818 17296 9840
rect 1104 9766 3680 9818
rect 3732 9766 3744 9818
rect 3796 9766 3808 9818
rect 3860 9766 3872 9818
rect 3924 9766 9078 9818
rect 9130 9766 9142 9818
rect 9194 9766 9206 9818
rect 9258 9766 9270 9818
rect 9322 9766 14475 9818
rect 14527 9766 14539 9818
rect 14591 9766 14603 9818
rect 14655 9766 14667 9818
rect 14719 9766 17296 9818
rect 1104 9744 17296 9766
rect 3697 9707 3755 9713
rect 3697 9673 3709 9707
rect 3743 9704 3755 9707
rect 4062 9704 4068 9716
rect 3743 9676 4068 9704
rect 3743 9673 3755 9676
rect 3697 9667 3755 9673
rect 4062 9664 4068 9676
rect 4120 9664 4126 9716
rect 6730 9664 6736 9716
rect 6788 9704 6794 9716
rect 9309 9707 9367 9713
rect 9309 9704 9321 9707
rect 6788 9676 9321 9704
rect 6788 9664 6794 9676
rect 9309 9673 9321 9676
rect 9355 9704 9367 9707
rect 10042 9704 10048 9716
rect 9355 9676 10048 9704
rect 9355 9673 9367 9676
rect 9309 9667 9367 9673
rect 10042 9664 10048 9676
rect 10100 9664 10106 9716
rect 15562 9664 15568 9716
rect 15620 9704 15626 9716
rect 15657 9707 15715 9713
rect 15657 9704 15669 9707
rect 15620 9676 15669 9704
rect 15620 9664 15626 9676
rect 15657 9673 15669 9676
rect 15703 9673 15715 9707
rect 15657 9667 15715 9673
rect 15930 9664 15936 9716
rect 15988 9704 15994 9716
rect 16209 9707 16267 9713
rect 16209 9704 16221 9707
rect 15988 9676 16221 9704
rect 15988 9664 15994 9676
rect 16209 9673 16221 9676
rect 16255 9673 16267 9707
rect 16209 9667 16267 9673
rect 2590 9636 2596 9648
rect 2551 9608 2596 9636
rect 2590 9596 2596 9608
rect 2648 9596 2654 9648
rect 12250 9636 12256 9648
rect 2746 9608 12256 9636
rect 2038 9568 2044 9580
rect 1951 9540 2044 9568
rect 2038 9528 2044 9540
rect 2096 9568 2102 9580
rect 2406 9568 2412 9580
rect 2096 9540 2412 9568
rect 2096 9528 2102 9540
rect 2406 9528 2412 9540
rect 2464 9528 2470 9580
rect 2746 9512 2774 9608
rect 12250 9596 12256 9608
rect 12308 9596 12314 9648
rect 12728 9608 15056 9636
rect 12728 9580 12756 9608
rect 3510 9528 3516 9580
rect 3568 9568 3574 9580
rect 3568 9540 3740 9568
rect 3568 9528 3574 9540
rect 2682 9460 2688 9512
rect 2740 9472 2774 9512
rect 2740 9460 2746 9472
rect 3234 9460 3240 9512
rect 3292 9500 3298 9512
rect 3605 9503 3663 9509
rect 3605 9500 3617 9503
rect 3292 9472 3617 9500
rect 3292 9460 3298 9472
rect 3605 9469 3617 9472
rect 3651 9469 3663 9503
rect 3712 9500 3740 9540
rect 3970 9528 3976 9580
rect 4028 9568 4034 9580
rect 4249 9571 4307 9577
rect 4249 9568 4261 9571
rect 4028 9540 4261 9568
rect 4028 9528 4034 9540
rect 4249 9537 4261 9540
rect 4295 9537 4307 9571
rect 4249 9531 4307 9537
rect 4356 9540 5120 9568
rect 4356 9500 4384 9540
rect 4798 9500 4804 9512
rect 3712 9472 4384 9500
rect 4759 9472 4804 9500
rect 3605 9463 3663 9469
rect 1765 9435 1823 9441
rect 1765 9401 1777 9435
rect 1811 9432 1823 9435
rect 1811 9404 2176 9432
rect 1811 9401 1823 9404
rect 1765 9395 1823 9401
rect 1394 9364 1400 9376
rect 1355 9336 1400 9364
rect 1394 9324 1400 9336
rect 1452 9324 1458 9376
rect 1854 9364 1860 9376
rect 1815 9336 1860 9364
rect 1854 9324 1860 9336
rect 1912 9324 1918 9376
rect 2148 9364 2176 9404
rect 2222 9392 2228 9444
rect 2280 9432 2286 9444
rect 2777 9435 2835 9441
rect 2777 9432 2789 9435
rect 2280 9404 2789 9432
rect 2280 9392 2286 9404
rect 2777 9401 2789 9404
rect 2823 9401 2835 9435
rect 3620 9432 3648 9463
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 4982 9500 4988 9512
rect 4943 9472 4988 9500
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 5092 9500 5120 9540
rect 7466 9528 7472 9580
rect 7524 9568 7530 9580
rect 7742 9568 7748 9580
rect 7524 9540 7748 9568
rect 7524 9528 7530 9540
rect 7742 9528 7748 9540
rect 7800 9568 7806 9580
rect 9674 9568 9680 9580
rect 7800 9540 9680 9568
rect 7800 9528 7806 9540
rect 7926 9500 7932 9512
rect 5092 9472 7932 9500
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 8110 9500 8116 9512
rect 8071 9472 8116 9500
rect 8110 9460 8116 9472
rect 8168 9460 8174 9512
rect 8202 9460 8208 9512
rect 8260 9500 8266 9512
rect 8404 9509 8432 9540
rect 9674 9528 9680 9540
rect 9732 9528 9738 9580
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9568 10011 9571
rect 10134 9568 10140 9580
rect 9999 9540 10140 9568
rect 9999 9537 10011 9540
rect 9953 9531 10011 9537
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 10226 9528 10232 9580
rect 10284 9568 10290 9580
rect 10505 9571 10563 9577
rect 10505 9568 10517 9571
rect 10284 9540 10517 9568
rect 10284 9528 10290 9540
rect 10505 9537 10517 9540
rect 10551 9537 10563 9571
rect 10505 9531 10563 9537
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9568 10747 9571
rect 11054 9568 11060 9580
rect 10735 9540 11060 9568
rect 10735 9537 10747 9540
rect 10689 9531 10747 9537
rect 11054 9528 11060 9540
rect 11112 9528 11118 9580
rect 12710 9568 12716 9580
rect 12671 9540 12716 9568
rect 12710 9528 12716 9540
rect 12768 9528 12774 9580
rect 12897 9571 12955 9577
rect 12897 9537 12909 9571
rect 12943 9568 12955 9571
rect 13078 9568 13084 9580
rect 12943 9540 13084 9568
rect 12943 9537 12955 9540
rect 12897 9531 12955 9537
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 15028 9577 15056 9608
rect 15013 9571 15071 9577
rect 15013 9537 15025 9571
rect 15059 9537 15071 9571
rect 15013 9531 15071 9537
rect 8389 9503 8447 9509
rect 8260 9472 8305 9500
rect 8260 9460 8266 9472
rect 8389 9469 8401 9503
rect 8435 9469 8447 9503
rect 9582 9500 9588 9512
rect 8389 9463 8447 9469
rect 8496 9472 9588 9500
rect 5626 9432 5632 9444
rect 3620 9404 5632 9432
rect 2777 9395 2835 9401
rect 5626 9392 5632 9404
rect 5684 9432 5690 9444
rect 6825 9435 6883 9441
rect 6825 9432 6837 9435
rect 5684 9404 6837 9432
rect 5684 9392 5690 9404
rect 6825 9401 6837 9404
rect 6871 9401 6883 9435
rect 7006 9432 7012 9444
rect 6967 9404 7012 9432
rect 6825 9395 6883 9401
rect 7006 9392 7012 9404
rect 7064 9392 7070 9444
rect 7190 9432 7196 9444
rect 7103 9404 7196 9432
rect 7190 9392 7196 9404
rect 7248 9432 7254 9444
rect 8018 9432 8024 9444
rect 7248 9404 8024 9432
rect 7248 9392 7254 9404
rect 8018 9392 8024 9404
rect 8076 9392 8082 9444
rect 8220 9432 8248 9460
rect 8496 9432 8524 9472
rect 9582 9460 9588 9472
rect 9640 9460 9646 9512
rect 9766 9460 9772 9512
rect 9824 9500 9830 9512
rect 10778 9500 10784 9512
rect 9824 9472 10784 9500
rect 9824 9460 9830 9472
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 10870 9460 10876 9512
rect 10928 9500 10934 9512
rect 12161 9503 12219 9509
rect 12161 9500 12173 9503
rect 10928 9472 12173 9500
rect 10928 9460 10934 9472
rect 12161 9469 12173 9472
rect 12207 9469 12219 9503
rect 12161 9463 12219 9469
rect 12618 9460 12624 9512
rect 12676 9500 12682 9512
rect 12989 9503 13047 9509
rect 12989 9500 13001 9503
rect 12676 9472 13001 9500
rect 12676 9460 12682 9472
rect 12989 9469 13001 9472
rect 13035 9469 13047 9503
rect 12989 9463 13047 9469
rect 13262 9460 13268 9512
rect 13320 9500 13326 9512
rect 13817 9503 13875 9509
rect 13817 9500 13829 9503
rect 13320 9472 13829 9500
rect 13320 9460 13326 9472
rect 13817 9469 13829 9472
rect 13863 9469 13875 9503
rect 13817 9463 13875 9469
rect 14185 9503 14243 9509
rect 14185 9469 14197 9503
rect 14231 9500 14243 9503
rect 14734 9500 14740 9512
rect 14231 9472 14740 9500
rect 14231 9469 14243 9472
rect 14185 9463 14243 9469
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 15930 9460 15936 9512
rect 15988 9500 15994 9512
rect 16393 9503 16451 9509
rect 16393 9500 16405 9503
rect 15988 9472 16405 9500
rect 15988 9460 15994 9472
rect 16393 9469 16405 9472
rect 16439 9469 16451 9503
rect 16393 9463 16451 9469
rect 8220 9404 8524 9432
rect 9309 9435 9367 9441
rect 9309 9401 9321 9435
rect 9355 9432 9367 9435
rect 9401 9435 9459 9441
rect 9401 9432 9413 9435
rect 9355 9404 9413 9432
rect 9355 9401 9367 9404
rect 9309 9395 9367 9401
rect 9401 9401 9413 9404
rect 9447 9401 9459 9435
rect 9401 9395 9459 9401
rect 9490 9392 9496 9444
rect 9548 9432 9554 9444
rect 15289 9435 15347 9441
rect 15289 9432 15301 9435
rect 9548 9404 15301 9432
rect 9548 9392 9554 9404
rect 15289 9401 15301 9404
rect 15335 9401 15347 9435
rect 15289 9395 15347 9401
rect 3602 9364 3608 9376
rect 2148 9336 3608 9364
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 8570 9364 8576 9376
rect 8531 9336 8576 9364
rect 8570 9324 8576 9336
rect 8628 9324 8634 9376
rect 9030 9324 9036 9376
rect 9088 9364 9094 9376
rect 10318 9364 10324 9376
rect 9088 9336 10324 9364
rect 9088 9324 9094 9336
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 11146 9364 11152 9376
rect 11107 9336 11152 9364
rect 11146 9324 11152 9336
rect 11204 9324 11210 9376
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 11977 9367 12035 9373
rect 11977 9364 11989 9367
rect 11664 9336 11989 9364
rect 11664 9324 11670 9336
rect 11977 9333 11989 9336
rect 12023 9333 12035 9367
rect 13354 9364 13360 9376
rect 13315 9336 13360 9364
rect 11977 9327 12035 9333
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 13722 9324 13728 9376
rect 13780 9364 13786 9376
rect 14185 9367 14243 9373
rect 14185 9364 14197 9367
rect 13780 9336 14197 9364
rect 13780 9324 13786 9336
rect 14185 9333 14197 9336
rect 14231 9333 14243 9367
rect 15194 9364 15200 9376
rect 15155 9336 15200 9364
rect 14185 9327 14243 9333
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 1104 9274 17296 9296
rect 1104 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 6571 9274
rect 6623 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 11904 9274
rect 11956 9222 11968 9274
rect 12020 9222 17296 9274
rect 1104 9200 17296 9222
rect 2222 9160 2228 9172
rect 2183 9132 2228 9160
rect 2222 9120 2228 9132
rect 2280 9120 2286 9172
rect 3602 9120 3608 9172
rect 3660 9160 3666 9172
rect 5721 9163 5779 9169
rect 5721 9160 5733 9163
rect 3660 9132 5733 9160
rect 3660 9120 3666 9132
rect 5721 9129 5733 9132
rect 5767 9129 5779 9163
rect 5721 9123 5779 9129
rect 5810 9120 5816 9172
rect 5868 9160 5874 9172
rect 7098 9160 7104 9172
rect 5868 9132 7104 9160
rect 5868 9120 5874 9132
rect 7098 9120 7104 9132
rect 7156 9120 7162 9172
rect 8573 9163 8631 9169
rect 8573 9129 8585 9163
rect 8619 9160 8631 9163
rect 9490 9160 9496 9172
rect 8619 9132 9496 9160
rect 8619 9129 8631 9132
rect 8573 9123 8631 9129
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 12342 9160 12348 9172
rect 12303 9132 12348 9160
rect 12342 9120 12348 9132
rect 12400 9120 12406 9172
rect 12713 9163 12771 9169
rect 12713 9129 12725 9163
rect 12759 9160 12771 9163
rect 13262 9160 13268 9172
rect 12759 9132 13268 9160
rect 12759 9129 12771 9132
rect 12713 9123 12771 9129
rect 13262 9120 13268 9132
rect 13320 9120 13326 9172
rect 14734 9160 14740 9172
rect 14695 9132 14740 9160
rect 14734 9120 14740 9132
rect 14792 9120 14798 9172
rect 1854 9052 1860 9104
rect 1912 9092 1918 9104
rect 5077 9095 5135 9101
rect 1912 9064 2774 9092
rect 1912 9052 1918 9064
rect 2746 9024 2774 9064
rect 5077 9061 5089 9095
rect 5123 9092 5135 9095
rect 11333 9095 11391 9101
rect 5123 9064 10916 9092
rect 5123 9061 5135 9064
rect 5077 9055 5135 9061
rect 5810 9024 5816 9036
rect 2746 8996 5816 9024
rect 5810 8984 5816 8996
rect 5868 8984 5874 9036
rect 5905 9027 5963 9033
rect 5905 8993 5917 9027
rect 5951 8993 5963 9027
rect 5905 8987 5963 8993
rect 6089 9027 6147 9033
rect 6089 8993 6101 9027
rect 6135 9024 6147 9027
rect 6362 9024 6368 9036
rect 6135 8996 6368 9024
rect 6135 8993 6147 8996
rect 6089 8987 6147 8993
rect 1394 8916 1400 8968
rect 1452 8956 1458 8968
rect 1857 8959 1915 8965
rect 1857 8956 1869 8959
rect 1452 8928 1869 8956
rect 1452 8916 1458 8928
rect 1857 8925 1869 8928
rect 1903 8925 1915 8959
rect 1857 8919 1915 8925
rect 2774 8916 2780 8968
rect 2832 8956 2838 8968
rect 3142 8956 3148 8968
rect 2832 8928 2877 8956
rect 3103 8928 3148 8956
rect 2832 8916 2838 8928
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 5074 8956 5080 8968
rect 5035 8928 5080 8956
rect 5074 8916 5080 8928
rect 5132 8916 5138 8968
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 5350 8956 5356 8968
rect 5215 8928 5356 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 2225 8891 2283 8897
rect 2225 8857 2237 8891
rect 2271 8888 2283 8891
rect 2498 8888 2504 8900
rect 2271 8860 2504 8888
rect 2271 8857 2283 8860
rect 2225 8851 2283 8857
rect 2498 8848 2504 8860
rect 2556 8848 2562 8900
rect 5920 8888 5948 8987
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 6730 9024 6736 9036
rect 6691 8996 6736 9024
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 6914 9024 6920 9036
rect 6875 8996 6920 9024
rect 6914 8984 6920 8996
rect 6972 8984 6978 9036
rect 7098 8984 7104 9036
rect 7156 9024 7162 9036
rect 7377 9027 7435 9033
rect 7377 9024 7389 9027
rect 7156 8996 7389 9024
rect 7156 8984 7162 8996
rect 7377 8993 7389 8996
rect 7423 8993 7435 9027
rect 7377 8987 7435 8993
rect 8294 8984 8300 9036
rect 8352 9024 8358 9036
rect 8389 9027 8447 9033
rect 8389 9024 8401 9027
rect 8352 8996 8401 9024
rect 8352 8984 8358 8996
rect 8389 8993 8401 8996
rect 8435 8993 8447 9027
rect 8389 8987 8447 8993
rect 9398 8984 9404 9036
rect 9456 9024 9462 9036
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 9456 8996 9505 9024
rect 9456 8984 9462 8996
rect 9493 8993 9505 8996
rect 9539 8993 9551 9027
rect 9493 8987 9551 8993
rect 9674 8984 9680 9036
rect 9732 9024 9738 9036
rect 9769 9027 9827 9033
rect 9769 9024 9781 9027
rect 9732 8996 9781 9024
rect 9732 8984 9738 8996
rect 9769 8993 9781 8996
rect 9815 8993 9827 9027
rect 9950 9024 9956 9036
rect 9911 8996 9956 9024
rect 9769 8987 9827 8993
rect 9950 8984 9956 8996
rect 10008 8984 10014 9036
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8956 7711 8959
rect 7926 8956 7932 8968
rect 7699 8928 7932 8956
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 8018 8916 8024 8968
rect 8076 8956 8082 8968
rect 8113 8959 8171 8965
rect 8113 8956 8125 8959
rect 8076 8928 8125 8956
rect 8076 8916 8082 8928
rect 8113 8925 8125 8928
rect 8159 8925 8171 8959
rect 8113 8919 8171 8925
rect 6546 8888 6552 8900
rect 5828 8860 6408 8888
rect 6507 8860 6552 8888
rect 2590 8780 2596 8832
rect 2648 8820 2654 8832
rect 2777 8823 2835 8829
rect 2777 8820 2789 8823
rect 2648 8792 2789 8820
rect 2648 8780 2654 8792
rect 2777 8789 2789 8792
rect 2823 8789 2835 8823
rect 4614 8820 4620 8832
rect 4575 8792 4620 8820
rect 2777 8783 2835 8789
rect 4614 8780 4620 8792
rect 4672 8780 4678 8832
rect 5442 8780 5448 8832
rect 5500 8820 5506 8832
rect 5828 8820 5856 8860
rect 5994 8820 6000 8832
rect 5500 8792 5856 8820
rect 5955 8792 6000 8820
rect 5500 8780 5506 8792
rect 5994 8780 6000 8792
rect 6052 8780 6058 8832
rect 6380 8820 6408 8860
rect 6546 8848 6552 8860
rect 6604 8848 6610 8900
rect 6730 8820 6736 8832
rect 6380 8792 6736 8820
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 7466 8820 7472 8832
rect 7427 8792 7472 8820
rect 7466 8780 7472 8792
rect 7524 8780 7530 8832
rect 7561 8823 7619 8829
rect 7561 8789 7573 8823
rect 7607 8820 7619 8823
rect 8018 8820 8024 8832
rect 7607 8792 8024 8820
rect 7607 8789 7619 8792
rect 7561 8783 7619 8789
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 8128 8820 8156 8919
rect 8478 8916 8484 8968
rect 8536 8956 8542 8968
rect 10888 8956 10916 9064
rect 11333 9061 11345 9095
rect 11379 9092 11391 9095
rect 13538 9092 13544 9104
rect 11379 9064 13544 9092
rect 11379 9061 11391 9064
rect 11333 9055 11391 9061
rect 13538 9052 13544 9064
rect 13596 9052 13602 9104
rect 13722 9092 13728 9104
rect 13683 9064 13728 9092
rect 13722 9052 13728 9064
rect 13780 9052 13786 9104
rect 15838 9052 15844 9104
rect 15896 9092 15902 9104
rect 15933 9095 15991 9101
rect 15933 9092 15945 9095
rect 15896 9064 15945 9092
rect 15896 9052 15902 9064
rect 15933 9061 15945 9064
rect 15979 9061 15991 9095
rect 15933 9055 15991 9061
rect 12250 9024 12256 9036
rect 12211 8996 12256 9024
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 13262 9024 13268 9036
rect 13223 8996 13268 9024
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 13817 9027 13875 9033
rect 13817 8993 13829 9027
rect 13863 9024 13875 9027
rect 14921 9027 14979 9033
rect 14921 9024 14933 9027
rect 13863 8996 14933 9024
rect 13863 8993 13875 8996
rect 13817 8987 13875 8993
rect 14921 8993 14933 8996
rect 14967 9024 14979 9027
rect 15010 9024 15016 9036
rect 14967 8996 15016 9024
rect 14967 8993 14979 8996
rect 14921 8987 14979 8993
rect 15010 8984 15016 8996
rect 15068 8984 15074 9036
rect 15473 9027 15531 9033
rect 15473 8993 15485 9027
rect 15519 9024 15531 9027
rect 15562 9024 15568 9036
rect 15519 8996 15568 9024
rect 15519 8993 15531 8996
rect 15473 8987 15531 8993
rect 15562 8984 15568 8996
rect 15620 8984 15626 9036
rect 16025 9027 16083 9033
rect 16025 9024 16037 9027
rect 15948 8996 16037 9024
rect 15948 8968 15976 8996
rect 16025 8993 16037 8996
rect 16071 8993 16083 9027
rect 16025 8987 16083 8993
rect 11330 8956 11336 8968
rect 8536 8928 9996 8956
rect 10888 8928 11192 8956
rect 11291 8928 11336 8956
rect 8536 8916 8542 8928
rect 8205 8891 8263 8897
rect 8205 8857 8217 8891
rect 8251 8888 8263 8891
rect 8662 8888 8668 8900
rect 8251 8860 8668 8888
rect 8251 8857 8263 8860
rect 8205 8851 8263 8857
rect 8662 8848 8668 8860
rect 8720 8848 8726 8900
rect 9858 8888 9864 8900
rect 8772 8860 9864 8888
rect 8772 8820 8800 8860
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 8128 8792 8800 8820
rect 9677 8823 9735 8829
rect 9677 8789 9689 8823
rect 9723 8820 9735 8823
rect 9766 8820 9772 8832
rect 9723 8792 9772 8820
rect 9723 8789 9735 8792
rect 9677 8783 9735 8789
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 9968 8820 9996 8928
rect 10229 8891 10287 8897
rect 10229 8857 10241 8891
rect 10275 8888 10287 8891
rect 10778 8888 10784 8900
rect 10275 8860 10784 8888
rect 10275 8857 10287 8860
rect 10229 8851 10287 8857
rect 10778 8848 10784 8860
rect 10836 8848 10842 8900
rect 11164 8888 11192 8928
rect 11330 8916 11336 8928
rect 11388 8916 11394 8968
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8956 11483 8959
rect 12161 8959 12219 8965
rect 12161 8956 12173 8959
rect 11471 8928 12173 8956
rect 11471 8925 11483 8928
rect 11425 8919 11483 8925
rect 12161 8925 12173 8928
rect 12207 8956 12219 8959
rect 12710 8956 12716 8968
rect 12207 8928 12716 8956
rect 12207 8925 12219 8928
rect 12161 8919 12219 8925
rect 12710 8916 12716 8928
rect 12768 8956 12774 8968
rect 12986 8956 12992 8968
rect 12768 8928 12992 8956
rect 12768 8916 12774 8928
rect 12986 8916 12992 8928
rect 13044 8916 13050 8968
rect 15930 8916 15936 8968
rect 15988 8916 15994 8968
rect 14366 8888 14372 8900
rect 11164 8860 14372 8888
rect 14366 8848 14372 8860
rect 14424 8848 14430 8900
rect 10873 8823 10931 8829
rect 10873 8820 10885 8823
rect 9968 8792 10885 8820
rect 10873 8789 10885 8792
rect 10919 8789 10931 8823
rect 10873 8783 10931 8789
rect 1104 8730 17296 8752
rect 1104 8678 3680 8730
rect 3732 8678 3744 8730
rect 3796 8678 3808 8730
rect 3860 8678 3872 8730
rect 3924 8678 9078 8730
rect 9130 8678 9142 8730
rect 9194 8678 9206 8730
rect 9258 8678 9270 8730
rect 9322 8678 14475 8730
rect 14527 8678 14539 8730
rect 14591 8678 14603 8730
rect 14655 8678 14667 8730
rect 14719 8678 17296 8730
rect 1104 8656 17296 8678
rect 2590 8616 2596 8628
rect 2551 8588 2596 8616
rect 2590 8576 2596 8588
rect 2648 8576 2654 8628
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 5353 8619 5411 8625
rect 5353 8616 5365 8619
rect 5132 8588 5365 8616
rect 5132 8576 5138 8588
rect 5353 8585 5365 8588
rect 5399 8585 5411 8619
rect 5353 8579 5411 8585
rect 5810 8576 5816 8628
rect 5868 8616 5874 8628
rect 7834 8616 7840 8628
rect 5868 8588 7840 8616
rect 5868 8576 5874 8588
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 8018 8576 8024 8628
rect 8076 8616 8082 8628
rect 8076 8588 10456 8616
rect 8076 8576 8082 8588
rect 8294 8548 8300 8560
rect 4724 8520 8300 8548
rect 4430 8440 4436 8492
rect 4488 8480 4494 8492
rect 4617 8483 4675 8489
rect 4617 8480 4629 8483
rect 4488 8452 4629 8480
rect 4488 8440 4494 8452
rect 4617 8449 4629 8452
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 2593 8415 2651 8421
rect 2593 8381 2605 8415
rect 2639 8412 2651 8415
rect 2682 8412 2688 8424
rect 2639 8384 2688 8412
rect 2639 8381 2651 8384
rect 2593 8375 2651 8381
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 3142 8412 3148 8424
rect 3103 8384 3148 8412
rect 3142 8372 3148 8384
rect 3200 8372 3206 8424
rect 4525 8415 4583 8421
rect 4525 8381 4537 8415
rect 4571 8412 4583 8415
rect 4724 8412 4752 8520
rect 8294 8508 8300 8520
rect 8352 8508 8358 8560
rect 9582 8508 9588 8560
rect 9640 8548 9646 8560
rect 10428 8548 10456 8588
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 12437 8619 12495 8625
rect 12437 8616 12449 8619
rect 10560 8588 12449 8616
rect 10560 8576 10566 8588
rect 12437 8585 12449 8588
rect 12483 8585 12495 8619
rect 12437 8579 12495 8585
rect 13538 8576 13544 8628
rect 13596 8616 13602 8628
rect 14645 8619 14703 8625
rect 14645 8616 14657 8619
rect 13596 8588 14657 8616
rect 13596 8576 13602 8588
rect 14645 8585 14657 8588
rect 14691 8585 14703 8619
rect 14645 8579 14703 8585
rect 11238 8548 11244 8560
rect 9640 8520 10272 8548
rect 10428 8520 11244 8548
rect 9640 8508 9646 8520
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8480 4859 8483
rect 4982 8480 4988 8492
rect 4847 8452 4988 8480
rect 4847 8449 4859 8452
rect 4801 8443 4859 8449
rect 4982 8440 4988 8452
rect 5040 8480 5046 8492
rect 5350 8480 5356 8492
rect 5040 8452 5356 8480
rect 5040 8440 5046 8452
rect 5350 8440 5356 8452
rect 5408 8440 5414 8492
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 5813 8483 5871 8489
rect 5684 8452 5729 8480
rect 5684 8440 5690 8452
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 5902 8480 5908 8492
rect 5859 8452 5908 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 5902 8440 5908 8452
rect 5960 8480 5966 8492
rect 6546 8480 6552 8492
rect 5960 8452 6552 8480
rect 5960 8440 5966 8452
rect 6546 8440 6552 8452
rect 6604 8440 6610 8492
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 7653 8483 7711 8489
rect 7653 8480 7665 8483
rect 7156 8452 7665 8480
rect 7156 8440 7162 8452
rect 7653 8449 7665 8452
rect 7699 8480 7711 8483
rect 8110 8480 8116 8492
rect 7699 8452 8116 8480
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 8110 8440 8116 8452
rect 8168 8440 8174 8492
rect 9398 8480 9404 8492
rect 8588 8452 9404 8480
rect 5534 8412 5540 8424
rect 4571 8384 4752 8412
rect 5495 8384 5540 8412
rect 4571 8381 4583 8384
rect 4525 8375 4583 8381
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 5721 8415 5779 8421
rect 5721 8381 5733 8415
rect 5767 8412 5779 8415
rect 5994 8412 6000 8424
rect 5767 8384 6000 8412
rect 5767 8381 5779 8384
rect 5721 8375 5779 8381
rect 5994 8372 6000 8384
rect 6052 8412 6058 8424
rect 7006 8412 7012 8424
rect 6052 8384 7012 8412
rect 6052 8372 6058 8384
rect 7006 8372 7012 8384
rect 7064 8412 7070 8424
rect 7282 8412 7288 8424
rect 7064 8384 7288 8412
rect 7064 8372 7070 8384
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 7466 8412 7472 8424
rect 7427 8384 7472 8412
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8381 7619 8415
rect 7742 8412 7748 8424
rect 7703 8384 7748 8412
rect 7561 8375 7619 8381
rect 1394 8344 1400 8356
rect 1355 8316 1400 8344
rect 1394 8304 1400 8316
rect 1452 8304 1458 8356
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 2130 8344 2136 8356
rect 1627 8316 2136 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 2130 8304 2136 8316
rect 2188 8304 2194 8356
rect 6362 8304 6368 8356
rect 6420 8304 6426 8356
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7576 8344 7604 8375
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 7834 8372 7840 8424
rect 7892 8412 7898 8424
rect 8588 8412 8616 8452
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 9766 8440 9772 8492
rect 9824 8480 9830 8492
rect 10045 8483 10103 8489
rect 10045 8480 10057 8483
rect 9824 8452 10057 8480
rect 9824 8440 9830 8452
rect 10045 8449 10057 8452
rect 10091 8449 10103 8483
rect 10045 8443 10103 8449
rect 8754 8412 8760 8424
rect 7892 8384 8616 8412
rect 8715 8384 8760 8412
rect 7892 8372 7898 8384
rect 8754 8372 8760 8384
rect 8812 8412 8818 8424
rect 9674 8412 9680 8424
rect 8812 8384 9680 8412
rect 8812 8372 8818 8384
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 10244 8421 10272 8520
rect 11238 8508 11244 8520
rect 11296 8508 11302 8560
rect 11422 8508 11428 8560
rect 11480 8548 11486 8560
rect 11793 8551 11851 8557
rect 11793 8548 11805 8551
rect 11480 8520 11805 8548
rect 11480 8508 11486 8520
rect 11793 8517 11805 8520
rect 11839 8517 11851 8551
rect 11793 8511 11851 8517
rect 10318 8440 10324 8492
rect 10376 8480 10382 8492
rect 12986 8480 12992 8492
rect 10376 8452 10421 8480
rect 12947 8452 12992 8480
rect 10376 8440 10382 8452
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 14274 8480 14280 8492
rect 13648 8452 14280 8480
rect 10229 8415 10287 8421
rect 10229 8381 10241 8415
rect 10275 8381 10287 8415
rect 10229 8375 10287 8381
rect 10413 8415 10471 8421
rect 10413 8381 10425 8415
rect 10459 8381 10471 8415
rect 10413 8375 10471 8381
rect 10505 8415 10563 8421
rect 10505 8381 10517 8415
rect 10551 8381 10563 8415
rect 10505 8375 10563 8381
rect 11977 8415 12035 8421
rect 11977 8381 11989 8415
rect 12023 8412 12035 8415
rect 13648 8412 13676 8452
rect 14274 8440 14280 8452
rect 14332 8440 14338 8492
rect 12023 8384 13676 8412
rect 12023 8381 12035 8384
rect 11977 8375 12035 8381
rect 8202 8344 8208 8356
rect 6972 8316 8208 8344
rect 6972 8304 6978 8316
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 9401 8347 9459 8353
rect 9401 8313 9413 8347
rect 9447 8313 9459 8347
rect 9401 8307 9459 8313
rect 4157 8279 4215 8285
rect 4157 8245 4169 8279
rect 4203 8276 4215 8279
rect 4246 8276 4252 8288
rect 4203 8248 4252 8276
rect 4203 8245 4215 8248
rect 4157 8239 4215 8245
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 5994 8236 6000 8288
rect 6052 8276 6058 8288
rect 6380 8276 6408 8304
rect 7926 8276 7932 8288
rect 6052 8248 6408 8276
rect 7887 8248 7932 8276
rect 6052 8236 6058 8248
rect 7926 8236 7932 8248
rect 7984 8236 7990 8288
rect 8018 8236 8024 8288
rect 8076 8276 8082 8288
rect 9416 8276 9444 8307
rect 9858 8304 9864 8356
rect 9916 8344 9922 8356
rect 10042 8344 10048 8356
rect 9916 8316 10048 8344
rect 9916 8304 9922 8316
rect 10042 8304 10048 8316
rect 10100 8344 10106 8356
rect 10419 8344 10447 8375
rect 10100 8316 10447 8344
rect 10100 8304 10106 8316
rect 8076 8248 9444 8276
rect 8076 8236 8082 8248
rect 10226 8236 10232 8288
rect 10284 8276 10290 8288
rect 10520 8276 10548 8375
rect 13722 8372 13728 8424
rect 13780 8412 13786 8424
rect 14093 8415 14151 8421
rect 14093 8412 14105 8415
rect 13780 8384 14105 8412
rect 13780 8372 13786 8384
rect 14093 8381 14105 8384
rect 14139 8381 14151 8415
rect 14826 8412 14832 8424
rect 14787 8384 14832 8412
rect 14093 8375 14151 8381
rect 14826 8372 14832 8384
rect 14884 8372 14890 8424
rect 15286 8412 15292 8424
rect 15247 8384 15292 8412
rect 15286 8372 15292 8384
rect 15344 8372 15350 8424
rect 15657 8415 15715 8421
rect 15657 8381 15669 8415
rect 15703 8412 15715 8415
rect 16209 8415 16267 8421
rect 16209 8412 16221 8415
rect 15703 8384 16221 8412
rect 15703 8381 15715 8384
rect 15657 8375 15715 8381
rect 16209 8381 16221 8384
rect 16255 8381 16267 8415
rect 16209 8375 16267 8381
rect 12897 8347 12955 8353
rect 12897 8313 12909 8347
rect 12943 8344 12955 8347
rect 13906 8344 13912 8356
rect 12943 8316 13768 8344
rect 13867 8316 13912 8344
rect 12943 8313 12955 8316
rect 12897 8307 12955 8313
rect 12802 8276 12808 8288
rect 10284 8248 10548 8276
rect 12763 8248 12808 8276
rect 10284 8236 10290 8248
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 13740 8276 13768 8316
rect 13906 8304 13912 8316
rect 13964 8304 13970 8356
rect 15838 8304 15844 8356
rect 15896 8344 15902 8356
rect 16117 8347 16175 8353
rect 16117 8344 16129 8347
rect 15896 8316 16129 8344
rect 15896 8304 15902 8316
rect 16117 8313 16129 8316
rect 16163 8313 16175 8347
rect 16117 8307 16175 8313
rect 15102 8276 15108 8288
rect 13740 8248 15108 8276
rect 15102 8236 15108 8248
rect 15160 8236 15166 8288
rect 15654 8276 15660 8288
rect 15615 8248 15660 8276
rect 15654 8236 15660 8248
rect 15712 8236 15718 8288
rect 1104 8186 17296 8208
rect 1104 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 6571 8186
rect 6623 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 11904 8186
rect 11956 8134 11968 8186
rect 12020 8134 17296 8186
rect 1104 8112 17296 8134
rect 2590 8032 2596 8084
rect 2648 8072 2654 8084
rect 2685 8075 2743 8081
rect 2685 8072 2697 8075
rect 2648 8044 2697 8072
rect 2648 8032 2654 8044
rect 2685 8041 2697 8044
rect 2731 8041 2743 8075
rect 2685 8035 2743 8041
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 3145 8075 3203 8081
rect 3145 8072 3157 8075
rect 2832 8044 3157 8072
rect 2832 8032 2838 8044
rect 3145 8041 3157 8044
rect 3191 8041 3203 8075
rect 3145 8035 3203 8041
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 5813 8075 5871 8081
rect 5813 8072 5825 8075
rect 5776 8044 5825 8072
rect 5776 8032 5782 8044
rect 5813 8041 5825 8044
rect 5859 8041 5871 8075
rect 5813 8035 5871 8041
rect 7190 8032 7196 8084
rect 7248 8072 7254 8084
rect 11425 8075 11483 8081
rect 7248 8044 9996 8072
rect 7248 8032 7254 8044
rect 1857 8007 1915 8013
rect 1857 7973 1869 8007
rect 1903 8004 1915 8007
rect 2222 8004 2228 8016
rect 1903 7976 2228 8004
rect 1903 7973 1915 7976
rect 1857 7967 1915 7973
rect 2222 7964 2228 7976
rect 2280 7964 2286 8016
rect 2498 8004 2504 8016
rect 2459 7976 2504 8004
rect 2498 7964 2504 7976
rect 2556 7964 2562 8016
rect 6178 7964 6184 8016
rect 6236 8004 6242 8016
rect 6236 7976 7236 8004
rect 6236 7964 6242 7976
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1486 7936 1492 7948
rect 1443 7908 1492 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1486 7896 1492 7908
rect 1544 7896 1550 7948
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7936 2007 7939
rect 2682 7936 2688 7948
rect 1995 7908 2688 7936
rect 1995 7905 2007 7908
rect 1949 7899 2007 7905
rect 2682 7896 2688 7908
rect 2740 7936 2746 7948
rect 3329 7939 3387 7945
rect 3329 7936 3341 7939
rect 2740 7908 3341 7936
rect 2740 7896 2746 7908
rect 3329 7905 3341 7908
rect 3375 7905 3387 7939
rect 3329 7899 3387 7905
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 4249 7939 4307 7945
rect 4249 7936 4261 7939
rect 4212 7908 4261 7936
rect 4212 7896 4218 7908
rect 4249 7905 4261 7908
rect 4295 7905 4307 7939
rect 4249 7899 4307 7905
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7936 5227 7939
rect 5534 7936 5540 7948
rect 5215 7908 5540 7936
rect 5215 7905 5227 7908
rect 5169 7899 5227 7905
rect 5534 7896 5540 7908
rect 5592 7936 5598 7948
rect 5810 7936 5816 7948
rect 5592 7908 5816 7936
rect 5592 7896 5598 7908
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 7098 7936 7104 7948
rect 7059 7908 7104 7936
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 7208 7936 7236 7976
rect 7374 7964 7380 8016
rect 7432 8004 7438 8016
rect 8389 8007 8447 8013
rect 8389 8004 8401 8007
rect 7432 7976 8401 8004
rect 7432 7964 7438 7976
rect 8389 7973 8401 7976
rect 8435 7973 8447 8007
rect 8389 7967 8447 7973
rect 8662 7964 8668 8016
rect 8720 8004 8726 8016
rect 9645 8007 9703 8013
rect 9645 8004 9657 8007
rect 8720 7976 9657 8004
rect 8720 7964 8726 7976
rect 9645 7973 9657 7976
rect 9691 7973 9703 8007
rect 9645 7967 9703 7973
rect 9861 8007 9919 8013
rect 9861 7973 9873 8007
rect 9907 7973 9919 8007
rect 9968 8004 9996 8044
rect 11425 8041 11437 8075
rect 11471 8072 11483 8075
rect 12342 8072 12348 8084
rect 11471 8044 12348 8072
rect 11471 8041 11483 8044
rect 11425 8035 11483 8041
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 12713 8075 12771 8081
rect 12713 8041 12725 8075
rect 12759 8072 12771 8075
rect 12802 8072 12808 8084
rect 12759 8044 12808 8072
rect 12759 8041 12771 8044
rect 12713 8035 12771 8041
rect 12802 8032 12808 8044
rect 12860 8032 12866 8084
rect 14366 8032 14372 8084
rect 14424 8072 14430 8084
rect 14645 8075 14703 8081
rect 14645 8072 14657 8075
rect 14424 8044 14657 8072
rect 14424 8032 14430 8044
rect 14645 8041 14657 8044
rect 14691 8041 14703 8075
rect 14645 8035 14703 8041
rect 15194 8032 15200 8084
rect 15252 8072 15258 8084
rect 16393 8075 16451 8081
rect 16393 8072 16405 8075
rect 15252 8044 16405 8072
rect 15252 8032 15258 8044
rect 16393 8041 16405 8044
rect 16439 8041 16451 8075
rect 16393 8035 16451 8041
rect 9968 7976 15056 8004
rect 9861 7967 9919 7973
rect 7561 7939 7619 7945
rect 7561 7936 7573 7939
rect 7208 7908 7573 7936
rect 7561 7905 7573 7908
rect 7607 7936 7619 7939
rect 8481 7939 8539 7945
rect 7607 7908 7788 7936
rect 7607 7905 7619 7908
rect 7561 7899 7619 7905
rect 5350 7828 5356 7880
rect 5408 7868 5414 7880
rect 5718 7868 5724 7880
rect 5408 7840 5724 7868
rect 5408 7828 5414 7840
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 5902 7868 5908 7880
rect 5863 7840 5908 7868
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 7466 7868 7472 7880
rect 6871 7840 7472 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 1946 7760 1952 7812
rect 2004 7800 2010 7812
rect 2222 7800 2228 7812
rect 2004 7772 2228 7800
rect 2004 7760 2010 7772
rect 2222 7760 2228 7772
rect 2280 7760 2286 7812
rect 5077 7803 5135 7809
rect 5077 7769 5089 7803
rect 5123 7800 5135 7803
rect 6840 7800 6868 7831
rect 7466 7828 7472 7840
rect 7524 7868 7530 7880
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 7524 7840 7665 7868
rect 7524 7828 7530 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 5123 7772 6868 7800
rect 7009 7803 7067 7809
rect 5123 7769 5135 7772
rect 5077 7763 5135 7769
rect 7009 7769 7021 7803
rect 7055 7800 7067 7803
rect 7760 7800 7788 7908
rect 8481 7905 8493 7939
rect 8527 7936 8539 7939
rect 8941 7939 8999 7945
rect 8941 7936 8953 7939
rect 8527 7908 8953 7936
rect 8527 7905 8539 7908
rect 8481 7899 8539 7905
rect 8941 7905 8953 7908
rect 8987 7905 8999 7939
rect 9876 7936 9904 7967
rect 10226 7936 10232 7948
rect 9876 7908 10232 7936
rect 8941 7899 8999 7905
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 10321 7939 10379 7945
rect 10321 7905 10333 7939
rect 10367 7905 10379 7939
rect 11146 7936 11152 7948
rect 11107 7908 11152 7936
rect 10321 7899 10379 7905
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7868 7895 7871
rect 7926 7868 7932 7880
rect 7883 7840 7932 7868
rect 7883 7837 7895 7840
rect 7837 7831 7895 7837
rect 7926 7828 7932 7840
rect 7984 7868 7990 7880
rect 10336 7868 10364 7899
rect 11146 7896 11152 7908
rect 11204 7896 11210 7948
rect 11241 7939 11299 7945
rect 11241 7905 11253 7939
rect 11287 7936 11299 7939
rect 11330 7936 11336 7948
rect 11287 7908 11336 7936
rect 11287 7905 11299 7908
rect 11241 7899 11299 7905
rect 11330 7896 11336 7908
rect 11388 7896 11394 7948
rect 11514 7896 11520 7948
rect 11572 7936 11578 7948
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 11572 7908 12081 7936
rect 11572 7896 11578 7908
rect 12069 7905 12081 7908
rect 12115 7905 12127 7939
rect 12529 7939 12587 7945
rect 12529 7936 12541 7939
rect 12069 7899 12127 7905
rect 12406 7908 12541 7936
rect 7984 7840 10364 7868
rect 7984 7828 7990 7840
rect 10410 7828 10416 7880
rect 10468 7868 10474 7880
rect 12406 7868 12434 7908
rect 12529 7905 12541 7908
rect 12575 7936 12587 7939
rect 12710 7936 12716 7948
rect 12575 7908 12716 7936
rect 12575 7905 12587 7908
rect 12529 7899 12587 7905
rect 12710 7896 12716 7908
rect 12768 7896 12774 7948
rect 13170 7936 13176 7948
rect 13131 7908 13176 7936
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 13725 7939 13783 7945
rect 13725 7905 13737 7939
rect 13771 7905 13783 7939
rect 13725 7899 13783 7905
rect 14829 7939 14887 7945
rect 14829 7905 14841 7939
rect 14875 7936 14887 7939
rect 14918 7936 14924 7948
rect 14875 7908 14924 7936
rect 14875 7905 14887 7908
rect 14829 7899 14887 7905
rect 10468 7840 12434 7868
rect 13740 7868 13768 7899
rect 14918 7896 14924 7908
rect 14976 7896 14982 7948
rect 15028 7936 15056 7976
rect 15654 7964 15660 8016
rect 15712 8004 15718 8016
rect 15749 8007 15807 8013
rect 15749 8004 15761 8007
rect 15712 7976 15761 8004
rect 15712 7964 15718 7976
rect 15749 7973 15761 7976
rect 15795 7973 15807 8007
rect 15749 7967 15807 7973
rect 15286 7945 15292 7948
rect 15277 7939 15292 7945
rect 15277 7936 15289 7939
rect 15028 7908 15289 7936
rect 15277 7905 15289 7908
rect 15277 7899 15292 7905
rect 15286 7896 15292 7899
rect 15344 7896 15350 7948
rect 15838 7936 15844 7948
rect 15799 7908 15844 7936
rect 15838 7896 15844 7908
rect 15896 7896 15902 7948
rect 16577 7939 16635 7945
rect 16577 7905 16589 7939
rect 16623 7936 16635 7939
rect 17034 7936 17040 7948
rect 16623 7908 17040 7936
rect 16623 7905 16635 7908
rect 16577 7899 16635 7905
rect 17034 7896 17040 7908
rect 17092 7896 17098 7948
rect 15010 7868 15016 7880
rect 13740 7840 15016 7868
rect 10468 7828 10474 7840
rect 15010 7828 15016 7840
rect 15068 7828 15074 7880
rect 7055 7772 7788 7800
rect 9493 7803 9551 7809
rect 7055 7769 7067 7772
rect 7009 7763 7067 7769
rect 9493 7769 9505 7803
rect 9539 7800 9551 7803
rect 9539 7772 9812 7800
rect 9539 7769 9551 7772
rect 9493 7763 9551 7769
rect 4338 7732 4344 7744
rect 4299 7704 4344 7732
rect 4338 7692 4344 7704
rect 4396 7692 4402 7744
rect 6273 7735 6331 7741
rect 6273 7701 6285 7735
rect 6319 7732 6331 7735
rect 6730 7732 6736 7744
rect 6319 7704 6736 7732
rect 6319 7701 6331 7704
rect 6273 7695 6331 7701
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 6914 7732 6920 7744
rect 6875 7704 6920 7732
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 7742 7732 7748 7744
rect 7703 7704 7748 7732
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 8941 7735 8999 7741
rect 8941 7701 8953 7735
rect 8987 7732 8999 7735
rect 9582 7732 9588 7744
rect 8987 7704 9588 7732
rect 8987 7701 8999 7704
rect 8941 7695 8999 7701
rect 9582 7692 9588 7704
rect 9640 7732 9646 7744
rect 9677 7735 9735 7741
rect 9677 7732 9689 7735
rect 9640 7704 9689 7732
rect 9640 7692 9646 7704
rect 9677 7701 9689 7704
rect 9723 7701 9735 7735
rect 9784 7732 9812 7772
rect 9858 7760 9864 7812
rect 9916 7800 9922 7812
rect 11885 7803 11943 7809
rect 11885 7800 11897 7803
rect 9916 7772 11897 7800
rect 9916 7760 9922 7772
rect 11885 7769 11897 7772
rect 11931 7769 11943 7803
rect 11885 7763 11943 7769
rect 9950 7732 9956 7744
rect 9784 7704 9956 7732
rect 9677 7695 9735 7701
rect 9950 7692 9956 7704
rect 10008 7692 10014 7744
rect 10042 7692 10048 7744
rect 10100 7732 10106 7744
rect 10413 7735 10471 7741
rect 10413 7732 10425 7735
rect 10100 7704 10425 7732
rect 10100 7692 10106 7704
rect 10413 7701 10425 7704
rect 10459 7701 10471 7735
rect 13722 7732 13728 7744
rect 13683 7704 13728 7732
rect 10413 7695 10471 7701
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 1104 7642 17296 7664
rect 1104 7590 3680 7642
rect 3732 7590 3744 7642
rect 3796 7590 3808 7642
rect 3860 7590 3872 7642
rect 3924 7590 9078 7642
rect 9130 7590 9142 7642
rect 9194 7590 9206 7642
rect 9258 7590 9270 7642
rect 9322 7590 14475 7642
rect 14527 7590 14539 7642
rect 14591 7590 14603 7642
rect 14655 7590 14667 7642
rect 14719 7590 17296 7642
rect 1104 7568 17296 7590
rect 2501 7531 2559 7537
rect 2501 7497 2513 7531
rect 2547 7528 2559 7531
rect 2682 7528 2688 7540
rect 2547 7500 2688 7528
rect 2547 7497 2559 7500
rect 2501 7491 2559 7497
rect 2682 7488 2688 7500
rect 2740 7488 2746 7540
rect 5902 7488 5908 7540
rect 5960 7528 5966 7540
rect 6825 7531 6883 7537
rect 6825 7528 6837 7531
rect 5960 7500 6837 7528
rect 5960 7488 5966 7500
rect 6825 7497 6837 7500
rect 6871 7497 6883 7531
rect 6825 7491 6883 7497
rect 8481 7531 8539 7537
rect 8481 7497 8493 7531
rect 8527 7528 8539 7531
rect 8662 7528 8668 7540
rect 8527 7500 8668 7528
rect 8527 7497 8539 7500
rect 8481 7491 8539 7497
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 10134 7528 10140 7540
rect 9640 7500 10140 7528
rect 9640 7488 9646 7500
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 10321 7531 10379 7537
rect 10321 7497 10333 7531
rect 10367 7528 10379 7531
rect 12250 7528 12256 7540
rect 10367 7500 12256 7528
rect 10367 7497 10379 7500
rect 10321 7491 10379 7497
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 13170 7488 13176 7540
rect 13228 7528 13234 7540
rect 13265 7531 13323 7537
rect 13265 7528 13277 7531
rect 13228 7500 13277 7528
rect 13228 7488 13234 7500
rect 13265 7497 13277 7500
rect 13311 7497 13323 7531
rect 13265 7491 13323 7497
rect 15102 7488 15108 7540
rect 15160 7528 15166 7540
rect 16209 7531 16267 7537
rect 16209 7528 16221 7531
rect 15160 7500 16221 7528
rect 15160 7488 15166 7500
rect 16209 7497 16221 7500
rect 16255 7497 16267 7531
rect 16209 7491 16267 7497
rect 4246 7420 4252 7472
rect 4304 7420 4310 7472
rect 5813 7463 5871 7469
rect 5813 7429 5825 7463
rect 5859 7460 5871 7463
rect 7190 7460 7196 7472
rect 5859 7432 7196 7460
rect 5859 7429 5871 7432
rect 5813 7423 5871 7429
rect 7190 7420 7196 7432
rect 7248 7420 7254 7472
rect 10042 7460 10048 7472
rect 7300 7432 10048 7460
rect 4264 7392 4292 7420
rect 3712 7364 4292 7392
rect 5445 7395 5503 7401
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 2866 7324 2872 7336
rect 1443 7296 2872 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 2866 7284 2872 7296
rect 2924 7284 2930 7336
rect 3050 7284 3056 7336
rect 3108 7324 3114 7336
rect 3712 7333 3740 7364
rect 5445 7361 5457 7395
rect 5491 7392 5503 7395
rect 5534 7392 5540 7404
rect 5491 7364 5540 7392
rect 5491 7361 5503 7364
rect 5445 7355 5503 7361
rect 5534 7352 5540 7364
rect 5592 7392 5598 7404
rect 7300 7401 7328 7432
rect 10042 7420 10048 7432
rect 10100 7420 10106 7472
rect 12158 7460 12164 7472
rect 12119 7432 12164 7460
rect 12158 7420 12164 7432
rect 12216 7420 12222 7472
rect 15010 7460 15016 7472
rect 14971 7432 15016 7460
rect 15010 7420 15016 7432
rect 15068 7420 15074 7472
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 5592 7364 7021 7392
rect 5592 7352 5598 7364
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 7742 7352 7748 7404
rect 7800 7392 7806 7404
rect 12529 7395 12587 7401
rect 12529 7392 12541 7395
rect 7800 7364 12541 7392
rect 7800 7352 7806 7364
rect 12529 7361 12541 7364
rect 12575 7361 12587 7395
rect 12986 7392 12992 7404
rect 12529 7355 12587 7361
rect 12820 7364 12992 7392
rect 3697 7327 3755 7333
rect 3697 7324 3709 7327
rect 3108 7296 3709 7324
rect 3108 7284 3114 7296
rect 3697 7293 3709 7296
rect 3743 7293 3755 7327
rect 3697 7287 3755 7293
rect 4249 7327 4307 7333
rect 4249 7293 4261 7327
rect 4295 7324 4307 7327
rect 4706 7324 4712 7336
rect 4295 7296 4712 7324
rect 4295 7293 4307 7296
rect 4249 7287 4307 7293
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 5626 7284 5632 7336
rect 5684 7324 5690 7336
rect 5902 7324 5908 7336
rect 5684 7296 5908 7324
rect 5684 7284 5690 7296
rect 5902 7284 5908 7296
rect 5960 7324 5966 7336
rect 7101 7327 7159 7333
rect 7101 7324 7113 7327
rect 5960 7296 7113 7324
rect 5960 7284 5966 7296
rect 7101 7293 7113 7296
rect 7147 7293 7159 7327
rect 7101 7287 7159 7293
rect 7193 7327 7251 7333
rect 7193 7293 7205 7327
rect 7239 7324 7251 7327
rect 7374 7324 7380 7336
rect 7239 7296 7380 7324
rect 7239 7293 7251 7296
rect 7193 7287 7251 7293
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 8294 7324 8300 7336
rect 8255 7296 8300 7324
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 8570 7284 8576 7336
rect 8628 7324 8634 7336
rect 8628 7296 8673 7324
rect 8628 7284 8634 7296
rect 8938 7284 8944 7336
rect 8996 7324 9002 7336
rect 9033 7327 9091 7333
rect 9033 7324 9045 7327
rect 8996 7296 9045 7324
rect 8996 7284 9002 7296
rect 9033 7293 9045 7296
rect 9079 7293 9091 7327
rect 10873 7327 10931 7333
rect 9033 7287 9091 7293
rect 9140 7296 10180 7324
rect 2593 7259 2651 7265
rect 2593 7225 2605 7259
rect 2639 7256 2651 7259
rect 2682 7256 2688 7268
rect 2639 7228 2688 7256
rect 2639 7225 2651 7228
rect 2593 7219 2651 7225
rect 2682 7216 2688 7228
rect 2740 7216 2746 7268
rect 3326 7216 3332 7268
rect 3384 7256 3390 7268
rect 4154 7256 4160 7268
rect 3384 7228 4160 7256
rect 3384 7216 3390 7228
rect 4154 7216 4160 7228
rect 4212 7216 4218 7268
rect 5261 7259 5319 7265
rect 5261 7225 5273 7259
rect 5307 7256 5319 7259
rect 5718 7256 5724 7268
rect 5307 7228 5724 7256
rect 5307 7225 5319 7228
rect 5261 7219 5319 7225
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 2498 7148 2504 7200
rect 2556 7188 2562 7200
rect 5276 7188 5304 7219
rect 5718 7216 5724 7228
rect 5776 7216 5782 7268
rect 9140 7256 9168 7296
rect 8036 7228 9168 7256
rect 2556 7160 5304 7188
rect 5353 7191 5411 7197
rect 2556 7148 2562 7160
rect 5353 7157 5365 7191
rect 5399 7188 5411 7191
rect 8036 7188 8064 7228
rect 9674 7216 9680 7268
rect 9732 7256 9738 7268
rect 9769 7259 9827 7265
rect 9769 7256 9781 7259
rect 9732 7228 9781 7256
rect 9732 7216 9738 7228
rect 9769 7225 9781 7228
rect 9815 7225 9827 7259
rect 9769 7219 9827 7225
rect 5399 7160 8064 7188
rect 8113 7191 8171 7197
rect 5399 7157 5411 7160
rect 5353 7151 5411 7157
rect 8113 7157 8125 7191
rect 8159 7188 8171 7191
rect 8202 7188 8208 7200
rect 8159 7160 8208 7188
rect 8159 7157 8171 7160
rect 8113 7151 8171 7157
rect 8202 7148 8208 7160
rect 8260 7148 8266 7200
rect 8570 7148 8576 7200
rect 8628 7188 8634 7200
rect 9125 7191 9183 7197
rect 9125 7188 9137 7191
rect 8628 7160 9137 7188
rect 8628 7148 8634 7160
rect 9125 7157 9137 7160
rect 9171 7157 9183 7191
rect 9784 7188 9812 7219
rect 9858 7216 9864 7268
rect 9916 7256 9922 7268
rect 10042 7256 10048 7268
rect 9916 7228 9961 7256
rect 10003 7228 10048 7256
rect 9916 7216 9922 7228
rect 10042 7216 10048 7228
rect 10100 7216 10106 7268
rect 10152 7256 10180 7296
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 10962 7324 10968 7336
rect 10919 7296 10968 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 12820 7268 12848 7364
rect 12986 7352 12992 7364
rect 13044 7392 13050 7404
rect 13817 7395 13875 7401
rect 13817 7392 13829 7395
rect 13044 7364 13829 7392
rect 13044 7352 13050 7364
rect 13817 7361 13829 7364
rect 13863 7361 13875 7395
rect 13817 7355 13875 7361
rect 15197 7327 15255 7333
rect 15197 7293 15209 7327
rect 15243 7324 15255 7327
rect 15654 7324 15660 7336
rect 15243 7296 15660 7324
rect 15243 7293 15255 7296
rect 15197 7287 15255 7293
rect 15654 7284 15660 7296
rect 15712 7284 15718 7336
rect 16390 7324 16396 7336
rect 16351 7296 16396 7324
rect 16390 7284 16396 7296
rect 16448 7284 16454 7336
rect 12526 7256 12532 7268
rect 10152 7228 12532 7256
rect 12526 7216 12532 7228
rect 12584 7216 12590 7268
rect 12713 7259 12771 7265
rect 12713 7225 12725 7259
rect 12759 7256 12771 7259
rect 12802 7256 12808 7268
rect 12759 7228 12808 7256
rect 12759 7225 12771 7228
rect 12713 7219 12771 7225
rect 12802 7216 12808 7228
rect 12860 7216 12866 7268
rect 14918 7256 14924 7268
rect 13464 7228 14924 7256
rect 10318 7188 10324 7200
rect 9784 7160 10324 7188
rect 9125 7151 9183 7157
rect 10318 7148 10324 7160
rect 10376 7148 10382 7200
rect 11054 7188 11060 7200
rect 11015 7160 11060 7188
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 12621 7191 12679 7197
rect 12621 7157 12633 7191
rect 12667 7188 12679 7191
rect 13464 7188 13492 7228
rect 14918 7216 14924 7228
rect 14976 7216 14982 7268
rect 13630 7188 13636 7200
rect 12667 7160 13492 7188
rect 13591 7160 13636 7188
rect 12667 7157 12679 7160
rect 12621 7151 12679 7157
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 13725 7191 13783 7197
rect 13725 7157 13737 7191
rect 13771 7188 13783 7191
rect 14182 7188 14188 7200
rect 13771 7160 14188 7188
rect 13771 7157 13783 7160
rect 13725 7151 13783 7157
rect 14182 7148 14188 7160
rect 14240 7148 14246 7200
rect 1104 7098 17296 7120
rect 1104 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 6571 7098
rect 6623 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 11904 7098
rect 11956 7046 11968 7098
rect 12020 7046 17296 7098
rect 1104 7024 17296 7046
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 2041 6987 2099 6993
rect 2041 6984 2053 6987
rect 1636 6956 2053 6984
rect 1636 6944 1642 6956
rect 2041 6953 2053 6956
rect 2087 6953 2099 6987
rect 5442 6984 5448 6996
rect 2041 6947 2099 6953
rect 2746 6956 5448 6984
rect 1949 6919 2007 6925
rect 1949 6885 1961 6919
rect 1995 6916 2007 6919
rect 2746 6916 2774 6956
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 8202 6984 8208 6996
rect 8163 6956 8208 6984
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 8294 6944 8300 6996
rect 8352 6984 8358 6996
rect 8938 6984 8944 6996
rect 8352 6956 8944 6984
rect 8352 6944 8358 6956
rect 8938 6944 8944 6956
rect 8996 6944 9002 6996
rect 10318 6944 10324 6996
rect 10376 6984 10382 6996
rect 12802 6984 12808 6996
rect 10376 6956 12808 6984
rect 10376 6944 10382 6956
rect 12802 6944 12808 6956
rect 12860 6944 12866 6996
rect 12897 6987 12955 6993
rect 12897 6953 12909 6987
rect 12943 6984 12955 6987
rect 13630 6984 13636 6996
rect 12943 6956 13636 6984
rect 12943 6953 12955 6956
rect 12897 6947 12955 6953
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 13722 6944 13728 6996
rect 13780 6984 13786 6996
rect 13817 6987 13875 6993
rect 13817 6984 13829 6987
rect 13780 6956 13829 6984
rect 13780 6944 13786 6956
rect 13817 6953 13829 6956
rect 13863 6953 13875 6987
rect 13817 6947 13875 6953
rect 15838 6944 15844 6996
rect 15896 6984 15902 6996
rect 16393 6987 16451 6993
rect 16393 6984 16405 6987
rect 15896 6956 16405 6984
rect 15896 6944 15902 6956
rect 16393 6953 16405 6956
rect 16439 6953 16451 6987
rect 16393 6947 16451 6953
rect 6914 6916 6920 6928
rect 1995 6888 2774 6916
rect 6564 6888 6920 6916
rect 1995 6885 2007 6888
rect 1949 6879 2007 6885
rect 2961 6851 3019 6857
rect 2961 6817 2973 6851
rect 3007 6848 3019 6851
rect 3050 6848 3056 6860
rect 3007 6820 3056 6848
rect 3007 6817 3019 6820
rect 2961 6811 3019 6817
rect 3050 6808 3056 6820
rect 3108 6808 3114 6860
rect 4614 6808 4620 6860
rect 4672 6848 4678 6860
rect 4801 6851 4859 6857
rect 4801 6848 4813 6851
rect 4672 6820 4813 6848
rect 4672 6808 4678 6820
rect 4801 6817 4813 6820
rect 4847 6817 4859 6851
rect 4801 6811 4859 6817
rect 5721 6851 5779 6857
rect 5721 6817 5733 6851
rect 5767 6817 5779 6851
rect 5902 6848 5908 6860
rect 5863 6820 5908 6848
rect 5721 6811 5779 6817
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2498 6780 2504 6792
rect 2271 6752 2504 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2498 6740 2504 6752
rect 2556 6740 2562 6792
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6780 3387 6783
rect 4062 6780 4068 6792
rect 3375 6752 4068 6780
rect 3375 6749 3387 6752
rect 3329 6743 3387 6749
rect 4062 6740 4068 6752
rect 4120 6740 4126 6792
rect 4246 6780 4252 6792
rect 4207 6752 4252 6780
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 5736 6780 5764 6811
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 5994 6808 6000 6860
rect 6052 6848 6058 6860
rect 6052 6820 6097 6848
rect 6052 6808 6058 6820
rect 6564 6780 6592 6888
rect 6914 6876 6920 6888
rect 6972 6876 6978 6928
rect 8478 6916 8484 6928
rect 7300 6888 8484 6916
rect 6641 6851 6699 6857
rect 6641 6817 6653 6851
rect 6687 6848 6699 6851
rect 7300 6848 7328 6888
rect 8478 6876 8484 6888
rect 8536 6876 8542 6928
rect 12158 6916 12164 6928
rect 11256 6888 12164 6916
rect 6687 6820 7328 6848
rect 7377 6851 7435 6857
rect 6687 6817 6699 6820
rect 6641 6811 6699 6817
rect 7377 6817 7389 6851
rect 7423 6848 7435 6851
rect 7558 6848 7564 6860
rect 7423 6820 7564 6848
rect 7423 6817 7435 6820
rect 7377 6811 7435 6817
rect 7558 6808 7564 6820
rect 7616 6808 7622 6860
rect 9674 6848 9680 6860
rect 9635 6820 9680 6848
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 10870 6848 10876 6860
rect 9784 6820 10876 6848
rect 8018 6780 8024 6792
rect 5736 6752 6592 6780
rect 7979 6752 8024 6780
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 1946 6672 1952 6724
rect 2004 6712 2010 6724
rect 4338 6712 4344 6724
rect 2004 6684 3464 6712
rect 4299 6684 4344 6712
rect 2004 6672 2010 6684
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 3326 6644 3332 6656
rect 3287 6616 3332 6644
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 3436 6644 3464 6684
rect 4338 6672 4344 6684
rect 4396 6672 4402 6724
rect 4706 6672 4712 6724
rect 4764 6712 4770 6724
rect 6457 6715 6515 6721
rect 6457 6712 6469 6715
rect 4764 6684 6469 6712
rect 4764 6672 4770 6684
rect 6457 6681 6469 6684
rect 6503 6681 6515 6715
rect 6457 6675 6515 6681
rect 7006 6672 7012 6724
rect 7064 6712 7070 6724
rect 8128 6712 8156 6743
rect 8202 6740 8208 6792
rect 8260 6780 8266 6792
rect 9784 6780 9812 6820
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 10962 6808 10968 6860
rect 11020 6848 11026 6860
rect 11149 6851 11207 6857
rect 11149 6848 11161 6851
rect 11020 6820 11161 6848
rect 11020 6808 11026 6820
rect 11149 6817 11161 6820
rect 11195 6817 11207 6851
rect 11149 6811 11207 6817
rect 8260 6752 9812 6780
rect 10137 6783 10195 6789
rect 8260 6740 8266 6752
rect 10137 6749 10149 6783
rect 10183 6780 10195 6783
rect 10594 6780 10600 6792
rect 10183 6752 10600 6780
rect 10183 6749 10195 6752
rect 10137 6743 10195 6749
rect 10594 6740 10600 6752
rect 10652 6740 10658 6792
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6780 10747 6783
rect 11256 6780 11284 6888
rect 12084 6857 12112 6888
rect 12158 6876 12164 6888
rect 12216 6876 12222 6928
rect 12710 6916 12716 6928
rect 12671 6888 12716 6916
rect 12710 6876 12716 6888
rect 12768 6876 12774 6928
rect 11333 6851 11391 6857
rect 11333 6817 11345 6851
rect 11379 6817 11391 6851
rect 11333 6811 11391 6817
rect 12069 6851 12127 6857
rect 12069 6817 12081 6851
rect 12115 6817 12127 6851
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 12069 6811 12127 6817
rect 12406 6820 12541 6848
rect 10735 6752 11284 6780
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 7064 6684 8156 6712
rect 7064 6672 7070 6684
rect 8478 6672 8484 6724
rect 8536 6712 8542 6724
rect 10229 6715 10287 6721
rect 10229 6712 10241 6715
rect 8536 6684 10241 6712
rect 8536 6672 8542 6684
rect 10229 6681 10241 6684
rect 10275 6712 10287 6715
rect 11348 6712 11376 6811
rect 10275 6684 11376 6712
rect 10275 6681 10287 6684
rect 10229 6675 10287 6681
rect 5537 6647 5595 6653
rect 5537 6644 5549 6647
rect 3436 6616 5549 6644
rect 5537 6613 5549 6616
rect 5583 6613 5595 6647
rect 5537 6607 5595 6613
rect 7193 6647 7251 6653
rect 7193 6613 7205 6647
rect 7239 6644 7251 6647
rect 7282 6644 7288 6656
rect 7239 6616 7288 6644
rect 7239 6613 7251 6616
rect 7193 6607 7251 6613
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 8570 6644 8576 6656
rect 8531 6616 8576 6644
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 8846 6604 8852 6656
rect 8904 6644 8910 6656
rect 9493 6647 9551 6653
rect 9493 6644 9505 6647
rect 8904 6616 9505 6644
rect 8904 6604 8910 6616
rect 9493 6613 9505 6616
rect 9539 6613 9551 6647
rect 9493 6607 9551 6613
rect 10134 6604 10140 6656
rect 10192 6644 10198 6656
rect 12406 6644 12434 6820
rect 12529 6817 12541 6820
rect 12575 6817 12587 6851
rect 12529 6811 12587 6817
rect 13170 6808 13176 6860
rect 13228 6848 13234 6860
rect 13449 6851 13507 6857
rect 13449 6848 13461 6851
rect 13228 6820 13461 6848
rect 13228 6808 13234 6820
rect 13449 6817 13461 6820
rect 13495 6817 13507 6851
rect 13449 6811 13507 6817
rect 13817 6851 13875 6857
rect 13817 6817 13829 6851
rect 13863 6848 13875 6851
rect 13906 6848 13912 6860
rect 13863 6820 13912 6848
rect 13863 6817 13875 6820
rect 13817 6811 13875 6817
rect 13906 6808 13912 6820
rect 13964 6808 13970 6860
rect 14826 6848 14832 6860
rect 14787 6820 14832 6848
rect 14826 6808 14832 6820
rect 14884 6808 14890 6860
rect 15194 6808 15200 6860
rect 15252 6848 15258 6860
rect 15657 6851 15715 6857
rect 15657 6848 15669 6851
rect 15252 6820 15669 6848
rect 15252 6808 15258 6820
rect 15657 6817 15669 6820
rect 15703 6817 15715 6851
rect 15657 6811 15715 6817
rect 16206 6808 16212 6860
rect 16264 6848 16270 6860
rect 16301 6851 16359 6857
rect 16301 6848 16313 6851
rect 16264 6820 16313 6848
rect 16264 6808 16270 6820
rect 16301 6817 16313 6820
rect 16347 6817 16359 6851
rect 16301 6811 16359 6817
rect 15013 6715 15071 6721
rect 15013 6681 15025 6715
rect 15059 6712 15071 6715
rect 15378 6712 15384 6724
rect 15059 6684 15384 6712
rect 15059 6681 15071 6684
rect 15013 6675 15071 6681
rect 15378 6672 15384 6684
rect 15436 6672 15442 6724
rect 10192 6616 12434 6644
rect 10192 6604 10198 6616
rect 15286 6604 15292 6656
rect 15344 6644 15350 6656
rect 15473 6647 15531 6653
rect 15473 6644 15485 6647
rect 15344 6616 15485 6644
rect 15344 6604 15350 6616
rect 15473 6613 15485 6616
rect 15519 6613 15531 6647
rect 15473 6607 15531 6613
rect 1104 6554 17296 6576
rect 1104 6502 3680 6554
rect 3732 6502 3744 6554
rect 3796 6502 3808 6554
rect 3860 6502 3872 6554
rect 3924 6502 9078 6554
rect 9130 6502 9142 6554
rect 9194 6502 9206 6554
rect 9258 6502 9270 6554
rect 9322 6502 14475 6554
rect 14527 6502 14539 6554
rect 14591 6502 14603 6554
rect 14655 6502 14667 6554
rect 14719 6502 17296 6554
rect 1104 6480 17296 6502
rect 4062 6400 4068 6452
rect 4120 6440 4126 6452
rect 4433 6443 4491 6449
rect 4433 6440 4445 6443
rect 4120 6412 4445 6440
rect 4120 6400 4126 6412
rect 4433 6409 4445 6412
rect 4479 6409 4491 6443
rect 5442 6440 5448 6452
rect 5403 6412 5448 6440
rect 4433 6403 4491 6409
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 8202 6440 8208 6452
rect 5552 6412 8208 6440
rect 4890 6332 4896 6384
rect 4948 6372 4954 6384
rect 5552 6372 5580 6412
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 8386 6440 8392 6452
rect 8347 6412 8392 6440
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 8662 6400 8668 6452
rect 8720 6440 8726 6452
rect 9033 6443 9091 6449
rect 9033 6440 9045 6443
rect 8720 6412 9045 6440
rect 8720 6400 8726 6412
rect 9033 6409 9045 6412
rect 9079 6409 9091 6443
rect 9033 6403 9091 6409
rect 10410 6400 10416 6452
rect 10468 6440 10474 6452
rect 10962 6440 10968 6452
rect 10468 6412 10968 6440
rect 10468 6400 10474 6412
rect 10962 6400 10968 6412
rect 11020 6440 11026 6452
rect 13449 6443 13507 6449
rect 13449 6440 13461 6443
rect 11020 6412 13461 6440
rect 11020 6400 11026 6412
rect 13449 6409 13461 6412
rect 13495 6409 13507 6443
rect 14182 6440 14188 6452
rect 14143 6412 14188 6440
rect 13449 6403 13507 6409
rect 14182 6400 14188 6412
rect 14240 6400 14246 6452
rect 15381 6443 15439 6449
rect 15381 6409 15393 6443
rect 15427 6440 15439 6443
rect 16206 6440 16212 6452
rect 15427 6412 16212 6440
rect 15427 6409 15439 6412
rect 15381 6403 15439 6409
rect 16206 6400 16212 6412
rect 16264 6400 16270 6452
rect 7374 6372 7380 6384
rect 4948 6344 5580 6372
rect 5920 6344 7380 6372
rect 4948 6332 4954 6344
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6304 1823 6307
rect 2498 6304 2504 6316
rect 1811 6276 2504 6304
rect 1811 6273 1823 6276
rect 1765 6267 1823 6273
rect 2498 6264 2504 6276
rect 2556 6264 2562 6316
rect 4338 6304 4344 6316
rect 3252 6276 4344 6304
rect 1946 6236 1952 6248
rect 1907 6208 1952 6236
rect 1946 6196 1952 6208
rect 2004 6196 2010 6248
rect 2682 6196 2688 6248
rect 2740 6236 2746 6248
rect 3252 6245 3280 6276
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 5920 6313 5948 6344
rect 7374 6332 7380 6344
rect 7432 6332 7438 6384
rect 10134 6372 10140 6384
rect 8312 6344 10140 6372
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6273 5963 6307
rect 7282 6304 7288 6316
rect 7243 6276 7288 6304
rect 5905 6267 5963 6273
rect 7282 6264 7288 6276
rect 7340 6264 7346 6316
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6304 7527 6307
rect 8018 6304 8024 6316
rect 7515 6276 8024 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 3237 6239 3295 6245
rect 3237 6236 3249 6239
rect 2740 6208 3249 6236
rect 2740 6196 2746 6208
rect 3237 6205 3249 6208
rect 3283 6205 3295 6239
rect 3237 6199 3295 6205
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 4522 6236 4528 6248
rect 3927 6208 4528 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 4522 6196 4528 6208
rect 4580 6196 4586 6248
rect 4617 6239 4675 6245
rect 4617 6205 4629 6239
rect 4663 6236 4675 6239
rect 4706 6236 4712 6248
rect 4663 6208 4712 6236
rect 4663 6205 4675 6208
rect 4617 6199 4675 6205
rect 1857 6171 1915 6177
rect 1857 6137 1869 6171
rect 1903 6168 1915 6171
rect 2961 6171 3019 6177
rect 1903 6140 2774 6168
rect 1903 6137 1915 6140
rect 1857 6131 1915 6137
rect 1946 6060 1952 6112
rect 2004 6100 2010 6112
rect 2317 6103 2375 6109
rect 2317 6100 2329 6103
rect 2004 6072 2329 6100
rect 2004 6060 2010 6072
rect 2317 6069 2329 6072
rect 2363 6069 2375 6103
rect 2746 6100 2774 6140
rect 2961 6137 2973 6171
rect 3007 6168 3019 6171
rect 4632 6168 4660 6199
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 5626 6236 5632 6248
rect 5587 6208 5632 6236
rect 5626 6196 5632 6208
rect 5684 6196 5690 6248
rect 5813 6239 5871 6245
rect 5813 6205 5825 6239
rect 5859 6236 5871 6239
rect 5994 6236 6000 6248
rect 5859 6208 6000 6236
rect 5859 6205 5871 6208
rect 5813 6199 5871 6205
rect 5994 6196 6000 6208
rect 6052 6236 6058 6248
rect 7742 6236 7748 6248
rect 6052 6208 7748 6236
rect 6052 6196 6058 6208
rect 7742 6196 7748 6208
rect 7800 6236 7806 6248
rect 8312 6245 8340 6344
rect 10134 6332 10140 6344
rect 10192 6332 10198 6384
rect 11054 6332 11060 6384
rect 11112 6372 11118 6384
rect 12069 6375 12127 6381
rect 12069 6372 12081 6375
rect 11112 6344 12081 6372
rect 11112 6332 11118 6344
rect 12069 6341 12081 6344
rect 12115 6341 12127 6375
rect 12069 6335 12127 6341
rect 12250 6332 12256 6384
rect 12308 6372 12314 6384
rect 12308 6344 14872 6372
rect 12308 6332 12314 6344
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 8628 6276 12449 6304
rect 8628 6264 8634 6276
rect 8297 6239 8355 6245
rect 8297 6236 8309 6239
rect 7800 6208 8309 6236
rect 7800 6196 7806 6208
rect 8297 6205 8309 6208
rect 8343 6205 8355 6239
rect 8297 6199 8355 6205
rect 8478 6196 8484 6248
rect 8536 6236 8542 6248
rect 8941 6239 8999 6245
rect 8536 6208 8581 6236
rect 8536 6196 8542 6208
rect 8941 6205 8953 6239
rect 8987 6205 8999 6239
rect 8941 6199 8999 6205
rect 3007 6140 4660 6168
rect 3007 6137 3019 6140
rect 2961 6131 3019 6137
rect 7374 6128 7380 6180
rect 7432 6168 7438 6180
rect 8956 6168 8984 6199
rect 9030 6196 9036 6248
rect 9088 6236 9094 6248
rect 9876 6245 9904 6276
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 14844 6304 14872 6344
rect 15841 6307 15899 6313
rect 15841 6304 15853 6307
rect 14844 6276 15853 6304
rect 9217 6239 9275 6245
rect 9217 6236 9229 6239
rect 9088 6208 9229 6236
rect 9088 6196 9094 6208
rect 9217 6205 9229 6208
rect 9263 6205 9275 6239
rect 9217 6199 9275 6205
rect 9861 6239 9919 6245
rect 9861 6205 9873 6239
rect 9907 6205 9919 6239
rect 10410 6236 10416 6248
rect 10371 6208 10416 6236
rect 9861 6199 9919 6205
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 10594 6196 10600 6248
rect 10652 6236 10658 6248
rect 10965 6239 11023 6245
rect 10965 6236 10977 6239
rect 10652 6208 10977 6236
rect 10652 6196 10658 6208
rect 10965 6205 10977 6208
rect 11011 6205 11023 6239
rect 10965 6199 11023 6205
rect 13541 6239 13599 6245
rect 13541 6205 13553 6239
rect 13587 6236 13599 6239
rect 13722 6236 13728 6248
rect 13587 6208 13728 6236
rect 13587 6205 13599 6208
rect 13541 6199 13599 6205
rect 13722 6196 13728 6208
rect 13780 6196 13786 6248
rect 14366 6236 14372 6248
rect 14327 6208 14372 6236
rect 14366 6196 14372 6208
rect 14424 6196 14430 6248
rect 14844 6245 14872 6276
rect 15841 6273 15853 6276
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6205 14887 6239
rect 15378 6236 15384 6248
rect 15339 6208 15384 6236
rect 14829 6199 14887 6205
rect 15378 6196 15384 6208
rect 15436 6196 15442 6248
rect 16206 6236 16212 6248
rect 16167 6208 16212 6236
rect 16206 6196 16212 6208
rect 16264 6196 16270 6248
rect 10226 6168 10232 6180
rect 7432 6140 8984 6168
rect 9048 6140 10232 6168
rect 7432 6128 7438 6140
rect 4246 6100 4252 6112
rect 2746 6072 4252 6100
rect 2317 6063 2375 6069
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 6822 6100 6828 6112
rect 6783 6072 6828 6100
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 7193 6103 7251 6109
rect 7193 6069 7205 6103
rect 7239 6100 7251 6103
rect 7282 6100 7288 6112
rect 7239 6072 7288 6100
rect 7239 6069 7251 6072
rect 7193 6063 7251 6069
rect 7282 6060 7288 6072
rect 7340 6060 7346 6112
rect 8110 6100 8116 6112
rect 8071 6072 8116 6100
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 8478 6060 8484 6112
rect 8536 6100 8542 6112
rect 9048 6100 9076 6140
rect 10226 6128 10232 6140
rect 10284 6128 10290 6180
rect 10321 6171 10379 6177
rect 10321 6137 10333 6171
rect 10367 6168 10379 6171
rect 10367 6140 11192 6168
rect 10367 6137 10379 6140
rect 10321 6131 10379 6137
rect 8536 6072 9076 6100
rect 9401 6103 9459 6109
rect 8536 6060 8542 6072
rect 9401 6069 9413 6103
rect 9447 6100 9459 6103
rect 9858 6100 9864 6112
rect 9447 6072 9864 6100
rect 9447 6069 9459 6072
rect 9401 6063 9459 6069
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 11164 6109 11192 6140
rect 11149 6103 11207 6109
rect 11149 6069 11161 6103
rect 11195 6100 11207 6103
rect 12069 6103 12127 6109
rect 12069 6100 12081 6103
rect 11195 6072 12081 6100
rect 11195 6069 11207 6072
rect 11149 6063 11207 6069
rect 12069 6069 12081 6072
rect 12115 6069 12127 6103
rect 12069 6063 12127 6069
rect 1104 6010 17296 6032
rect 1104 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 6571 6010
rect 6623 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 11904 6010
rect 11956 5958 11968 6010
rect 12020 5958 17296 6010
rect 1104 5936 17296 5958
rect 2225 5899 2283 5905
rect 2225 5865 2237 5899
rect 2271 5896 2283 5899
rect 2314 5896 2320 5908
rect 2271 5868 2320 5896
rect 2271 5865 2283 5868
rect 2225 5859 2283 5865
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 4525 5899 4583 5905
rect 4525 5865 4537 5899
rect 4571 5896 4583 5899
rect 4798 5896 4804 5908
rect 4571 5868 4804 5896
rect 4571 5865 4583 5868
rect 4525 5859 4583 5865
rect 4798 5856 4804 5868
rect 4856 5856 4862 5908
rect 6273 5899 6331 5905
rect 6273 5865 6285 5899
rect 6319 5896 6331 5899
rect 6914 5896 6920 5908
rect 6319 5868 6920 5896
rect 6319 5865 6331 5868
rect 6273 5859 6331 5865
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 7300 5868 7512 5896
rect 4890 5828 4896 5840
rect 4816 5800 4896 5828
rect 1578 5720 1584 5772
rect 1636 5760 1642 5772
rect 1857 5763 1915 5769
rect 1857 5760 1869 5763
rect 1636 5732 1869 5760
rect 1636 5720 1642 5732
rect 1857 5729 1869 5732
rect 1903 5729 1915 5763
rect 1857 5723 1915 5729
rect 2685 5763 2743 5769
rect 2685 5729 2697 5763
rect 2731 5760 2743 5763
rect 2866 5760 2872 5772
rect 2731 5732 2872 5760
rect 2731 5729 2743 5732
rect 2685 5723 2743 5729
rect 2866 5720 2872 5732
rect 2924 5720 2930 5772
rect 4614 5760 4620 5772
rect 4575 5732 4620 5760
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 4816 5769 4844 5800
rect 4890 5788 4896 5800
rect 4948 5788 4954 5840
rect 6365 5831 6423 5837
rect 6365 5797 6377 5831
rect 6411 5828 6423 5831
rect 7300 5828 7328 5868
rect 6411 5800 7328 5828
rect 7484 5828 7512 5868
rect 7650 5856 7656 5908
rect 7708 5896 7714 5908
rect 11606 5896 11612 5908
rect 7708 5868 11612 5896
rect 7708 5856 7714 5868
rect 11606 5856 11612 5868
rect 11664 5856 11670 5908
rect 12526 5856 12532 5908
rect 12584 5896 12590 5908
rect 13633 5899 13691 5905
rect 13633 5896 13645 5899
rect 12584 5868 13645 5896
rect 12584 5856 12590 5868
rect 13633 5865 13645 5868
rect 13679 5865 13691 5899
rect 13633 5859 13691 5865
rect 7484 5800 11100 5828
rect 6411 5797 6423 5800
rect 6365 5791 6423 5797
rect 4801 5763 4859 5769
rect 4801 5729 4813 5763
rect 4847 5729 4859 5763
rect 4801 5723 4859 5729
rect 5626 5720 5632 5772
rect 5684 5760 5690 5772
rect 7469 5763 7527 5769
rect 7469 5760 7481 5763
rect 5684 5732 7481 5760
rect 5684 5720 5690 5732
rect 7469 5729 7481 5732
rect 7515 5760 7527 5763
rect 8202 5760 8208 5772
rect 7515 5732 7880 5760
rect 8163 5732 8208 5760
rect 7515 5729 7527 5732
rect 7469 5723 7527 5729
rect 5258 5692 5264 5704
rect 5219 5664 5264 5692
rect 5258 5652 5264 5664
rect 5316 5652 5322 5704
rect 5718 5652 5724 5704
rect 5776 5692 5782 5704
rect 6454 5692 6460 5704
rect 5776 5664 6460 5692
rect 5776 5652 5782 5664
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 7742 5692 7748 5704
rect 7703 5664 7748 5692
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 7852 5692 7880 5732
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5760 9551 5763
rect 10962 5760 10968 5772
rect 9539 5732 10968 5760
rect 9539 5729 9551 5732
rect 9493 5723 9551 5729
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 8478 5692 8484 5704
rect 7852 5664 8484 5692
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5661 10195 5695
rect 10502 5692 10508 5704
rect 10463 5664 10508 5692
rect 10137 5655 10195 5661
rect 2225 5627 2283 5633
rect 2225 5593 2237 5627
rect 2271 5624 2283 5627
rect 2774 5624 2780 5636
rect 2271 5596 2780 5624
rect 2271 5593 2283 5596
rect 2225 5587 2283 5593
rect 2774 5584 2780 5596
rect 2832 5584 2838 5636
rect 2869 5627 2927 5633
rect 2869 5593 2881 5627
rect 2915 5624 2927 5627
rect 7006 5624 7012 5636
rect 2915 5596 7012 5624
rect 2915 5593 2927 5596
rect 2869 5587 2927 5593
rect 7006 5584 7012 5596
rect 7064 5584 7070 5636
rect 7558 5584 7564 5636
rect 7616 5624 7622 5636
rect 8297 5627 8355 5633
rect 8297 5624 8309 5627
rect 7616 5596 8309 5624
rect 7616 5584 7622 5596
rect 8297 5593 8309 5596
rect 8343 5593 8355 5627
rect 10152 5624 10180 5655
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 10965 5627 11023 5633
rect 10965 5624 10977 5627
rect 10152 5596 10977 5624
rect 8297 5587 8355 5593
rect 10965 5593 10977 5596
rect 11011 5593 11023 5627
rect 11072 5624 11100 5800
rect 12250 5788 12256 5840
rect 12308 5828 12314 5840
rect 12989 5831 13047 5837
rect 12989 5828 13001 5831
rect 12308 5800 13001 5828
rect 12308 5788 12314 5800
rect 12989 5797 13001 5800
rect 13035 5797 13047 5831
rect 12989 5791 13047 5797
rect 13354 5788 13360 5840
rect 13412 5828 13418 5840
rect 15562 5828 15568 5840
rect 13412 5800 14780 5828
rect 13412 5788 13418 5800
rect 11146 5720 11152 5772
rect 11204 5760 11210 5772
rect 11606 5760 11612 5772
rect 11204 5732 11249 5760
rect 11567 5732 11612 5760
rect 11204 5720 11210 5732
rect 11606 5720 11612 5732
rect 11664 5720 11670 5772
rect 12066 5720 12072 5772
rect 12124 5760 12130 5772
rect 12161 5763 12219 5769
rect 12161 5760 12173 5763
rect 12124 5732 12173 5760
rect 12124 5720 12130 5732
rect 12161 5729 12173 5732
rect 12207 5729 12219 5763
rect 13814 5760 13820 5772
rect 13775 5732 13820 5760
rect 12161 5723 12219 5729
rect 13814 5720 13820 5732
rect 13872 5720 13878 5772
rect 14752 5769 14780 5800
rect 14844 5800 15568 5828
rect 14737 5763 14795 5769
rect 14737 5729 14749 5763
rect 14783 5729 14795 5763
rect 14737 5723 14795 5729
rect 13081 5695 13139 5701
rect 13081 5661 13093 5695
rect 13127 5692 13139 5695
rect 14369 5695 14427 5701
rect 14369 5692 14381 5695
rect 13127 5664 14381 5692
rect 13127 5661 13139 5664
rect 13081 5655 13139 5661
rect 14369 5661 14381 5664
rect 14415 5661 14427 5695
rect 14369 5655 14427 5661
rect 14844 5624 14872 5800
rect 15562 5788 15568 5800
rect 15620 5788 15626 5840
rect 15197 5763 15255 5769
rect 15197 5729 15209 5763
rect 15243 5760 15255 5763
rect 15378 5760 15384 5772
rect 15243 5732 15384 5760
rect 15243 5729 15255 5732
rect 15197 5723 15255 5729
rect 15378 5720 15384 5732
rect 15436 5720 15442 5772
rect 15841 5695 15899 5701
rect 15841 5692 15853 5695
rect 15396 5664 15853 5692
rect 15396 5633 15424 5664
rect 15841 5661 15853 5664
rect 15887 5661 15899 5695
rect 15841 5655 15899 5661
rect 15930 5652 15936 5704
rect 15988 5692 15994 5704
rect 16209 5695 16267 5701
rect 16209 5692 16221 5695
rect 15988 5664 16221 5692
rect 15988 5652 15994 5664
rect 16209 5661 16221 5664
rect 16255 5661 16267 5695
rect 16209 5655 16267 5661
rect 11072 5596 14872 5624
rect 15381 5627 15439 5633
rect 10965 5587 11023 5593
rect 15381 5593 15393 5627
rect 15427 5593 15439 5627
rect 15381 5587 15439 5593
rect 5902 5556 5908 5568
rect 5863 5528 5908 5556
rect 5902 5516 5908 5528
rect 5960 5516 5966 5568
rect 7282 5556 7288 5568
rect 7243 5528 7288 5556
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 7653 5559 7711 5565
rect 7653 5525 7665 5559
rect 7699 5556 7711 5559
rect 8386 5556 8392 5568
rect 7699 5528 8392 5556
rect 7699 5525 7711 5528
rect 7653 5519 7711 5525
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 9677 5559 9735 5565
rect 9677 5525 9689 5559
rect 9723 5556 9735 5559
rect 9950 5556 9956 5568
rect 9723 5528 9956 5556
rect 9723 5525 9735 5528
rect 9677 5519 9735 5525
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 10134 5556 10140 5568
rect 10095 5528 10140 5556
rect 10134 5516 10140 5528
rect 10192 5516 10198 5568
rect 12158 5556 12164 5568
rect 12119 5528 12164 5556
rect 12158 5516 12164 5528
rect 12216 5516 12222 5568
rect 14366 5556 14372 5568
rect 14327 5528 14372 5556
rect 14366 5516 14372 5528
rect 14424 5556 14430 5568
rect 14826 5556 14832 5568
rect 14424 5528 14832 5556
rect 14424 5516 14430 5528
rect 14826 5516 14832 5528
rect 14884 5516 14890 5568
rect 15470 5516 15476 5568
rect 15528 5556 15534 5568
rect 15841 5559 15899 5565
rect 15841 5556 15853 5559
rect 15528 5528 15853 5556
rect 15528 5516 15534 5528
rect 15841 5525 15853 5528
rect 15887 5525 15899 5559
rect 15841 5519 15899 5525
rect 1104 5466 17296 5488
rect 1104 5414 3680 5466
rect 3732 5414 3744 5466
rect 3796 5414 3808 5466
rect 3860 5414 3872 5466
rect 3924 5414 9078 5466
rect 9130 5414 9142 5466
rect 9194 5414 9206 5466
rect 9258 5414 9270 5466
rect 9322 5414 14475 5466
rect 14527 5414 14539 5466
rect 14591 5414 14603 5466
rect 14655 5414 14667 5466
rect 14719 5414 17296 5466
rect 1104 5392 17296 5414
rect 2314 5352 2320 5364
rect 2275 5324 2320 5352
rect 2314 5312 2320 5324
rect 2372 5312 2378 5364
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 2832 5324 2877 5352
rect 2832 5312 2838 5324
rect 7190 5312 7196 5364
rect 7248 5352 7254 5364
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 7248 5324 7389 5352
rect 7248 5312 7254 5324
rect 7377 5321 7389 5324
rect 7423 5352 7435 5355
rect 8202 5352 8208 5364
rect 7423 5324 8208 5352
rect 7423 5321 7435 5324
rect 7377 5315 7435 5321
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 10134 5312 10140 5364
rect 10192 5352 10198 5364
rect 10229 5355 10287 5361
rect 10229 5352 10241 5355
rect 10192 5324 10241 5352
rect 10192 5312 10198 5324
rect 10229 5321 10241 5324
rect 10275 5321 10287 5355
rect 10229 5315 10287 5321
rect 12713 5355 12771 5361
rect 12713 5321 12725 5355
rect 12759 5352 12771 5355
rect 14366 5352 14372 5364
rect 12759 5324 14372 5352
rect 12759 5321 12771 5324
rect 12713 5315 12771 5321
rect 14366 5312 14372 5324
rect 14424 5312 14430 5364
rect 9769 5287 9827 5293
rect 9769 5253 9781 5287
rect 9815 5284 9827 5287
rect 11606 5284 11612 5296
rect 9815 5256 11612 5284
rect 9815 5253 9827 5256
rect 9769 5247 9827 5253
rect 11606 5244 11612 5256
rect 11664 5244 11670 5296
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5216 4491 5219
rect 4798 5216 4804 5228
rect 4479 5188 4804 5216
rect 4479 5185 4491 5188
rect 4433 5179 4491 5185
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 6454 5176 6460 5228
rect 6512 5216 6518 5228
rect 8018 5216 8024 5228
rect 6512 5188 8024 5216
rect 6512 5176 6518 5188
rect 8018 5176 8024 5188
rect 8076 5216 8082 5228
rect 8938 5216 8944 5228
rect 8076 5188 8944 5216
rect 8076 5176 8082 5188
rect 8938 5176 8944 5188
rect 8996 5216 9002 5228
rect 9125 5219 9183 5225
rect 9125 5216 9137 5219
rect 8996 5188 9137 5216
rect 8996 5176 9002 5188
rect 9125 5185 9137 5188
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 13078 5176 13084 5228
rect 13136 5216 13142 5228
rect 14369 5219 14427 5225
rect 14369 5216 14381 5219
rect 13136 5188 14381 5216
rect 13136 5176 13142 5188
rect 14369 5185 14381 5188
rect 14415 5185 14427 5219
rect 15470 5216 15476 5228
rect 15431 5188 15476 5216
rect 14369 5179 14427 5185
rect 15470 5176 15476 5188
rect 15528 5176 15534 5228
rect 1578 5108 1584 5160
rect 1636 5148 1642 5160
rect 1765 5151 1823 5157
rect 1765 5148 1777 5151
rect 1636 5120 1777 5148
rect 1636 5108 1642 5120
rect 1765 5117 1777 5120
rect 1811 5117 1823 5151
rect 1765 5111 1823 5117
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5148 2375 5151
rect 2406 5148 2412 5160
rect 2363 5120 2412 5148
rect 2363 5117 2375 5120
rect 2317 5111 2375 5117
rect 2406 5108 2412 5120
rect 2464 5148 2470 5160
rect 2961 5151 3019 5157
rect 2961 5148 2973 5151
rect 2464 5120 2973 5148
rect 2464 5108 2470 5120
rect 2961 5117 2973 5120
rect 3007 5117 3019 5151
rect 2961 5111 3019 5117
rect 3973 5151 4031 5157
rect 3973 5117 3985 5151
rect 4019 5117 4031 5151
rect 5258 5148 5264 5160
rect 5219 5120 5264 5148
rect 3973 5111 4031 5117
rect 3988 5080 4016 5111
rect 5258 5108 5264 5120
rect 5316 5108 5322 5160
rect 6822 5148 6828 5160
rect 6783 5120 6828 5148
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 7374 5148 7380 5160
rect 7335 5120 7380 5148
rect 7374 5108 7380 5120
rect 7432 5108 7438 5160
rect 8110 5108 8116 5160
rect 8168 5148 8174 5160
rect 8205 5151 8263 5157
rect 8205 5148 8217 5151
rect 8168 5120 8217 5148
rect 8168 5108 8174 5120
rect 8205 5117 8217 5120
rect 8251 5117 8263 5151
rect 8205 5111 8263 5117
rect 9401 5151 9459 5157
rect 9401 5117 9413 5151
rect 9447 5148 9459 5151
rect 9766 5148 9772 5160
rect 9447 5120 9772 5148
rect 9447 5117 9459 5120
rect 9401 5111 9459 5117
rect 9766 5108 9772 5120
rect 9824 5108 9830 5160
rect 10229 5151 10287 5157
rect 10229 5117 10241 5151
rect 10275 5117 10287 5151
rect 10229 5111 10287 5117
rect 5074 5080 5080 5092
rect 3988 5052 5080 5080
rect 5074 5040 5080 5052
rect 5132 5040 5138 5092
rect 8018 5040 8024 5092
rect 8076 5080 8082 5092
rect 10244 5080 10272 5111
rect 10502 5108 10508 5160
rect 10560 5148 10566 5160
rect 10781 5151 10839 5157
rect 10781 5148 10793 5151
rect 10560 5120 10793 5148
rect 10560 5108 10566 5120
rect 10781 5117 10793 5120
rect 10827 5117 10839 5151
rect 10781 5111 10839 5117
rect 11238 5108 11244 5160
rect 11296 5148 11302 5160
rect 12066 5148 12072 5160
rect 11296 5120 12072 5148
rect 11296 5108 11302 5120
rect 12066 5108 12072 5120
rect 12124 5148 12130 5160
rect 12253 5151 12311 5157
rect 12253 5148 12265 5151
rect 12124 5120 12265 5148
rect 12124 5108 12130 5120
rect 12253 5117 12265 5120
rect 12299 5148 12311 5151
rect 12713 5151 12771 5157
rect 12713 5148 12725 5151
rect 12299 5120 12725 5148
rect 12299 5117 12311 5120
rect 12253 5111 12311 5117
rect 12713 5117 12725 5120
rect 12759 5117 12771 5151
rect 12713 5111 12771 5117
rect 13265 5151 13323 5157
rect 13265 5117 13277 5151
rect 13311 5148 13323 5151
rect 13354 5148 13360 5160
rect 13311 5120 13360 5148
rect 13311 5117 13323 5120
rect 13265 5111 13323 5117
rect 13354 5108 13360 5120
rect 13412 5108 13418 5160
rect 14274 5108 14280 5160
rect 14332 5148 14338 5160
rect 14461 5151 14519 5157
rect 14461 5148 14473 5151
rect 14332 5120 14473 5148
rect 14332 5108 14338 5120
rect 14461 5117 14473 5120
rect 14507 5117 14519 5151
rect 14461 5111 14519 5117
rect 14737 5151 14795 5157
rect 14737 5117 14749 5151
rect 14783 5117 14795 5151
rect 14737 5111 14795 5117
rect 15289 5151 15347 5157
rect 15289 5117 15301 5151
rect 15335 5148 15347 5151
rect 15378 5148 15384 5160
rect 15335 5120 15384 5148
rect 15335 5117 15347 5120
rect 15289 5111 15347 5117
rect 11146 5080 11152 5092
rect 8076 5052 11152 5080
rect 8076 5040 8082 5052
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 14182 5080 14188 5092
rect 14143 5052 14188 5080
rect 14182 5040 14188 5052
rect 14240 5040 14246 5092
rect 3789 5015 3847 5021
rect 3789 4981 3801 5015
rect 3835 5012 3847 5015
rect 4154 5012 4160 5024
rect 3835 4984 4160 5012
rect 3835 4981 3847 4984
rect 3789 4975 3847 4981
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 7742 4972 7748 5024
rect 7800 5012 7806 5024
rect 8113 5015 8171 5021
rect 8113 5012 8125 5015
rect 7800 4984 8125 5012
rect 7800 4972 7806 4984
rect 8113 4981 8125 4984
rect 8159 4981 8171 5015
rect 8570 5012 8576 5024
rect 8531 4984 8576 5012
rect 8113 4975 8171 4981
rect 8570 4972 8576 4984
rect 8628 4972 8634 5024
rect 8662 4972 8668 5024
rect 8720 5012 8726 5024
rect 9309 5015 9367 5021
rect 9309 5012 9321 5015
rect 8720 4984 9321 5012
rect 8720 4972 8726 4984
rect 9309 4981 9321 4984
rect 9355 4981 9367 5015
rect 12066 5012 12072 5024
rect 12027 4984 12072 5012
rect 9309 4975 9367 4981
rect 12066 4972 12072 4984
rect 12124 4972 12130 5024
rect 13998 4972 14004 5024
rect 14056 5012 14062 5024
rect 14752 5012 14780 5111
rect 15378 5108 15384 5120
rect 15436 5108 15442 5160
rect 15841 5151 15899 5157
rect 15841 5117 15853 5151
rect 15887 5148 15899 5151
rect 15930 5148 15936 5160
rect 15887 5120 15936 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 15930 5108 15936 5120
rect 15988 5108 15994 5160
rect 14056 4984 14780 5012
rect 14056 4972 14062 4984
rect 1104 4922 17296 4944
rect 1104 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 6571 4922
rect 6623 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 11904 4922
rect 11956 4870 11968 4922
rect 12020 4870 17296 4922
rect 1104 4848 17296 4870
rect 3510 4768 3516 4820
rect 3568 4808 3574 4820
rect 9398 4808 9404 4820
rect 3568 4780 7696 4808
rect 9359 4780 9404 4808
rect 3568 4768 3574 4780
rect 4617 4743 4675 4749
rect 1964 4712 3188 4740
rect 1964 4684 1992 4712
rect 1765 4675 1823 4681
rect 1765 4641 1777 4675
rect 1811 4672 1823 4675
rect 1946 4672 1952 4684
rect 1811 4644 1952 4672
rect 1811 4641 1823 4644
rect 1765 4635 1823 4641
rect 1946 4632 1952 4644
rect 2004 4632 2010 4684
rect 2317 4675 2375 4681
rect 2317 4641 2329 4675
rect 2363 4672 2375 4675
rect 2406 4672 2412 4684
rect 2363 4644 2412 4672
rect 2363 4641 2375 4644
rect 2317 4635 2375 4641
rect 2406 4632 2412 4644
rect 2464 4632 2470 4684
rect 3160 4681 3188 4712
rect 4617 4709 4629 4743
rect 4663 4740 4675 4743
rect 7374 4740 7380 4752
rect 4663 4712 7380 4740
rect 4663 4709 4675 4712
rect 4617 4703 4675 4709
rect 7374 4700 7380 4712
rect 7432 4740 7438 4752
rect 7668 4740 7696 4780
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 10134 4768 10140 4820
rect 10192 4808 10198 4820
rect 10229 4811 10287 4817
rect 10229 4808 10241 4811
rect 10192 4780 10241 4808
rect 10192 4768 10198 4780
rect 10229 4777 10241 4780
rect 10275 4777 10287 4811
rect 10229 4771 10287 4777
rect 10778 4768 10784 4820
rect 10836 4808 10842 4820
rect 12069 4811 12127 4817
rect 10836 4780 12020 4808
rect 10836 4768 10842 4780
rect 11238 4740 11244 4752
rect 7432 4712 7604 4740
rect 7668 4712 9628 4740
rect 11199 4712 11244 4740
rect 7432 4700 7438 4712
rect 3145 4675 3203 4681
rect 3145 4641 3157 4675
rect 3191 4641 3203 4675
rect 3145 4635 3203 4641
rect 4893 4675 4951 4681
rect 4893 4641 4905 4675
rect 4939 4641 4951 4675
rect 5534 4672 5540 4684
rect 5495 4644 5540 4672
rect 4893 4635 4951 4641
rect 2774 4564 2780 4616
rect 2832 4604 2838 4616
rect 4908 4604 4936 4635
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 5902 4632 5908 4684
rect 5960 4672 5966 4684
rect 5997 4675 6055 4681
rect 5997 4672 6009 4675
rect 5960 4644 6009 4672
rect 5960 4632 5966 4644
rect 5997 4641 6009 4644
rect 6043 4641 6055 4675
rect 5997 4635 6055 4641
rect 6825 4675 6883 4681
rect 6825 4641 6837 4675
rect 6871 4672 6883 4675
rect 7466 4672 7472 4684
rect 6871 4644 7472 4672
rect 6871 4641 6883 4644
rect 6825 4635 6883 4641
rect 7466 4632 7472 4644
rect 7524 4632 7530 4684
rect 7576 4681 7604 4712
rect 7561 4675 7619 4681
rect 7561 4641 7573 4675
rect 7607 4641 7619 4675
rect 8018 4672 8024 4684
rect 7979 4644 8024 4672
rect 7561 4635 7619 4641
rect 8018 4632 8024 4644
rect 8076 4632 8082 4684
rect 8570 4672 8576 4684
rect 8531 4644 8576 4672
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 9600 4681 9628 4712
rect 11238 4700 11244 4712
rect 11296 4700 11302 4752
rect 11992 4740 12020 4780
rect 12069 4777 12081 4811
rect 12115 4808 12127 4811
rect 12158 4808 12164 4820
rect 12115 4780 12164 4808
rect 12115 4777 12127 4780
rect 12069 4771 12127 4777
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 15013 4811 15071 4817
rect 15013 4777 15025 4811
rect 15059 4808 15071 4811
rect 15286 4808 15292 4820
rect 15059 4780 15292 4808
rect 15059 4777 15071 4780
rect 15013 4771 15071 4777
rect 15286 4768 15292 4780
rect 15344 4768 15350 4820
rect 15473 4811 15531 4817
rect 15473 4777 15485 4811
rect 15519 4808 15531 4811
rect 15930 4808 15936 4820
rect 15519 4780 15936 4808
rect 15519 4777 15531 4780
rect 15473 4771 15531 4777
rect 15930 4768 15936 4780
rect 15988 4768 15994 4820
rect 16206 4768 16212 4820
rect 16264 4808 16270 4820
rect 16301 4811 16359 4817
rect 16301 4808 16313 4811
rect 16264 4780 16313 4808
rect 16264 4768 16270 4780
rect 16301 4777 16313 4780
rect 16347 4777 16359 4811
rect 16301 4771 16359 4777
rect 15105 4743 15163 4749
rect 15105 4740 15117 4743
rect 11992 4712 15117 4740
rect 15105 4709 15117 4712
rect 15151 4709 15163 4743
rect 15746 4740 15752 4752
rect 15105 4703 15163 4709
rect 15212 4712 15752 4740
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4641 9643 4675
rect 9585 4635 9643 4641
rect 11057 4675 11115 4681
rect 11057 4641 11069 4675
rect 11103 4641 11115 4675
rect 11057 4635 11115 4641
rect 5074 4604 5080 4616
rect 2832 4576 2877 4604
rect 4908 4576 5080 4604
rect 2832 4564 2838 4576
rect 5074 4564 5080 4576
rect 5132 4604 5138 4616
rect 6733 4607 6791 4613
rect 6733 4604 6745 4607
rect 5132 4576 6745 4604
rect 5132 4564 5138 4576
rect 6733 4573 6745 4576
rect 6779 4604 6791 4607
rect 11072 4604 11100 4635
rect 11606 4632 11612 4684
rect 11664 4672 11670 4684
rect 11701 4675 11759 4681
rect 11701 4672 11713 4675
rect 11664 4644 11713 4672
rect 11664 4632 11670 4644
rect 11701 4641 11713 4644
rect 11747 4641 11759 4675
rect 12066 4672 12072 4684
rect 12027 4644 12072 4672
rect 11701 4635 11759 4641
rect 12066 4632 12072 4644
rect 12124 4632 12130 4684
rect 13265 4675 13323 4681
rect 13265 4641 13277 4675
rect 13311 4641 13323 4675
rect 13265 4635 13323 4641
rect 13541 4675 13599 4681
rect 13541 4641 13553 4675
rect 13587 4672 13599 4675
rect 13998 4672 14004 4684
rect 13587 4644 14004 4672
rect 13587 4641 13599 4644
rect 13541 4635 13599 4641
rect 12894 4604 12900 4616
rect 6779 4576 11100 4604
rect 12855 4576 12900 4604
rect 6779 4573 6791 4576
rect 6733 4567 6791 4573
rect 12894 4564 12900 4576
rect 12952 4564 12958 4616
rect 13078 4604 13084 4616
rect 13039 4576 13084 4604
rect 13078 4564 13084 4576
rect 13136 4564 13142 4616
rect 13280 4604 13308 4635
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 15212 4672 15240 4712
rect 15746 4700 15752 4712
rect 15804 4700 15810 4752
rect 14108 4644 15240 4672
rect 13722 4604 13728 4616
rect 13280 4576 13728 4604
rect 13722 4564 13728 4576
rect 13780 4604 13786 4616
rect 14108 4604 14136 4644
rect 15470 4632 15476 4684
rect 15528 4672 15534 4684
rect 16209 4675 16267 4681
rect 16209 4672 16221 4675
rect 15528 4644 16221 4672
rect 15528 4632 15534 4644
rect 16209 4641 16221 4644
rect 16255 4641 16267 4675
rect 16209 4635 16267 4641
rect 14826 4604 14832 4616
rect 13780 4576 14136 4604
rect 14787 4576 14832 4604
rect 13780 4564 13786 4576
rect 14826 4564 14832 4576
rect 14884 4564 14890 4616
rect 2317 4471 2375 4477
rect 2317 4437 2329 4471
rect 2363 4468 2375 4471
rect 2777 4471 2835 4477
rect 2777 4468 2789 4471
rect 2363 4440 2789 4468
rect 2363 4437 2375 4440
rect 2317 4431 2375 4437
rect 2777 4437 2789 4440
rect 2823 4468 2835 4471
rect 3142 4468 3148 4480
rect 2823 4440 3148 4468
rect 2823 4437 2835 4440
rect 2777 4431 2835 4437
rect 3142 4428 3148 4440
rect 3200 4428 3206 4480
rect 7374 4468 7380 4480
rect 7335 4440 7380 4468
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 8018 4468 8024 4480
rect 7979 4440 8024 4468
rect 8018 4428 8024 4440
rect 8076 4428 8082 4480
rect 10134 4468 10140 4480
rect 10095 4440 10140 4468
rect 10134 4428 10140 4440
rect 10192 4428 10198 4480
rect 1104 4378 17296 4400
rect 1104 4326 3680 4378
rect 3732 4326 3744 4378
rect 3796 4326 3808 4378
rect 3860 4326 3872 4378
rect 3924 4326 9078 4378
rect 9130 4326 9142 4378
rect 9194 4326 9206 4378
rect 9258 4326 9270 4378
rect 9322 4326 14475 4378
rect 14527 4326 14539 4378
rect 14591 4326 14603 4378
rect 14655 4326 14667 4378
rect 14719 4326 17296 4378
rect 1104 4304 17296 4326
rect 7576 4236 10180 4264
rect 7193 4199 7251 4205
rect 5184 4168 6132 4196
rect 1394 4128 1400 4140
rect 1355 4100 1400 4128
rect 1394 4088 1400 4100
rect 1452 4088 1458 4140
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 2774 4128 2780 4140
rect 2731 4100 2780 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 4430 4088 4436 4140
rect 4488 4128 4494 4140
rect 4709 4131 4767 4137
rect 4709 4128 4721 4131
rect 4488 4100 4721 4128
rect 4488 4088 4494 4100
rect 4709 4097 4721 4100
rect 4755 4128 4767 4131
rect 5184 4128 5212 4168
rect 4755 4100 5212 4128
rect 5261 4131 5319 4137
rect 4755 4097 4767 4100
rect 4709 4091 4767 4097
rect 5261 4097 5273 4131
rect 5307 4128 5319 4131
rect 5534 4128 5540 4140
rect 5307 4100 5540 4128
rect 5307 4097 5319 4100
rect 5261 4091 5319 4097
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 6104 4128 6132 4168
rect 6656 4168 6960 4196
rect 6656 4128 6684 4168
rect 6822 4128 6828 4140
rect 6104 4100 6684 4128
rect 6783 4100 6828 4128
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 6932 4128 6960 4168
rect 7193 4165 7205 4199
rect 7239 4196 7251 4199
rect 7374 4196 7380 4208
rect 7239 4168 7380 4196
rect 7239 4165 7251 4168
rect 7193 4159 7251 4165
rect 7374 4156 7380 4168
rect 7432 4156 7438 4208
rect 7576 4128 7604 4236
rect 7837 4199 7895 4205
rect 7837 4165 7849 4199
rect 7883 4196 7895 4199
rect 7926 4196 7932 4208
rect 7883 4168 7932 4196
rect 7883 4165 7895 4168
rect 7837 4159 7895 4165
rect 7926 4156 7932 4168
rect 7984 4196 7990 4208
rect 9582 4196 9588 4208
rect 7984 4168 9588 4196
rect 7984 4156 7990 4168
rect 9582 4156 9588 4168
rect 9640 4156 9646 4208
rect 10152 4196 10180 4236
rect 15010 4224 15016 4276
rect 15068 4264 15074 4276
rect 16114 4264 16120 4276
rect 15068 4236 16120 4264
rect 15068 4224 15074 4236
rect 16114 4224 16120 4236
rect 16172 4264 16178 4276
rect 16285 4267 16343 4273
rect 16285 4264 16297 4267
rect 16172 4236 16297 4264
rect 16172 4224 16178 4236
rect 16285 4233 16297 4236
rect 16331 4233 16343 4267
rect 16285 4227 16343 4233
rect 12894 4196 12900 4208
rect 10152 4168 10272 4196
rect 8570 4128 8576 4140
rect 6932 4100 7604 4128
rect 8531 4100 8576 4128
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 8941 4131 8999 4137
rect 8941 4097 8953 4131
rect 8987 4128 8999 4131
rect 10134 4128 10140 4140
rect 8987 4100 10140 4128
rect 8987 4097 8999 4100
rect 8941 4091 8999 4097
rect 10134 4088 10140 4100
rect 10192 4088 10198 4140
rect 10244 4128 10272 4168
rect 10980 4168 11284 4196
rect 10980 4128 11008 4168
rect 11146 4128 11152 4140
rect 10244 4100 11008 4128
rect 11107 4100 11152 4128
rect 11146 4088 11152 4100
rect 11204 4088 11210 4140
rect 11256 4128 11284 4168
rect 12728 4168 12900 4196
rect 12728 4137 12756 4168
rect 12894 4156 12900 4168
rect 12952 4156 12958 4208
rect 12529 4131 12587 4137
rect 12529 4128 12541 4131
rect 11256 4100 12541 4128
rect 12529 4097 12541 4100
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 12713 4131 12771 4137
rect 12713 4097 12725 4131
rect 12759 4097 12771 4131
rect 13814 4128 13820 4140
rect 12713 4091 12771 4097
rect 13096 4100 13820 4128
rect 2314 4020 2320 4072
rect 2372 4060 2378 4072
rect 2593 4063 2651 4069
rect 2593 4060 2605 4063
rect 2372 4032 2605 4060
rect 2372 4020 2378 4032
rect 2593 4029 2605 4032
rect 2639 4029 2651 4063
rect 4154 4060 4160 4072
rect 4115 4032 4160 4060
rect 2593 4023 2651 4029
rect 4154 4020 4160 4032
rect 4212 4020 4218 4072
rect 4798 4020 4804 4072
rect 4856 4060 4862 4072
rect 5445 4063 5503 4069
rect 5445 4060 5457 4063
rect 4856 4032 5457 4060
rect 4856 4020 4862 4032
rect 5445 4029 5457 4032
rect 5491 4029 5503 4063
rect 5445 4023 5503 4029
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4060 5687 4063
rect 5902 4060 5908 4072
rect 5675 4032 5908 4060
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 5902 4020 5908 4032
rect 5960 4020 5966 4072
rect 8018 4060 8024 4072
rect 7979 4032 8024 4060
rect 8018 4020 8024 4032
rect 8076 4020 8082 4072
rect 9582 4060 9588 4072
rect 9543 4032 9588 4060
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 10226 4060 10232 4072
rect 10187 4032 10232 4060
rect 10226 4020 10232 4032
rect 10284 4020 10290 4072
rect 10318 4020 10324 4072
rect 10376 4060 10382 4072
rect 13096 4060 13124 4100
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 14553 4131 14611 4137
rect 14553 4097 14565 4131
rect 14599 4128 14611 4131
rect 15010 4128 15016 4140
rect 14599 4100 15016 4128
rect 14599 4097 14611 4100
rect 14553 4091 14611 4097
rect 15010 4088 15016 4100
rect 15068 4088 15074 4140
rect 10376 4032 13124 4060
rect 13725 4063 13783 4069
rect 10376 4020 10382 4032
rect 13725 4029 13737 4063
rect 13771 4029 13783 4063
rect 13725 4023 13783 4029
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 3510 3992 3516 4004
rect 1627 3964 3516 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 3510 3952 3516 3964
rect 3568 3952 3574 4004
rect 8662 3992 8668 4004
rect 6012 3964 8668 3992
rect 1762 3884 1768 3936
rect 1820 3924 1826 3936
rect 6012 3924 6040 3964
rect 8662 3952 8668 3964
rect 8720 3952 8726 4004
rect 8754 3952 8760 4004
rect 8812 3992 8818 4004
rect 8812 3964 10180 3992
rect 8812 3952 8818 3964
rect 7190 3924 7196 3936
rect 1820 3896 6040 3924
rect 7151 3896 7196 3924
rect 1820 3884 1826 3896
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 8018 3884 8024 3936
rect 8076 3924 8082 3936
rect 8941 3927 8999 3933
rect 8941 3924 8953 3927
rect 8076 3896 8953 3924
rect 8076 3884 8082 3896
rect 8941 3893 8953 3896
rect 8987 3893 8999 3927
rect 8941 3887 8999 3893
rect 9030 3884 9036 3936
rect 9088 3924 9094 3936
rect 9401 3927 9459 3933
rect 9401 3924 9413 3927
rect 9088 3896 9413 3924
rect 9088 3884 9094 3896
rect 9401 3893 9413 3896
rect 9447 3893 9459 3927
rect 10042 3924 10048 3936
rect 10003 3896 10048 3924
rect 9401 3887 9459 3893
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10152 3924 10180 3964
rect 10778 3952 10784 4004
rect 10836 3992 10842 4004
rect 10965 3995 11023 4001
rect 10965 3992 10977 3995
rect 10836 3964 10977 3992
rect 10836 3952 10842 3964
rect 10965 3961 10977 3964
rect 11011 3961 11023 3995
rect 12986 3992 12992 4004
rect 10965 3955 11023 3961
rect 11072 3964 12992 3992
rect 11072 3924 11100 3964
rect 12986 3952 12992 3964
rect 13044 3952 13050 4004
rect 13078 3952 13084 4004
rect 13136 3992 13142 4004
rect 13740 3992 13768 4023
rect 13906 4020 13912 4072
rect 13964 4060 13970 4072
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 13964 4032 14289 4060
rect 13964 4020 13970 4032
rect 14277 4029 14289 4032
rect 14323 4029 14335 4063
rect 14277 4023 14335 4029
rect 15654 4020 15660 4072
rect 15712 4020 15718 4072
rect 13136 3964 13768 3992
rect 13136 3952 13142 3964
rect 10152 3896 11100 3924
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 12069 3927 12127 3933
rect 12069 3924 12081 3927
rect 11204 3896 12081 3924
rect 11204 3884 11210 3896
rect 12069 3893 12081 3896
rect 12115 3893 12127 3927
rect 12069 3887 12127 3893
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 13630 3924 13636 3936
rect 12492 3896 12537 3924
rect 13543 3896 13636 3924
rect 12492 3884 12498 3896
rect 13630 3884 13636 3896
rect 13688 3924 13694 3936
rect 16390 3924 16396 3936
rect 13688 3896 16396 3924
rect 13688 3884 13694 3896
rect 16390 3884 16396 3896
rect 16448 3884 16454 3936
rect 1104 3834 17296 3856
rect 1104 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 6571 3834
rect 6623 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 11904 3834
rect 11956 3782 11968 3834
rect 12020 3782 17296 3834
rect 1104 3760 17296 3782
rect 1762 3720 1768 3732
rect 1723 3692 1768 3720
rect 1762 3680 1768 3692
rect 1820 3680 1826 3732
rect 11146 3720 11152 3732
rect 3252 3692 11152 3720
rect 3142 3652 3148 3664
rect 3103 3624 3148 3652
rect 3142 3612 3148 3624
rect 3200 3612 3206 3664
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3553 1639 3587
rect 1581 3547 1639 3553
rect 2374 3587 2432 3593
rect 2374 3553 2386 3587
rect 2420 3584 2432 3587
rect 2682 3584 2688 3596
rect 2420 3556 2688 3584
rect 2420 3553 2432 3556
rect 2374 3547 2432 3553
rect 1596 3516 1624 3547
rect 2682 3544 2688 3556
rect 2740 3544 2746 3596
rect 2774 3516 2780 3528
rect 1596 3488 2780 3516
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 2130 3408 2136 3460
rect 2188 3448 2194 3460
rect 3252 3448 3280 3692
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 11422 3720 11428 3732
rect 11383 3692 11428 3720
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 12492 3692 12537 3720
rect 12492 3680 12498 3692
rect 12986 3680 12992 3732
rect 13044 3720 13050 3732
rect 15654 3720 15660 3732
rect 13044 3692 15660 3720
rect 13044 3680 13050 3692
rect 15654 3680 15660 3692
rect 15712 3680 15718 3732
rect 16025 3723 16083 3729
rect 16025 3689 16037 3723
rect 16071 3689 16083 3723
rect 16025 3683 16083 3689
rect 3326 3612 3332 3664
rect 3384 3652 3390 3664
rect 3384 3624 3429 3652
rect 3384 3612 3390 3624
rect 5626 3612 5632 3664
rect 5684 3652 5690 3664
rect 6914 3652 6920 3664
rect 5684 3624 6920 3652
rect 5684 3612 5690 3624
rect 6914 3612 6920 3624
rect 6972 3612 6978 3664
rect 7466 3652 7472 3664
rect 7427 3624 7472 3652
rect 7466 3612 7472 3624
rect 7524 3612 7530 3664
rect 7745 3655 7803 3661
rect 7745 3621 7757 3655
rect 7791 3652 7803 3655
rect 7926 3652 7932 3664
rect 7791 3624 7932 3652
rect 7791 3621 7803 3624
rect 7745 3615 7803 3621
rect 7926 3612 7932 3624
rect 7984 3612 7990 3664
rect 8386 3612 8392 3664
rect 8444 3652 8450 3664
rect 10226 3652 10232 3664
rect 8444 3624 10232 3652
rect 8444 3612 8450 3624
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 6825 3587 6883 3593
rect 6825 3584 6837 3587
rect 6788 3556 6837 3584
rect 6788 3544 6794 3556
rect 6825 3553 6837 3556
rect 6871 3553 6883 3587
rect 8202 3584 8208 3596
rect 8163 3556 8208 3584
rect 6825 3547 6883 3553
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 8573 3587 8631 3593
rect 8573 3553 8585 3587
rect 8619 3584 8631 3587
rect 9030 3584 9036 3596
rect 8619 3556 9036 3584
rect 8619 3553 8631 3556
rect 8573 3547 8631 3553
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 9490 3584 9496 3596
rect 9451 3556 9496 3584
rect 9490 3544 9496 3556
rect 9548 3544 9554 3596
rect 10060 3593 10088 3624
rect 10226 3612 10232 3624
rect 10284 3612 10290 3664
rect 11330 3652 11336 3664
rect 11291 3624 11336 3652
rect 11330 3612 11336 3624
rect 11388 3612 11394 3664
rect 12897 3655 12955 3661
rect 12897 3652 12909 3655
rect 11440 3624 12909 3652
rect 10045 3587 10103 3593
rect 9692 3556 9996 3584
rect 6089 3519 6147 3525
rect 6089 3485 6101 3519
rect 6135 3516 6147 3519
rect 6135 3488 6316 3516
rect 6135 3485 6147 3488
rect 6089 3479 6147 3485
rect 2188 3420 3280 3448
rect 6288 3448 6316 3488
rect 6362 3476 6368 3528
rect 6420 3516 6426 3528
rect 9692 3516 9720 3556
rect 6420 3488 9720 3516
rect 6420 3476 6426 3488
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9824 3488 9873 3516
rect 9824 3476 9830 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9968 3516 9996 3556
rect 10045 3553 10057 3587
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 11440 3516 11468 3624
rect 12897 3621 12909 3624
rect 12943 3621 12955 3655
rect 12897 3615 12955 3621
rect 13998 3612 14004 3664
rect 14056 3652 14062 3664
rect 14056 3624 15976 3652
rect 14056 3612 14062 3624
rect 12805 3587 12863 3593
rect 12805 3553 12817 3587
rect 12851 3584 12863 3587
rect 13170 3584 13176 3596
rect 12851 3556 13176 3584
rect 12851 3553 12863 3556
rect 12805 3547 12863 3553
rect 13170 3544 13176 3556
rect 13228 3544 13234 3596
rect 13633 3587 13691 3593
rect 13633 3584 13645 3587
rect 13280 3556 13645 3584
rect 11606 3516 11612 3528
rect 9968 3488 11468 3516
rect 11567 3488 11612 3516
rect 9861 3479 9919 3485
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 12986 3516 12992 3528
rect 12947 3488 12992 3516
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 6288 3420 11100 3448
rect 2188 3408 2194 3420
rect 1854 3340 1860 3392
rect 1912 3380 1918 3392
rect 2271 3383 2329 3389
rect 2271 3380 2283 3383
rect 1912 3352 2283 3380
rect 1912 3340 1918 3352
rect 2271 3349 2283 3352
rect 2317 3349 2329 3383
rect 2271 3343 2329 3349
rect 3510 3340 3516 3392
rect 3568 3380 3574 3392
rect 4357 3383 4415 3389
rect 4357 3380 4369 3383
rect 3568 3352 4369 3380
rect 3568 3340 3574 3352
rect 4357 3349 4369 3352
rect 4403 3380 4415 3383
rect 6288 3380 6316 3420
rect 4403 3352 6316 3380
rect 4403 3349 4415 3352
rect 4357 3343 4415 3349
rect 7650 3340 7656 3392
rect 7708 3380 7714 3392
rect 8573 3383 8631 3389
rect 8573 3380 8585 3383
rect 7708 3352 8585 3380
rect 7708 3340 7714 3352
rect 8573 3349 8585 3352
rect 8619 3349 8631 3383
rect 8573 3343 8631 3349
rect 8662 3340 8668 3392
rect 8720 3380 8726 3392
rect 10318 3380 10324 3392
rect 8720 3352 10324 3380
rect 8720 3340 8726 3352
rect 10318 3340 10324 3352
rect 10376 3340 10382 3392
rect 10962 3380 10968 3392
rect 10923 3352 10968 3380
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 11072 3380 11100 3420
rect 12434 3408 12440 3460
rect 12492 3448 12498 3460
rect 13280 3448 13308 3556
rect 13633 3553 13645 3556
rect 13679 3584 13691 3587
rect 13722 3584 13728 3596
rect 13679 3556 13728 3584
rect 13679 3553 13691 3556
rect 13633 3547 13691 3553
rect 13722 3544 13728 3556
rect 13780 3544 13786 3596
rect 15105 3587 15163 3593
rect 15105 3553 15117 3587
rect 15151 3584 15163 3587
rect 15286 3584 15292 3596
rect 15151 3556 15292 3584
rect 15151 3553 15163 3556
rect 15105 3547 15163 3553
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 15948 3593 15976 3624
rect 15933 3587 15991 3593
rect 15933 3553 15945 3587
rect 15979 3553 15991 3587
rect 15933 3547 15991 3553
rect 13906 3516 13912 3528
rect 12492 3420 13308 3448
rect 13464 3488 13912 3516
rect 12492 3408 12498 3420
rect 13464 3380 13492 3488
rect 13906 3476 13912 3488
rect 13964 3476 13970 3528
rect 15010 3476 15016 3528
rect 15068 3516 15074 3528
rect 15197 3519 15255 3525
rect 15197 3516 15209 3519
rect 15068 3488 15209 3516
rect 15068 3476 15074 3488
rect 15197 3485 15209 3488
rect 15243 3485 15255 3519
rect 15197 3479 15255 3485
rect 15381 3519 15439 3525
rect 15381 3485 15393 3519
rect 15427 3516 15439 3519
rect 16040 3516 16068 3683
rect 16209 3587 16267 3593
rect 16209 3553 16221 3587
rect 16255 3553 16267 3587
rect 16390 3584 16396 3596
rect 16351 3556 16396 3584
rect 16209 3547 16267 3553
rect 15427 3488 16068 3516
rect 15427 3485 15439 3488
rect 15381 3479 15439 3485
rect 13725 3451 13783 3457
rect 13725 3417 13737 3451
rect 13771 3448 13783 3451
rect 14274 3448 14280 3460
rect 13771 3420 14280 3448
rect 13771 3417 13783 3420
rect 13725 3411 13783 3417
rect 14274 3408 14280 3420
rect 14332 3448 14338 3460
rect 16224 3448 16252 3547
rect 16390 3544 16396 3556
rect 16448 3544 16454 3596
rect 14332 3420 16252 3448
rect 14332 3408 14338 3420
rect 11072 3352 13492 3380
rect 13814 3340 13820 3392
rect 13872 3380 13878 3392
rect 14737 3383 14795 3389
rect 14737 3380 14749 3383
rect 13872 3352 14749 3380
rect 13872 3340 13878 3352
rect 14737 3349 14749 3352
rect 14783 3349 14795 3383
rect 14737 3343 14795 3349
rect 1104 3290 17296 3312
rect 1104 3238 3680 3290
rect 3732 3238 3744 3290
rect 3796 3238 3808 3290
rect 3860 3238 3872 3290
rect 3924 3238 9078 3290
rect 9130 3238 9142 3290
rect 9194 3238 9206 3290
rect 9258 3238 9270 3290
rect 9322 3238 14475 3290
rect 14527 3238 14539 3290
rect 14591 3238 14603 3290
rect 14655 3238 14667 3290
rect 14719 3238 17296 3290
rect 1104 3216 17296 3238
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 6086 3176 6092 3188
rect 5592 3148 6092 3176
rect 5592 3136 5598 3148
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 6178 3136 6184 3188
rect 6236 3176 6242 3188
rect 8662 3176 8668 3188
rect 6236 3148 8668 3176
rect 6236 3136 6242 3148
rect 8662 3136 8668 3148
rect 8720 3136 8726 3188
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 9585 3179 9643 3185
rect 9585 3176 9597 3179
rect 9548 3148 9597 3176
rect 9548 3136 9554 3148
rect 9585 3145 9597 3148
rect 9631 3145 9643 3179
rect 10778 3176 10784 3188
rect 10739 3148 10784 3176
rect 9585 3139 9643 3145
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 13170 3176 13176 3188
rect 13131 3148 13176 3176
rect 13170 3136 13176 3148
rect 13228 3136 13234 3188
rect 5169 3111 5227 3117
rect 5169 3077 5181 3111
rect 5215 3108 5227 3111
rect 5215 3080 10824 3108
rect 5215 3077 5227 3080
rect 5169 3071 5227 3077
rect 1578 3000 1584 3052
rect 1636 3040 1642 3052
rect 1765 3043 1823 3049
rect 1765 3040 1777 3043
rect 1636 3012 1777 3040
rect 1636 3000 1642 3012
rect 1765 3009 1777 3012
rect 1811 3040 1823 3043
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 1811 3012 2513 3040
rect 1811 3009 1823 3012
rect 1765 3003 1823 3009
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 5813 3043 5871 3049
rect 4212 3012 4660 3040
rect 4212 3000 4218 3012
rect 1854 2972 1860 2984
rect 1815 2944 1860 2972
rect 1854 2932 1860 2944
rect 1912 2932 1918 2984
rect 4632 2972 4660 3012
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 8846 3040 8852 3052
rect 5859 3012 7604 3040
rect 8807 3012 8852 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 6178 2972 6184 2984
rect 4632 2944 6184 2972
rect 6178 2932 6184 2944
rect 6236 2932 6242 2984
rect 6730 2932 6736 2984
rect 6788 2972 6794 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6788 2944 6837 2972
rect 6788 2932 6794 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 7466 2972 7472 2984
rect 7427 2944 7472 2972
rect 6825 2935 6883 2941
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 7576 2981 7604 3012
rect 8846 3000 8852 3012
rect 8904 3000 8910 3052
rect 8938 3000 8944 3052
rect 8996 3040 9002 3052
rect 9033 3043 9091 3049
rect 9033 3040 9045 3043
rect 8996 3012 9045 3040
rect 8996 3000 9002 3012
rect 9033 3009 9045 3012
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2941 7619 2975
rect 9048 2972 9076 3003
rect 9950 3000 9956 3052
rect 10008 3040 10014 3052
rect 10796 3049 10824 3080
rect 10045 3043 10103 3049
rect 10045 3040 10057 3043
rect 10008 3012 10057 3040
rect 10008 3000 10014 3012
rect 10045 3009 10057 3012
rect 10091 3009 10103 3043
rect 10045 3003 10103 3009
rect 10137 3043 10195 3049
rect 10137 3009 10149 3043
rect 10183 3009 10195 3043
rect 10137 3003 10195 3009
rect 10781 3043 10839 3049
rect 10781 3009 10793 3043
rect 10827 3009 10839 3043
rect 10781 3003 10839 3009
rect 10152 2972 10180 3003
rect 10962 3000 10968 3052
rect 11020 3040 11026 3052
rect 11149 3043 11207 3049
rect 11149 3040 11161 3043
rect 11020 3012 11161 3040
rect 11020 3000 11026 3012
rect 11149 3009 11161 3012
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 12253 3043 12311 3049
rect 12253 3009 12265 3043
rect 12299 3040 12311 3043
rect 13630 3040 13636 3052
rect 12299 3012 13636 3040
rect 12299 3009 12311 3012
rect 12253 3003 12311 3009
rect 13630 3000 13636 3012
rect 13688 3000 13694 3052
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3040 13783 3043
rect 14182 3040 14188 3052
rect 13771 3012 14188 3040
rect 13771 3009 13783 3012
rect 13725 3003 13783 3009
rect 14182 3000 14188 3012
rect 14240 3000 14246 3052
rect 14369 3043 14427 3049
rect 14369 3009 14381 3043
rect 14415 3040 14427 3043
rect 15010 3040 15016 3052
rect 14415 3012 15016 3040
rect 14415 3009 14427 3012
rect 14369 3003 14427 3009
rect 15010 3000 15016 3012
rect 15068 3000 15074 3052
rect 9048 2944 10180 2972
rect 7561 2935 7619 2941
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12713 2975 12771 2981
rect 12492 2944 12537 2972
rect 12492 2932 12498 2944
rect 12713 2941 12725 2975
rect 12759 2941 12771 2975
rect 12713 2935 12771 2941
rect 13541 2975 13599 2981
rect 13541 2941 13553 2975
rect 13587 2972 13599 2975
rect 13814 2972 13820 2984
rect 13587 2944 13820 2972
rect 13587 2941 13599 2944
rect 13541 2935 13599 2941
rect 2777 2907 2835 2913
rect 2777 2873 2789 2907
rect 2823 2904 2835 2907
rect 5074 2904 5080 2916
rect 2823 2876 3004 2904
rect 4002 2876 5080 2904
rect 2823 2873 2835 2876
rect 2777 2867 2835 2873
rect 2976 2848 3004 2876
rect 5074 2864 5080 2876
rect 5132 2864 5138 2916
rect 5261 2907 5319 2913
rect 5261 2873 5273 2907
rect 5307 2904 5319 2907
rect 9766 2904 9772 2916
rect 5307 2876 7420 2904
rect 5307 2873 5319 2876
rect 5261 2867 5319 2873
rect 2958 2796 2964 2848
rect 3016 2836 3022 2848
rect 4501 2839 4559 2845
rect 4501 2836 4513 2839
rect 3016 2808 4513 2836
rect 3016 2796 3022 2808
rect 4501 2805 4513 2808
rect 4547 2836 4559 2839
rect 5810 2836 5816 2848
rect 4547 2808 5816 2836
rect 4547 2805 4559 2808
rect 4501 2799 4559 2805
rect 5810 2796 5816 2808
rect 5868 2796 5874 2848
rect 5905 2839 5963 2845
rect 5905 2805 5917 2839
rect 5951 2836 5963 2839
rect 7190 2836 7196 2848
rect 5951 2808 7196 2836
rect 5951 2805 5963 2808
rect 5905 2799 5963 2805
rect 7190 2796 7196 2808
rect 7248 2796 7254 2848
rect 7392 2836 7420 2876
rect 7760 2876 9772 2904
rect 7760 2836 7788 2876
rect 9766 2864 9772 2876
rect 9824 2864 9830 2916
rect 9858 2864 9864 2916
rect 9916 2904 9922 2916
rect 9953 2907 10011 2913
rect 9953 2904 9965 2907
rect 9916 2876 9965 2904
rect 9916 2864 9922 2876
rect 9953 2873 9965 2876
rect 9999 2873 10011 2907
rect 9953 2867 10011 2873
rect 10134 2864 10140 2916
rect 10192 2864 10198 2916
rect 12728 2904 12756 2935
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 15654 2932 15660 2984
rect 15712 2972 15718 2984
rect 15712 2944 15778 2972
rect 15712 2932 15718 2944
rect 13633 2907 13691 2913
rect 12728 2876 13584 2904
rect 7392 2808 7788 2836
rect 7834 2796 7840 2848
rect 7892 2836 7898 2848
rect 8202 2836 8208 2848
rect 7892 2808 8208 2836
rect 7892 2796 7898 2808
rect 8202 2796 8208 2808
rect 8260 2836 8266 2848
rect 8389 2839 8447 2845
rect 8389 2836 8401 2839
rect 8260 2808 8401 2836
rect 8260 2796 8266 2808
rect 8389 2805 8401 2808
rect 8435 2805 8447 2839
rect 8389 2799 8447 2805
rect 8757 2839 8815 2845
rect 8757 2805 8769 2839
rect 8803 2836 8815 2839
rect 10152 2836 10180 2864
rect 8803 2808 10180 2836
rect 12621 2839 12679 2845
rect 8803 2805 8815 2808
rect 8757 2799 8815 2805
rect 12621 2805 12633 2839
rect 12667 2836 12679 2839
rect 12986 2836 12992 2848
rect 12667 2808 12992 2836
rect 12667 2805 12679 2808
rect 12621 2799 12679 2805
rect 12986 2796 12992 2808
rect 13044 2796 13050 2848
rect 13556 2836 13584 2876
rect 13633 2873 13645 2907
rect 13679 2904 13691 2907
rect 13906 2904 13912 2916
rect 13679 2876 13912 2904
rect 13679 2873 13691 2876
rect 13633 2867 13691 2873
rect 13906 2864 13912 2876
rect 13964 2864 13970 2916
rect 14645 2907 14703 2913
rect 14645 2873 14657 2907
rect 14691 2873 14703 2907
rect 14645 2867 14703 2873
rect 13814 2836 13820 2848
rect 13556 2808 13820 2836
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 14660 2836 14688 2867
rect 15286 2836 15292 2848
rect 14660 2808 15292 2836
rect 15286 2796 15292 2808
rect 15344 2836 15350 2848
rect 16390 2836 16396 2848
rect 15344 2808 16396 2836
rect 15344 2796 15350 2808
rect 16390 2796 16396 2808
rect 16448 2796 16454 2848
rect 1104 2746 17296 2768
rect 1104 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 6571 2746
rect 6623 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 11904 2746
rect 11956 2694 11968 2746
rect 12020 2694 17296 2746
rect 1104 2672 17296 2694
rect 2222 2632 2228 2644
rect 2183 2604 2228 2632
rect 2222 2592 2228 2604
rect 2280 2592 2286 2644
rect 2777 2635 2835 2641
rect 2777 2601 2789 2635
rect 2823 2601 2835 2635
rect 2777 2595 2835 2601
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 4246 2632 4252 2644
rect 4203 2604 4252 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 1578 2564 1584 2576
rect 1539 2536 1584 2564
rect 1578 2524 1584 2536
rect 1636 2524 1642 2576
rect 2317 2499 2375 2505
rect 2317 2465 2329 2499
rect 2363 2496 2375 2499
rect 2792 2496 2820 2595
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 5074 2632 5080 2644
rect 4987 2604 5080 2632
rect 5074 2592 5080 2604
rect 5132 2632 5138 2644
rect 5626 2632 5632 2644
rect 5132 2604 5632 2632
rect 5132 2592 5138 2604
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 6270 2592 6276 2644
rect 6328 2632 6334 2644
rect 6641 2635 6699 2641
rect 6641 2632 6653 2635
rect 6328 2604 6653 2632
rect 6328 2592 6334 2604
rect 6641 2601 6653 2604
rect 6687 2601 6699 2635
rect 6641 2595 6699 2601
rect 9766 2592 9772 2644
rect 9824 2632 9830 2644
rect 9953 2635 10011 2641
rect 9953 2632 9965 2635
rect 9824 2604 9965 2632
rect 9824 2592 9830 2604
rect 9953 2601 9965 2604
rect 9999 2601 10011 2635
rect 13906 2632 13912 2644
rect 13867 2604 13912 2632
rect 9953 2595 10011 2601
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 14918 2592 14924 2644
rect 14976 2632 14982 2644
rect 15013 2635 15071 2641
rect 15013 2632 15025 2635
rect 14976 2604 15025 2632
rect 14976 2592 14982 2604
rect 15013 2601 15025 2604
rect 15059 2601 15071 2635
rect 15654 2632 15660 2644
rect 15615 2604 15660 2632
rect 15013 2595 15071 2601
rect 15654 2592 15660 2604
rect 15712 2592 15718 2644
rect 7926 2564 7932 2576
rect 7300 2536 7932 2564
rect 2363 2468 2820 2496
rect 2961 2499 3019 2505
rect 2363 2465 2375 2468
rect 2317 2459 2375 2465
rect 2961 2465 2973 2499
rect 3007 2465 3019 2499
rect 2961 2459 3019 2465
rect 474 2388 480 2440
rect 532 2428 538 2440
rect 2976 2428 3004 2459
rect 3050 2456 3056 2508
rect 3108 2496 3114 2508
rect 4341 2499 4399 2505
rect 4341 2496 4353 2499
rect 3108 2468 4353 2496
rect 3108 2456 3114 2468
rect 4341 2465 4353 2468
rect 4387 2465 4399 2499
rect 4341 2459 4399 2465
rect 4798 2456 4804 2508
rect 4856 2496 4862 2508
rect 7300 2505 7328 2536
rect 7926 2524 7932 2536
rect 7984 2524 7990 2576
rect 10505 2567 10563 2573
rect 10505 2533 10517 2567
rect 10551 2564 10563 2567
rect 10778 2564 10784 2576
rect 10551 2536 10784 2564
rect 10551 2533 10563 2536
rect 10505 2527 10563 2533
rect 10778 2524 10784 2536
rect 10836 2524 10842 2576
rect 11606 2524 11612 2576
rect 11664 2564 11670 2576
rect 12802 2564 12808 2576
rect 11664 2536 12808 2564
rect 11664 2524 11670 2536
rect 12802 2524 12808 2536
rect 12860 2564 12866 2576
rect 12897 2567 12955 2573
rect 12897 2564 12909 2567
rect 12860 2536 12909 2564
rect 12860 2524 12866 2536
rect 12897 2533 12909 2536
rect 12943 2564 12955 2567
rect 14826 2564 14832 2576
rect 12943 2536 14832 2564
rect 12943 2533 12955 2536
rect 12897 2527 12955 2533
rect 14826 2524 14832 2536
rect 14884 2524 14890 2576
rect 15102 2524 15108 2576
rect 15160 2564 15166 2576
rect 16390 2564 16396 2576
rect 15160 2536 15884 2564
rect 16351 2536 16396 2564
rect 15160 2524 15166 2536
rect 4893 2499 4951 2505
rect 4893 2496 4905 2499
rect 4856 2468 4905 2496
rect 4856 2456 4862 2468
rect 4893 2465 4905 2468
rect 4939 2465 4951 2499
rect 4893 2459 4951 2465
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2465 5871 2499
rect 5813 2459 5871 2465
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2496 6607 2499
rect 6825 2499 6883 2505
rect 6825 2496 6837 2499
rect 6595 2468 6837 2496
rect 6595 2465 6607 2468
rect 6549 2459 6607 2465
rect 6825 2465 6837 2468
rect 6871 2465 6883 2499
rect 6825 2459 6883 2465
rect 7285 2499 7343 2505
rect 7285 2465 7297 2499
rect 7331 2465 7343 2499
rect 7834 2496 7840 2508
rect 7795 2468 7840 2496
rect 7285 2459 7343 2465
rect 532 2400 3004 2428
rect 5828 2428 5856 2459
rect 7834 2456 7840 2468
rect 7892 2456 7898 2508
rect 8294 2456 8300 2508
rect 8352 2496 8358 2508
rect 8389 2499 8447 2505
rect 8389 2496 8401 2499
rect 8352 2468 8401 2496
rect 8352 2456 8358 2468
rect 8389 2465 8401 2468
rect 8435 2465 8447 2499
rect 8389 2459 8447 2465
rect 9490 2456 9496 2508
rect 9548 2496 9554 2508
rect 9585 2499 9643 2505
rect 9585 2496 9597 2499
rect 9548 2468 9597 2496
rect 9548 2456 9554 2468
rect 9585 2465 9597 2468
rect 9631 2465 9643 2499
rect 9585 2459 9643 2465
rect 9953 2499 10011 2505
rect 9953 2465 9965 2499
rect 9999 2496 10011 2499
rect 10042 2496 10048 2508
rect 9999 2468 10048 2496
rect 9999 2465 10011 2468
rect 9953 2459 10011 2465
rect 10042 2456 10048 2468
rect 10100 2456 10106 2508
rect 10134 2456 10140 2508
rect 10192 2496 10198 2508
rect 10413 2499 10471 2505
rect 10413 2496 10425 2499
rect 10192 2468 10425 2496
rect 10192 2456 10198 2468
rect 10413 2465 10425 2468
rect 10459 2465 10471 2499
rect 10962 2496 10968 2508
rect 10923 2468 10968 2496
rect 10413 2459 10471 2465
rect 10962 2456 10968 2468
rect 11020 2456 11026 2508
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 12529 2499 12587 2505
rect 12529 2496 12541 2499
rect 12492 2468 12541 2496
rect 12492 2456 12498 2468
rect 12529 2465 12541 2468
rect 12575 2465 12587 2499
rect 13814 2496 13820 2508
rect 13775 2468 13820 2496
rect 12529 2459 12587 2465
rect 13814 2456 13820 2468
rect 13872 2456 13878 2508
rect 15197 2499 15255 2505
rect 15197 2465 15209 2499
rect 15243 2496 15255 2499
rect 15746 2496 15752 2508
rect 15243 2468 15752 2496
rect 15243 2465 15255 2468
rect 15197 2459 15255 2465
rect 15746 2456 15752 2468
rect 15804 2456 15810 2508
rect 15856 2505 15884 2536
rect 16390 2524 16396 2536
rect 16448 2524 16454 2576
rect 15841 2499 15899 2505
rect 15841 2465 15853 2499
rect 15887 2465 15899 2499
rect 15841 2459 15899 2465
rect 6914 2428 6920 2440
rect 5828 2400 6920 2428
rect 532 2388 538 2400
rect 6914 2388 6920 2400
rect 6972 2388 6978 2440
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7248 2400 7481 2428
rect 7248 2388 7254 2400
rect 7469 2397 7481 2400
rect 7515 2428 7527 2431
rect 7650 2428 7656 2440
rect 7515 2400 7656 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 13078 2428 13084 2440
rect 8619 2400 13084 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 13078 2388 13084 2400
rect 13136 2388 13142 2440
rect 1394 2360 1400 2372
rect 1355 2332 1400 2360
rect 1394 2320 1400 2332
rect 1452 2320 1458 2372
rect 5997 2363 6055 2369
rect 5997 2329 6009 2363
rect 6043 2360 6055 2363
rect 7742 2360 7748 2372
rect 6043 2332 7748 2360
rect 6043 2329 6055 2332
rect 5997 2323 6055 2329
rect 7742 2320 7748 2332
rect 7800 2320 7806 2372
rect 16574 2320 16580 2372
rect 16632 2360 16638 2372
rect 16632 2332 16677 2360
rect 16632 2320 16638 2332
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 6549 2295 6607 2301
rect 6549 2292 6561 2295
rect 1360 2264 6561 2292
rect 1360 2252 1366 2264
rect 6549 2261 6561 2264
rect 6595 2261 6607 2295
rect 6549 2255 6607 2261
rect 1104 2202 17296 2224
rect 1104 2150 3680 2202
rect 3732 2150 3744 2202
rect 3796 2150 3808 2202
rect 3860 2150 3872 2202
rect 3924 2150 9078 2202
rect 9130 2150 9142 2202
rect 9194 2150 9206 2202
rect 9258 2150 9270 2202
rect 9322 2150 14475 2202
rect 14527 2150 14539 2202
rect 14591 2150 14603 2202
rect 14655 2150 14667 2202
rect 14719 2150 17296 2202
rect 1104 2128 17296 2150
<< via1 >>
rect 2320 18028 2372 18080
rect 8760 18028 8812 18080
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 6571 17926 6623 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 11904 17926 11956 17978
rect 11968 17926 12020 17978
rect 1492 17867 1544 17876
rect 1492 17833 1501 17867
rect 1501 17833 1535 17867
rect 1535 17833 1544 17867
rect 1492 17824 1544 17833
rect 3424 17824 3476 17876
rect 6000 17756 6052 17808
rect 1768 17620 1820 17672
rect 5356 17620 5408 17672
rect 5540 17688 5592 17740
rect 15660 17824 15712 17876
rect 7656 17731 7708 17740
rect 7656 17697 7665 17731
rect 7665 17697 7699 17731
rect 7699 17697 7708 17731
rect 7656 17688 7708 17697
rect 8484 17731 8536 17740
rect 8484 17697 8493 17731
rect 8493 17697 8527 17731
rect 8527 17697 8536 17731
rect 8484 17688 8536 17697
rect 9588 17731 9640 17740
rect 9588 17697 9597 17731
rect 9597 17697 9631 17731
rect 9631 17697 9640 17731
rect 9588 17688 9640 17697
rect 9772 17731 9824 17740
rect 9772 17697 9781 17731
rect 9781 17697 9815 17731
rect 9815 17697 9824 17731
rect 9772 17688 9824 17697
rect 14280 17756 14332 17808
rect 14924 17756 14976 17808
rect 17040 17756 17092 17808
rect 5724 17620 5776 17672
rect 12440 17620 12492 17672
rect 13084 17620 13136 17672
rect 14832 17731 14884 17740
rect 14832 17697 14841 17731
rect 14841 17697 14875 17731
rect 14875 17697 14884 17731
rect 14832 17688 14884 17697
rect 16028 17688 16080 17740
rect 15568 17620 15620 17672
rect 5632 17552 5684 17604
rect 4804 17527 4856 17536
rect 4804 17493 4813 17527
rect 4813 17493 4847 17527
rect 4847 17493 4856 17527
rect 4804 17484 4856 17493
rect 5264 17527 5316 17536
rect 5264 17493 5273 17527
rect 5273 17493 5307 17527
rect 5307 17493 5316 17527
rect 5264 17484 5316 17493
rect 7840 17527 7892 17536
rect 7840 17493 7849 17527
rect 7849 17493 7883 17527
rect 7883 17493 7892 17527
rect 7840 17484 7892 17493
rect 8392 17527 8444 17536
rect 8392 17493 8401 17527
rect 8401 17493 8435 17527
rect 8435 17493 8444 17527
rect 8392 17484 8444 17493
rect 9680 17527 9732 17536
rect 9680 17493 9689 17527
rect 9689 17493 9723 17527
rect 9723 17493 9732 17527
rect 9680 17484 9732 17493
rect 15108 17552 15160 17604
rect 16120 17552 16172 17604
rect 11060 17484 11112 17536
rect 11336 17527 11388 17536
rect 11336 17493 11345 17527
rect 11345 17493 11379 17527
rect 11379 17493 11388 17527
rect 11336 17484 11388 17493
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 13176 17527 13228 17536
rect 13176 17493 13185 17527
rect 13185 17493 13219 17527
rect 13219 17493 13228 17527
rect 13176 17484 13228 17493
rect 15016 17527 15068 17536
rect 15016 17493 15025 17527
rect 15025 17493 15059 17527
rect 15059 17493 15068 17527
rect 15016 17484 15068 17493
rect 15752 17527 15804 17536
rect 15752 17493 15761 17527
rect 15761 17493 15795 17527
rect 15795 17493 15804 17527
rect 15752 17484 15804 17493
rect 3680 17382 3732 17434
rect 3744 17382 3796 17434
rect 3808 17382 3860 17434
rect 3872 17382 3924 17434
rect 9078 17382 9130 17434
rect 9142 17382 9194 17434
rect 9206 17382 9258 17434
rect 9270 17382 9322 17434
rect 14475 17382 14527 17434
rect 14539 17382 14591 17434
rect 14603 17382 14655 17434
rect 14667 17382 14719 17434
rect 6920 17280 6972 17332
rect 10416 17280 10468 17332
rect 12532 17280 12584 17332
rect 2964 17212 3016 17264
rect 5724 17212 5776 17264
rect 1768 17119 1820 17128
rect 1768 17085 1777 17119
rect 1777 17085 1811 17119
rect 1811 17085 1820 17119
rect 1768 17076 1820 17085
rect 3332 17144 3384 17196
rect 5264 17144 5316 17196
rect 15016 17144 15068 17196
rect 1676 17008 1728 17060
rect 3056 17076 3108 17128
rect 3424 17119 3476 17128
rect 3424 17085 3433 17119
rect 3433 17085 3467 17119
rect 3467 17085 3476 17119
rect 3424 17076 3476 17085
rect 5356 17076 5408 17128
rect 7656 17076 7708 17128
rect 7840 17076 7892 17128
rect 10416 17119 10468 17128
rect 2872 17008 2924 17060
rect 1952 16983 2004 16992
rect 1952 16949 1961 16983
rect 1961 16949 1995 16983
rect 1995 16949 2004 16983
rect 1952 16940 2004 16949
rect 10416 17085 10425 17119
rect 10425 17085 10459 17119
rect 10459 17085 10468 17119
rect 10416 17076 10468 17085
rect 10508 17119 10560 17128
rect 10508 17085 10517 17119
rect 10517 17085 10551 17119
rect 10551 17085 10560 17119
rect 10508 17076 10560 17085
rect 10876 17076 10928 17128
rect 14372 17119 14424 17128
rect 14372 17085 14381 17119
rect 14381 17085 14415 17119
rect 14415 17085 14424 17119
rect 14372 17076 14424 17085
rect 7564 16940 7616 16992
rect 9864 17008 9916 17060
rect 11152 17008 11204 17060
rect 13176 17008 13228 17060
rect 15108 17008 15160 17060
rect 12256 16940 12308 16992
rect 14832 16940 14884 16992
rect 15384 16940 15436 16992
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 6571 16838 6623 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 11904 16838 11956 16890
rect 11968 16838 12020 16890
rect 9772 16779 9824 16788
rect 1676 16711 1728 16720
rect 1676 16677 1685 16711
rect 1685 16677 1719 16711
rect 1719 16677 1728 16711
rect 1676 16668 1728 16677
rect 1952 16668 2004 16720
rect 2964 16668 3016 16720
rect 5724 16668 5776 16720
rect 9772 16745 9781 16779
rect 9781 16745 9815 16779
rect 9815 16745 9824 16779
rect 9772 16736 9824 16745
rect 7564 16668 7616 16720
rect 11152 16711 11204 16720
rect 11152 16677 11161 16711
rect 11161 16677 11195 16711
rect 11195 16677 11204 16711
rect 11152 16668 11204 16677
rect 3332 16600 3384 16652
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 6092 16532 6144 16584
rect 5540 16464 5592 16516
rect 6000 16464 6052 16516
rect 3056 16396 3108 16448
rect 9864 16600 9916 16652
rect 10508 16600 10560 16652
rect 10968 16600 11020 16652
rect 9956 16575 10008 16584
rect 9956 16541 9965 16575
rect 9965 16541 9999 16575
rect 9999 16541 10008 16575
rect 9956 16532 10008 16541
rect 10416 16575 10468 16584
rect 10416 16541 10425 16575
rect 10425 16541 10459 16575
rect 10459 16541 10468 16575
rect 10416 16532 10468 16541
rect 12256 16736 12308 16788
rect 13084 16736 13136 16788
rect 11336 16668 11388 16720
rect 11244 16643 11296 16652
rect 11244 16609 11253 16643
rect 11253 16609 11287 16643
rect 11287 16609 11296 16643
rect 11428 16643 11480 16652
rect 11244 16600 11296 16609
rect 11428 16609 11437 16643
rect 11437 16609 11471 16643
rect 11471 16609 11480 16643
rect 11428 16600 11480 16609
rect 12716 16643 12768 16652
rect 12716 16609 12725 16643
rect 12725 16609 12759 16643
rect 12759 16609 12768 16643
rect 12716 16600 12768 16609
rect 12808 16600 12860 16652
rect 12164 16532 12216 16584
rect 14372 16532 14424 16584
rect 15384 16532 15436 16584
rect 10232 16464 10284 16516
rect 12348 16464 12400 16516
rect 12440 16464 12492 16516
rect 6920 16396 6972 16448
rect 8024 16439 8076 16448
rect 8024 16405 8033 16439
rect 8033 16405 8067 16439
rect 8067 16405 8076 16439
rect 8024 16396 8076 16405
rect 10140 16396 10192 16448
rect 11520 16396 11572 16448
rect 13452 16396 13504 16448
rect 16488 16439 16540 16448
rect 16488 16405 16497 16439
rect 16497 16405 16531 16439
rect 16531 16405 16540 16439
rect 16488 16396 16540 16405
rect 3680 16294 3732 16346
rect 3744 16294 3796 16346
rect 3808 16294 3860 16346
rect 3872 16294 3924 16346
rect 9078 16294 9130 16346
rect 9142 16294 9194 16346
rect 9206 16294 9258 16346
rect 9270 16294 9322 16346
rect 14475 16294 14527 16346
rect 14539 16294 14591 16346
rect 14603 16294 14655 16346
rect 14667 16294 14719 16346
rect 2872 16235 2924 16244
rect 2872 16201 2881 16235
rect 2881 16201 2915 16235
rect 2915 16201 2924 16235
rect 2872 16192 2924 16201
rect 8300 16192 8352 16244
rect 9772 16192 9824 16244
rect 1860 15988 1912 16040
rect 3424 16056 3476 16108
rect 4252 16056 4304 16108
rect 3056 15988 3108 16040
rect 480 15920 532 15972
rect 1308 15920 1360 15972
rect 4160 15963 4212 15972
rect 4160 15929 4169 15963
rect 4169 15929 4203 15963
rect 4203 15929 4212 15963
rect 4160 15920 4212 15929
rect 4804 15920 4856 15972
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 9588 16124 9640 16176
rect 6092 16056 6144 16108
rect 6276 16056 6328 16108
rect 5724 15988 5776 16040
rect 7288 16031 7340 16040
rect 6184 15920 6236 15972
rect 7288 15997 7297 16031
rect 7297 15997 7331 16031
rect 7331 15997 7340 16031
rect 7288 15988 7340 15997
rect 8668 16099 8720 16108
rect 8024 15988 8076 16040
rect 8668 16065 8677 16099
rect 8677 16065 8711 16099
rect 8711 16065 8720 16099
rect 8668 16056 8720 16065
rect 9680 16056 9732 16108
rect 11428 16192 11480 16244
rect 12716 16192 12768 16244
rect 13176 16192 13228 16244
rect 8484 16031 8536 16040
rect 8484 15997 8493 16031
rect 8493 15997 8527 16031
rect 8527 15997 8536 16031
rect 9772 16031 9824 16040
rect 8484 15988 8536 15997
rect 9772 15997 9781 16031
rect 9781 15997 9815 16031
rect 9815 15997 9824 16031
rect 9772 15988 9824 15997
rect 11244 16124 11296 16176
rect 6092 15852 6144 15904
rect 13912 16056 13964 16108
rect 10968 16031 11020 16040
rect 10968 15997 10977 16031
rect 10977 15997 11011 16031
rect 11011 15997 11020 16031
rect 10968 15988 11020 15997
rect 10692 15920 10744 15972
rect 11244 15852 11296 15904
rect 15200 15988 15252 16040
rect 16488 16124 16540 16176
rect 12716 15963 12768 15972
rect 12716 15929 12725 15963
rect 12725 15929 12759 15963
rect 12759 15929 12768 15963
rect 12716 15920 12768 15929
rect 13452 15920 13504 15972
rect 15016 15920 15068 15972
rect 16580 15988 16632 16040
rect 14372 15852 14424 15904
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 6571 15750 6623 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 11904 15750 11956 15802
rect 11968 15750 12020 15802
rect 1676 15648 1728 15700
rect 4160 15648 4212 15700
rect 1768 15512 1820 15564
rect 5724 15580 5776 15632
rect 6184 15623 6236 15632
rect 2872 15555 2924 15564
rect 2872 15521 2881 15555
rect 2881 15521 2915 15555
rect 2915 15521 2924 15555
rect 2872 15512 2924 15521
rect 3976 15512 4028 15564
rect 6184 15589 6193 15623
rect 6193 15589 6227 15623
rect 6227 15589 6236 15623
rect 6184 15580 6236 15589
rect 6000 15555 6052 15564
rect 6000 15521 6009 15555
rect 6009 15521 6043 15555
rect 6043 15521 6052 15555
rect 6000 15512 6052 15521
rect 2780 15444 2832 15496
rect 3332 15444 3384 15496
rect 6920 15512 6972 15564
rect 7196 15555 7248 15564
rect 6276 15444 6328 15496
rect 7196 15521 7205 15555
rect 7205 15521 7239 15555
rect 7239 15521 7248 15555
rect 7196 15512 7248 15521
rect 2964 15376 3016 15428
rect 7380 15444 7432 15496
rect 2136 15308 2188 15360
rect 2228 15308 2280 15360
rect 4344 15351 4396 15360
rect 4344 15317 4353 15351
rect 4353 15317 4387 15351
rect 4387 15317 4396 15351
rect 4344 15308 4396 15317
rect 6736 15376 6788 15428
rect 9772 15648 9824 15700
rect 10416 15691 10468 15700
rect 10416 15657 10425 15691
rect 10425 15657 10459 15691
rect 10459 15657 10468 15691
rect 10416 15648 10468 15657
rect 10600 15648 10652 15700
rect 10876 15648 10928 15700
rect 12716 15691 12768 15700
rect 9956 15580 10008 15632
rect 10232 15623 10284 15632
rect 10232 15589 10241 15623
rect 10241 15589 10275 15623
rect 10275 15589 10284 15623
rect 10232 15580 10284 15589
rect 8116 15444 8168 15496
rect 8300 15512 8352 15564
rect 11612 15580 11664 15632
rect 12716 15657 12725 15691
rect 12725 15657 12759 15691
rect 12759 15657 12768 15691
rect 12716 15648 12768 15657
rect 16580 15691 16632 15700
rect 16580 15657 16589 15691
rect 16589 15657 16623 15691
rect 16623 15657 16632 15691
rect 16580 15648 16632 15657
rect 12164 15555 12216 15564
rect 8668 15444 8720 15496
rect 8760 15376 8812 15428
rect 9680 15376 9732 15428
rect 12164 15521 12173 15555
rect 12173 15521 12207 15555
rect 12207 15521 12216 15555
rect 12164 15512 12216 15521
rect 13084 15580 13136 15632
rect 15200 15580 15252 15632
rect 15568 15580 15620 15632
rect 12440 15512 12492 15564
rect 13176 15512 13228 15564
rect 13268 15512 13320 15564
rect 13820 15555 13872 15564
rect 13820 15521 13829 15555
rect 13829 15521 13863 15555
rect 13863 15521 13872 15555
rect 13820 15512 13872 15521
rect 13084 15444 13136 15496
rect 14372 15444 14424 15496
rect 6276 15308 6328 15360
rect 10692 15308 10744 15360
rect 13636 15308 13688 15360
rect 3680 15206 3732 15258
rect 3744 15206 3796 15258
rect 3808 15206 3860 15258
rect 3872 15206 3924 15258
rect 9078 15206 9130 15258
rect 9142 15206 9194 15258
rect 9206 15206 9258 15258
rect 9270 15206 9322 15258
rect 14475 15206 14527 15258
rect 14539 15206 14591 15258
rect 14603 15206 14655 15258
rect 14667 15206 14719 15258
rect 2780 15036 2832 15088
rect 2228 14968 2280 15020
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 3976 14968 4028 15020
rect 7196 15104 7248 15156
rect 9956 15104 10008 15156
rect 13268 15104 13320 15156
rect 7288 15036 7340 15088
rect 5172 14968 5224 15020
rect 10968 15036 11020 15088
rect 11060 15036 11112 15088
rect 14924 15104 14976 15156
rect 2136 14832 2188 14884
rect 4344 14900 4396 14952
rect 5632 14900 5684 14952
rect 6736 14900 6788 14952
rect 6920 14943 6972 14952
rect 6920 14909 6929 14943
rect 6929 14909 6963 14943
rect 6963 14909 6972 14943
rect 6920 14900 6972 14909
rect 8392 14943 8444 14952
rect 8392 14909 8401 14943
rect 8401 14909 8435 14943
rect 8435 14909 8444 14943
rect 8392 14900 8444 14909
rect 9772 14968 9824 15020
rect 9956 14968 10008 15020
rect 8760 14943 8812 14952
rect 8760 14909 8769 14943
rect 8769 14909 8803 14943
rect 8803 14909 8812 14943
rect 8760 14900 8812 14909
rect 7932 14875 7984 14884
rect 7932 14841 7941 14875
rect 7941 14841 7975 14875
rect 7975 14841 7984 14875
rect 7932 14832 7984 14841
rect 8024 14832 8076 14884
rect 9680 14900 9732 14952
rect 10324 14943 10376 14952
rect 10324 14909 10330 14943
rect 10330 14909 10364 14943
rect 10364 14909 10376 14943
rect 10324 14900 10376 14909
rect 10692 14943 10744 14952
rect 10692 14909 10701 14943
rect 10701 14909 10735 14943
rect 10735 14909 10744 14943
rect 10692 14900 10744 14909
rect 12624 14900 12676 14952
rect 13820 15036 13872 15088
rect 13636 15011 13688 15020
rect 13636 14977 13645 15011
rect 13645 14977 13679 15011
rect 13679 14977 13688 15011
rect 13636 14968 13688 14977
rect 3332 14764 3384 14816
rect 4160 14764 4212 14816
rect 5080 14764 5132 14816
rect 10232 14764 10284 14816
rect 12440 14832 12492 14884
rect 13912 14900 13964 14952
rect 14924 14943 14976 14952
rect 14924 14909 14933 14943
rect 14933 14909 14967 14943
rect 14967 14909 14976 14943
rect 14924 14900 14976 14909
rect 15108 14943 15160 14952
rect 15108 14909 15117 14943
rect 15117 14909 15151 14943
rect 15151 14909 15160 14943
rect 15108 14900 15160 14909
rect 15936 14900 15988 14952
rect 16212 14832 16264 14884
rect 13176 14764 13228 14816
rect 15108 14764 15160 14816
rect 15844 14807 15896 14816
rect 15844 14773 15853 14807
rect 15853 14773 15887 14807
rect 15887 14773 15896 14807
rect 15844 14764 15896 14773
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 6571 14662 6623 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 11904 14662 11956 14714
rect 11968 14662 12020 14714
rect 2780 14560 2832 14612
rect 2964 14603 3016 14612
rect 2964 14569 2973 14603
rect 2973 14569 3007 14603
rect 3007 14569 3016 14603
rect 2964 14560 3016 14569
rect 3332 14535 3384 14544
rect 1768 14424 1820 14476
rect 3332 14501 3341 14535
rect 3341 14501 3375 14535
rect 3375 14501 3384 14535
rect 3332 14492 3384 14501
rect 3056 14424 3108 14476
rect 1952 14356 2004 14408
rect 8024 14560 8076 14612
rect 8760 14560 8812 14612
rect 10324 14560 10376 14612
rect 8392 14535 8444 14544
rect 8392 14501 8401 14535
rect 8401 14501 8435 14535
rect 8435 14501 8444 14535
rect 8392 14492 8444 14501
rect 10968 14535 11020 14544
rect 10968 14501 10977 14535
rect 10977 14501 11011 14535
rect 11011 14501 11020 14535
rect 10968 14492 11020 14501
rect 8024 14424 8076 14476
rect 8208 14467 8260 14476
rect 8208 14433 8217 14467
rect 8217 14433 8251 14467
rect 8251 14433 8260 14467
rect 8208 14424 8260 14433
rect 9956 14467 10008 14476
rect 9956 14433 9965 14467
rect 9965 14433 9999 14467
rect 9999 14433 10008 14467
rect 9956 14424 10008 14433
rect 10232 14467 10284 14476
rect 10232 14433 10241 14467
rect 10241 14433 10275 14467
rect 10275 14433 10284 14467
rect 10232 14424 10284 14433
rect 12440 14603 12492 14612
rect 12440 14569 12449 14603
rect 12449 14569 12483 14603
rect 12483 14569 12492 14603
rect 12440 14560 12492 14569
rect 13176 14560 13228 14612
rect 12532 14492 12584 14544
rect 15936 14560 15988 14612
rect 16212 14560 16264 14612
rect 4252 14356 4304 14408
rect 5264 14356 5316 14408
rect 7196 14356 7248 14408
rect 8484 14356 8536 14408
rect 9864 14356 9916 14408
rect 11336 14356 11388 14408
rect 12440 14424 12492 14476
rect 12624 14424 12676 14476
rect 13084 14467 13136 14476
rect 13084 14433 13093 14467
rect 13093 14433 13127 14467
rect 13127 14433 13136 14467
rect 13084 14424 13136 14433
rect 13176 14467 13228 14476
rect 13176 14433 13185 14467
rect 13185 14433 13219 14467
rect 13219 14433 13228 14467
rect 14832 14492 14884 14544
rect 13176 14424 13228 14433
rect 12348 14356 12400 14408
rect 14280 14424 14332 14476
rect 15016 14424 15068 14476
rect 14096 14356 14148 14408
rect 4988 14220 5040 14272
rect 6092 14220 6144 14272
rect 7380 14263 7432 14272
rect 7380 14229 7389 14263
rect 7389 14229 7423 14263
rect 7423 14229 7432 14263
rect 7380 14220 7432 14229
rect 9772 14263 9824 14272
rect 9772 14229 9781 14263
rect 9781 14229 9815 14263
rect 9815 14229 9824 14263
rect 9772 14220 9824 14229
rect 11152 14220 11204 14272
rect 14740 14288 14792 14340
rect 15660 14424 15712 14476
rect 15844 14424 15896 14476
rect 16304 14424 16356 14476
rect 16488 14356 16540 14408
rect 12624 14220 12676 14272
rect 14924 14263 14976 14272
rect 14924 14229 14933 14263
rect 14933 14229 14967 14263
rect 14967 14229 14976 14263
rect 14924 14220 14976 14229
rect 3680 14118 3732 14170
rect 3744 14118 3796 14170
rect 3808 14118 3860 14170
rect 3872 14118 3924 14170
rect 9078 14118 9130 14170
rect 9142 14118 9194 14170
rect 9206 14118 9258 14170
rect 9270 14118 9322 14170
rect 14475 14118 14527 14170
rect 14539 14118 14591 14170
rect 14603 14118 14655 14170
rect 14667 14118 14719 14170
rect 3240 14016 3292 14068
rect 2596 13948 2648 14000
rect 5080 14016 5132 14068
rect 5264 14059 5316 14068
rect 5264 14025 5273 14059
rect 5273 14025 5307 14059
rect 5307 14025 5316 14059
rect 5264 14016 5316 14025
rect 6736 14016 6788 14068
rect 7932 14016 7984 14068
rect 8116 14059 8168 14068
rect 8116 14025 8125 14059
rect 8125 14025 8159 14059
rect 8159 14025 8168 14059
rect 8116 14016 8168 14025
rect 9772 14016 9824 14068
rect 10968 14016 11020 14068
rect 14096 14059 14148 14068
rect 14096 14025 14105 14059
rect 14105 14025 14139 14059
rect 14139 14025 14148 14059
rect 14096 14016 14148 14025
rect 15936 14016 15988 14068
rect 4344 13948 4396 14000
rect 5908 13948 5960 14000
rect 8208 13948 8260 14000
rect 3976 13880 4028 13932
rect 3516 13855 3568 13864
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 3516 13812 3568 13821
rect 2780 13676 2832 13728
rect 2964 13744 3016 13796
rect 4068 13812 4120 13864
rect 4344 13855 4396 13864
rect 4344 13821 4353 13855
rect 4353 13821 4387 13855
rect 4387 13821 4396 13855
rect 4344 13812 4396 13821
rect 3332 13719 3384 13728
rect 3332 13685 3341 13719
rect 3341 13685 3375 13719
rect 3375 13685 3384 13719
rect 3332 13676 3384 13685
rect 4160 13744 4212 13796
rect 6000 13812 6052 13864
rect 4620 13676 4672 13728
rect 5632 13787 5684 13796
rect 5632 13753 5641 13787
rect 5641 13753 5675 13787
rect 5675 13753 5684 13787
rect 5632 13744 5684 13753
rect 6092 13744 6144 13796
rect 7196 13880 7248 13932
rect 11060 13948 11112 14000
rect 11336 13948 11388 14000
rect 8392 13923 8444 13932
rect 8392 13889 8401 13923
rect 8401 13889 8435 13923
rect 8435 13889 8444 13923
rect 8760 13923 8812 13932
rect 8392 13880 8444 13889
rect 8760 13889 8769 13923
rect 8769 13889 8803 13923
rect 8803 13889 8812 13923
rect 8760 13880 8812 13889
rect 10692 13880 10744 13932
rect 10968 13855 11020 13864
rect 10968 13821 10977 13855
rect 10977 13821 11011 13855
rect 11011 13821 11020 13855
rect 10968 13812 11020 13821
rect 7012 13744 7064 13796
rect 10232 13744 10284 13796
rect 12624 13923 12676 13932
rect 12624 13889 12633 13923
rect 12633 13889 12667 13923
rect 12667 13889 12676 13923
rect 12624 13880 12676 13889
rect 14924 13923 14976 13932
rect 14924 13889 14933 13923
rect 14933 13889 14967 13923
rect 14967 13889 14976 13923
rect 14924 13880 14976 13889
rect 14372 13812 14424 13864
rect 12532 13744 12584 13796
rect 16212 13744 16264 13796
rect 7656 13676 7708 13728
rect 9772 13676 9824 13728
rect 12440 13676 12492 13728
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 6571 13574 6623 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 11904 13574 11956 13626
rect 11968 13574 12020 13626
rect 2872 13472 2924 13524
rect 4252 13515 4304 13524
rect 4252 13481 4261 13515
rect 4261 13481 4295 13515
rect 4295 13481 4304 13515
rect 4252 13472 4304 13481
rect 7196 13515 7248 13524
rect 7196 13481 7205 13515
rect 7205 13481 7239 13515
rect 7239 13481 7248 13515
rect 7196 13472 7248 13481
rect 7932 13515 7984 13524
rect 7932 13481 7941 13515
rect 7941 13481 7975 13515
rect 7975 13481 7984 13515
rect 7932 13472 7984 13481
rect 10692 13515 10744 13524
rect 10692 13481 10701 13515
rect 10701 13481 10735 13515
rect 10735 13481 10744 13515
rect 10692 13472 10744 13481
rect 10876 13515 10928 13524
rect 10876 13481 10885 13515
rect 10885 13481 10919 13515
rect 10919 13481 10928 13515
rect 10876 13472 10928 13481
rect 10968 13472 11020 13524
rect 3516 13404 3568 13456
rect 4804 13404 4856 13456
rect 7104 13404 7156 13456
rect 7656 13404 7708 13456
rect 1768 13336 1820 13388
rect 2780 13336 2832 13388
rect 3056 13379 3108 13388
rect 3056 13345 3065 13379
rect 3065 13345 3099 13379
rect 3099 13345 3108 13379
rect 4620 13379 4672 13388
rect 3056 13336 3108 13345
rect 3608 13268 3660 13320
rect 4620 13345 4629 13379
rect 4629 13345 4663 13379
rect 4663 13345 4672 13379
rect 4620 13336 4672 13345
rect 5080 13379 5132 13388
rect 5080 13345 5089 13379
rect 5089 13345 5123 13379
rect 5123 13345 5132 13379
rect 5080 13336 5132 13345
rect 5908 13336 5960 13388
rect 6092 13379 6144 13388
rect 6092 13345 6101 13379
rect 6101 13345 6135 13379
rect 6135 13345 6144 13379
rect 6092 13336 6144 13345
rect 6736 13336 6788 13388
rect 7012 13379 7064 13388
rect 5632 13268 5684 13320
rect 7012 13345 7021 13379
rect 7021 13345 7055 13379
rect 7055 13345 7064 13379
rect 7012 13336 7064 13345
rect 8208 13379 8260 13388
rect 8208 13345 8217 13379
rect 8217 13345 8251 13379
rect 8251 13345 8260 13379
rect 8208 13336 8260 13345
rect 12440 13404 12492 13456
rect 11612 13336 11664 13388
rect 12164 13336 12216 13388
rect 12348 13336 12400 13388
rect 13084 13472 13136 13524
rect 15016 13515 15068 13524
rect 15016 13481 15025 13515
rect 15025 13481 15059 13515
rect 15059 13481 15068 13515
rect 15016 13472 15068 13481
rect 13176 13404 13228 13456
rect 13268 13336 13320 13388
rect 15752 13404 15804 13456
rect 16304 13472 16356 13524
rect 15844 13379 15896 13388
rect 2228 13175 2280 13184
rect 2228 13141 2237 13175
rect 2237 13141 2271 13175
rect 2271 13141 2280 13175
rect 2228 13132 2280 13141
rect 2688 13175 2740 13184
rect 2688 13141 2697 13175
rect 2697 13141 2731 13175
rect 2731 13141 2740 13175
rect 2688 13132 2740 13141
rect 2964 13200 3016 13252
rect 4344 13200 4396 13252
rect 7840 13268 7892 13320
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 11336 13311 11388 13320
rect 11336 13277 11345 13311
rect 11345 13277 11379 13311
rect 11379 13277 11388 13311
rect 11336 13268 11388 13277
rect 12808 13268 12860 13320
rect 15844 13345 15853 13379
rect 15853 13345 15887 13379
rect 15887 13345 15896 13379
rect 15844 13336 15896 13345
rect 15568 13268 15620 13320
rect 5908 13200 5960 13252
rect 6184 13200 6236 13252
rect 7380 13200 7432 13252
rect 14832 13200 14884 13252
rect 16488 13336 16540 13388
rect 5816 13175 5868 13184
rect 5816 13141 5825 13175
rect 5825 13141 5859 13175
rect 5859 13141 5868 13175
rect 5816 13132 5868 13141
rect 6736 13132 6788 13184
rect 7196 13132 7248 13184
rect 11060 13132 11112 13184
rect 11796 13175 11848 13184
rect 11796 13141 11805 13175
rect 11805 13141 11839 13175
rect 11839 13141 11848 13175
rect 11796 13132 11848 13141
rect 13176 13175 13228 13184
rect 13176 13141 13185 13175
rect 13185 13141 13219 13175
rect 13219 13141 13228 13175
rect 13176 13132 13228 13141
rect 3680 13030 3732 13082
rect 3744 13030 3796 13082
rect 3808 13030 3860 13082
rect 3872 13030 3924 13082
rect 9078 13030 9130 13082
rect 9142 13030 9194 13082
rect 9206 13030 9258 13082
rect 9270 13030 9322 13082
rect 14475 13030 14527 13082
rect 14539 13030 14591 13082
rect 14603 13030 14655 13082
rect 14667 13030 14719 13082
rect 1400 12928 1452 12980
rect 3240 12928 3292 12980
rect 3516 12928 3568 12980
rect 7012 12928 7064 12980
rect 7840 12971 7892 12980
rect 7840 12937 7849 12971
rect 7849 12937 7883 12971
rect 7883 12937 7892 12971
rect 7840 12928 7892 12937
rect 11060 12971 11112 12980
rect 11060 12937 11069 12971
rect 11069 12937 11103 12971
rect 11103 12937 11112 12971
rect 11060 12928 11112 12937
rect 11336 12928 11388 12980
rect 13820 12928 13872 12980
rect 14832 12928 14884 12980
rect 16212 12971 16264 12980
rect 16212 12937 16221 12971
rect 16221 12937 16255 12971
rect 16255 12937 16264 12971
rect 16212 12928 16264 12937
rect 4988 12860 5040 12912
rect 5632 12860 5684 12912
rect 8116 12860 8168 12912
rect 2688 12792 2740 12844
rect 3148 12792 3200 12844
rect 3516 12792 3568 12844
rect 4804 12835 4856 12844
rect 4804 12801 4813 12835
rect 4813 12801 4847 12835
rect 4847 12801 4856 12835
rect 4804 12792 4856 12801
rect 6000 12792 6052 12844
rect 7932 12792 7984 12844
rect 10876 12792 10928 12844
rect 13636 12792 13688 12844
rect 3332 12724 3384 12776
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 4620 12724 4672 12733
rect 4712 12767 4764 12776
rect 4712 12733 4721 12767
rect 4721 12733 4755 12767
rect 4755 12733 4764 12767
rect 5080 12767 5132 12776
rect 4712 12724 4764 12733
rect 5080 12733 5089 12767
rect 5089 12733 5123 12767
rect 5123 12733 5132 12767
rect 5080 12724 5132 12733
rect 2228 12656 2280 12708
rect 6736 12724 6788 12776
rect 7380 12767 7432 12776
rect 7380 12733 7387 12767
rect 7387 12733 7432 12767
rect 7380 12724 7432 12733
rect 7656 12767 7708 12776
rect 7656 12733 7670 12767
rect 7670 12733 7704 12767
rect 7704 12733 7708 12767
rect 7656 12724 7708 12733
rect 7472 12699 7524 12708
rect 7472 12665 7481 12699
rect 7481 12665 7515 12699
rect 7515 12665 7524 12699
rect 7472 12656 7524 12665
rect 10784 12724 10836 12776
rect 12072 12767 12124 12776
rect 12072 12733 12081 12767
rect 12081 12733 12115 12767
rect 12115 12733 12124 12767
rect 12072 12724 12124 12733
rect 12256 12767 12308 12776
rect 12256 12733 12265 12767
rect 12265 12733 12299 12767
rect 12299 12733 12308 12767
rect 12256 12724 12308 12733
rect 12992 12767 13044 12776
rect 12992 12733 13001 12767
rect 13001 12733 13035 12767
rect 13035 12733 13044 12767
rect 12992 12724 13044 12733
rect 13176 12724 13228 12776
rect 14096 12724 14148 12776
rect 15384 12767 15436 12776
rect 15384 12733 15393 12767
rect 15393 12733 15427 12767
rect 15427 12733 15436 12767
rect 15384 12724 15436 12733
rect 15568 12767 15620 12776
rect 15568 12733 15577 12767
rect 15577 12733 15611 12767
rect 15611 12733 15620 12767
rect 15568 12724 15620 12733
rect 15752 12767 15804 12776
rect 15752 12733 15761 12767
rect 15761 12733 15795 12767
rect 15795 12733 15804 12767
rect 15752 12724 15804 12733
rect 16304 12724 16356 12776
rect 3332 12588 3384 12640
rect 8484 12656 8536 12708
rect 11796 12656 11848 12708
rect 13728 12699 13780 12708
rect 13728 12665 13737 12699
rect 13737 12665 13771 12699
rect 13771 12665 13780 12699
rect 13728 12656 13780 12665
rect 15476 12699 15528 12708
rect 15476 12665 15485 12699
rect 15485 12665 15519 12699
rect 15519 12665 15528 12699
rect 15476 12656 15528 12665
rect 7840 12588 7892 12640
rect 9496 12588 9548 12640
rect 12716 12631 12768 12640
rect 12716 12597 12725 12631
rect 12725 12597 12759 12631
rect 12759 12597 12768 12631
rect 12716 12588 12768 12597
rect 14096 12631 14148 12640
rect 14096 12597 14105 12631
rect 14105 12597 14139 12631
rect 14139 12597 14148 12631
rect 14096 12588 14148 12597
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 6571 12486 6623 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 11904 12486 11956 12538
rect 11968 12486 12020 12538
rect 3976 12384 4028 12436
rect 4252 12384 4304 12436
rect 2320 12316 2372 12368
rect 2044 12248 2096 12300
rect 3148 12291 3200 12300
rect 3148 12257 3157 12291
rect 3157 12257 3191 12291
rect 3191 12257 3200 12291
rect 3148 12248 3200 12257
rect 3332 12291 3384 12300
rect 3332 12257 3341 12291
rect 3341 12257 3375 12291
rect 3375 12257 3384 12291
rect 3332 12248 3384 12257
rect 4068 12112 4120 12164
rect 4712 12248 4764 12300
rect 5356 12248 5408 12300
rect 7288 12384 7340 12436
rect 7472 12427 7524 12436
rect 7472 12393 7481 12427
rect 7481 12393 7515 12427
rect 7515 12393 7524 12427
rect 7472 12384 7524 12393
rect 8668 12384 8720 12436
rect 6092 12316 6144 12368
rect 6644 12316 6696 12368
rect 6552 12291 6604 12300
rect 6552 12257 6561 12291
rect 6561 12257 6595 12291
rect 6595 12257 6604 12291
rect 6552 12248 6604 12257
rect 5080 12180 5132 12232
rect 7840 12316 7892 12368
rect 11336 12316 11388 12368
rect 7196 12248 7248 12300
rect 7656 12291 7708 12300
rect 7656 12257 7665 12291
rect 7665 12257 7699 12291
rect 7699 12257 7708 12291
rect 7656 12248 7708 12257
rect 7380 12180 7432 12232
rect 8208 12248 8260 12300
rect 9496 12291 9548 12300
rect 9496 12257 9505 12291
rect 9505 12257 9539 12291
rect 9539 12257 9548 12291
rect 9496 12248 9548 12257
rect 10784 12248 10836 12300
rect 5632 12112 5684 12164
rect 6368 12155 6420 12164
rect 6368 12121 6377 12155
rect 6377 12121 6411 12155
rect 6411 12121 6420 12155
rect 6368 12112 6420 12121
rect 6552 12112 6604 12164
rect 7472 12112 7524 12164
rect 11612 12248 11664 12300
rect 12256 12384 12308 12436
rect 12072 12291 12124 12300
rect 12072 12257 12081 12291
rect 12081 12257 12115 12291
rect 12115 12257 12124 12291
rect 12072 12248 12124 12257
rect 12716 12248 12768 12300
rect 13268 12316 13320 12368
rect 13176 12248 13228 12300
rect 15108 12384 15160 12436
rect 15384 12359 15436 12368
rect 15384 12325 15393 12359
rect 15393 12325 15427 12359
rect 15427 12325 15436 12359
rect 15384 12316 15436 12325
rect 15936 12316 15988 12368
rect 14280 12248 14332 12300
rect 15476 12291 15528 12300
rect 15476 12257 15485 12291
rect 15485 12257 15519 12291
rect 15519 12257 15528 12291
rect 15476 12248 15528 12257
rect 15660 12291 15712 12300
rect 15660 12257 15669 12291
rect 15669 12257 15703 12291
rect 15703 12257 15712 12291
rect 15660 12248 15712 12257
rect 16580 12291 16632 12300
rect 16580 12257 16589 12291
rect 16589 12257 16623 12291
rect 16623 12257 16632 12291
rect 16580 12248 16632 12257
rect 12808 12112 12860 12164
rect 14280 12112 14332 12164
rect 2228 12044 2280 12096
rect 2780 12044 2832 12096
rect 4252 12044 4304 12096
rect 4620 12044 4672 12096
rect 5816 12087 5868 12096
rect 5816 12053 5825 12087
rect 5825 12053 5859 12087
rect 5859 12053 5868 12087
rect 5816 12044 5868 12053
rect 6184 12044 6236 12096
rect 7748 12044 7800 12096
rect 12624 12087 12676 12096
rect 12624 12053 12633 12087
rect 12633 12053 12667 12087
rect 12667 12053 12676 12087
rect 12624 12044 12676 12053
rect 13084 12044 13136 12096
rect 13636 12044 13688 12096
rect 15108 12087 15160 12096
rect 15108 12053 15117 12087
rect 15117 12053 15151 12087
rect 15151 12053 15160 12087
rect 15108 12044 15160 12053
rect 3680 11942 3732 11994
rect 3744 11942 3796 11994
rect 3808 11942 3860 11994
rect 3872 11942 3924 11994
rect 9078 11942 9130 11994
rect 9142 11942 9194 11994
rect 9206 11942 9258 11994
rect 9270 11942 9322 11994
rect 14475 11942 14527 11994
rect 14539 11942 14591 11994
rect 14603 11942 14655 11994
rect 14667 11942 14719 11994
rect 4160 11840 4212 11892
rect 4528 11840 4580 11892
rect 4896 11840 4948 11892
rect 5356 11883 5408 11892
rect 5356 11849 5365 11883
rect 5365 11849 5399 11883
rect 5399 11849 5408 11883
rect 5356 11840 5408 11849
rect 6184 11840 6236 11892
rect 12532 11840 12584 11892
rect 2320 11704 2372 11756
rect 4160 11636 4212 11688
rect 4528 11704 4580 11756
rect 4620 11679 4672 11688
rect 2504 11568 2556 11620
rect 2596 11568 2648 11620
rect 4620 11645 4629 11679
rect 4629 11645 4663 11679
rect 4663 11645 4672 11679
rect 4620 11636 4672 11645
rect 13268 11772 13320 11824
rect 13728 11840 13780 11892
rect 15752 11840 15804 11892
rect 15844 11840 15896 11892
rect 16120 11840 16172 11892
rect 13820 11772 13872 11824
rect 5080 11704 5132 11756
rect 7380 11704 7432 11756
rect 12992 11747 13044 11756
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 14004 11747 14056 11756
rect 12992 11704 13044 11713
rect 5908 11679 5960 11688
rect 5356 11568 5408 11620
rect 5908 11645 5917 11679
rect 5917 11645 5951 11679
rect 5951 11645 5960 11679
rect 5908 11636 5960 11645
rect 6736 11636 6788 11688
rect 7012 11679 7064 11688
rect 7012 11645 7019 11679
rect 7019 11645 7064 11679
rect 7012 11636 7064 11645
rect 7288 11679 7340 11688
rect 7288 11645 7302 11679
rect 7302 11645 7336 11679
rect 7336 11645 7340 11679
rect 8484 11679 8536 11688
rect 7288 11636 7340 11645
rect 8484 11645 8493 11679
rect 8493 11645 8527 11679
rect 8527 11645 8536 11679
rect 8484 11636 8536 11645
rect 12164 11636 12216 11688
rect 13084 11679 13136 11688
rect 13084 11645 13093 11679
rect 13093 11645 13127 11679
rect 13127 11645 13136 11679
rect 14004 11713 14013 11747
rect 14013 11713 14047 11747
rect 14047 11713 14056 11747
rect 14004 11704 14056 11713
rect 13084 11636 13136 11645
rect 5816 11568 5868 11620
rect 6368 11568 6420 11620
rect 8760 11611 8812 11620
rect 2412 11500 2464 11552
rect 4896 11543 4948 11552
rect 4896 11509 4905 11543
rect 4905 11509 4939 11543
rect 4939 11509 4948 11543
rect 4896 11500 4948 11509
rect 6184 11500 6236 11552
rect 8760 11577 8769 11611
rect 8769 11577 8803 11611
rect 8803 11577 8812 11611
rect 8760 11568 8812 11577
rect 13820 11636 13872 11688
rect 14280 11679 14332 11688
rect 14280 11645 14289 11679
rect 14289 11645 14323 11679
rect 14323 11645 14332 11679
rect 14280 11636 14332 11645
rect 15476 11704 15528 11756
rect 15936 11679 15988 11688
rect 15936 11645 15945 11679
rect 15945 11645 15979 11679
rect 15979 11645 15988 11679
rect 15936 11636 15988 11645
rect 16028 11679 16080 11688
rect 16028 11645 16037 11679
rect 16037 11645 16071 11679
rect 16071 11645 16080 11679
rect 16028 11636 16080 11645
rect 8024 11500 8076 11552
rect 10232 11543 10284 11552
rect 10232 11509 10241 11543
rect 10241 11509 10275 11543
rect 10275 11509 10284 11543
rect 10232 11500 10284 11509
rect 15936 11500 15988 11552
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 6571 11398 6623 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 11904 11398 11956 11450
rect 11968 11398 12020 11450
rect 2596 11296 2648 11348
rect 7196 11296 7248 11348
rect 7472 11296 7524 11348
rect 4160 11228 4212 11280
rect 2044 11203 2096 11212
rect 2044 11169 2053 11203
rect 2053 11169 2087 11203
rect 2087 11169 2096 11203
rect 2044 11160 2096 11169
rect 2504 11203 2556 11212
rect 2504 11169 2513 11203
rect 2513 11169 2547 11203
rect 2547 11169 2556 11203
rect 2504 11160 2556 11169
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 7196 11160 7248 11169
rect 7380 11160 7432 11212
rect 2136 11092 2188 11144
rect 4528 11135 4580 11144
rect 4528 11101 4537 11135
rect 4537 11101 4571 11135
rect 4571 11101 4580 11135
rect 4528 11092 4580 11101
rect 7748 11228 7800 11280
rect 8760 11296 8812 11348
rect 10876 11296 10928 11348
rect 11612 11296 11664 11348
rect 8116 11160 8168 11212
rect 8484 11228 8536 11280
rect 9956 11228 10008 11280
rect 12072 11228 12124 11280
rect 12808 11228 12860 11280
rect 15936 11296 15988 11348
rect 15108 11271 15160 11280
rect 15108 11237 15117 11271
rect 15117 11237 15151 11271
rect 15151 11237 15160 11271
rect 15108 11228 15160 11237
rect 14372 11160 14424 11212
rect 16212 11160 16264 11212
rect 8024 11135 8076 11144
rect 7288 11024 7340 11076
rect 4344 10956 4396 11008
rect 4988 10956 5040 11008
rect 5816 10956 5868 11008
rect 6828 10956 6880 11008
rect 8024 11101 8033 11135
rect 8033 11101 8067 11135
rect 8067 11101 8076 11135
rect 8024 11092 8076 11101
rect 9864 11135 9916 11144
rect 9864 11101 9873 11135
rect 9873 11101 9907 11135
rect 9907 11101 9916 11135
rect 9864 11092 9916 11101
rect 9956 11092 10008 11144
rect 12624 11092 12676 11144
rect 14372 11024 14424 11076
rect 3680 10854 3732 10906
rect 3744 10854 3796 10906
rect 3808 10854 3860 10906
rect 3872 10854 3924 10906
rect 9078 10854 9130 10906
rect 9142 10854 9194 10906
rect 9206 10854 9258 10906
rect 9270 10854 9322 10906
rect 14475 10854 14527 10906
rect 14539 10854 14591 10906
rect 14603 10854 14655 10906
rect 14667 10854 14719 10906
rect 2136 10795 2188 10804
rect 2136 10761 2145 10795
rect 2145 10761 2179 10795
rect 2179 10761 2188 10795
rect 2136 10752 2188 10761
rect 4160 10752 4212 10804
rect 4528 10752 4580 10804
rect 6184 10752 6236 10804
rect 7104 10752 7156 10804
rect 9864 10752 9916 10804
rect 12072 10795 12124 10804
rect 12072 10761 12081 10795
rect 12081 10761 12115 10795
rect 12115 10761 12124 10795
rect 12072 10752 12124 10761
rect 12808 10752 12860 10804
rect 2780 10727 2832 10736
rect 2780 10693 2789 10727
rect 2789 10693 2823 10727
rect 2823 10693 2832 10727
rect 2780 10684 2832 10693
rect 1952 10616 2004 10668
rect 3148 10659 3200 10668
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 3056 10548 3108 10600
rect 4896 10616 4948 10668
rect 5540 10616 5592 10668
rect 6276 10616 6328 10668
rect 8668 10659 8720 10668
rect 8668 10625 8677 10659
rect 8677 10625 8711 10659
rect 8711 10625 8720 10659
rect 8668 10616 8720 10625
rect 8760 10659 8812 10668
rect 8760 10625 8769 10659
rect 8769 10625 8803 10659
rect 8803 10625 8812 10659
rect 8760 10616 8812 10625
rect 1768 10455 1820 10464
rect 1768 10421 1777 10455
rect 1777 10421 1811 10455
rect 1811 10421 1820 10455
rect 1768 10412 1820 10421
rect 2412 10412 2464 10464
rect 2964 10480 3016 10532
rect 3976 10548 4028 10600
rect 5632 10548 5684 10600
rect 5816 10548 5868 10600
rect 6736 10548 6788 10600
rect 10232 10548 10284 10600
rect 10968 10616 11020 10668
rect 14096 10659 14148 10668
rect 14096 10625 14105 10659
rect 14105 10625 14139 10659
rect 14139 10625 14148 10659
rect 14096 10616 14148 10625
rect 16028 10616 16080 10668
rect 5540 10412 5592 10464
rect 5908 10412 5960 10464
rect 6184 10412 6236 10464
rect 8576 10455 8628 10464
rect 8576 10421 8585 10455
rect 8585 10421 8619 10455
rect 8619 10421 8628 10455
rect 8576 10412 8628 10421
rect 9680 10412 9732 10464
rect 10600 10480 10652 10532
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 11152 10591 11204 10600
rect 10876 10548 10928 10557
rect 11152 10557 11161 10591
rect 11161 10557 11195 10591
rect 11195 10557 11204 10591
rect 11152 10548 11204 10557
rect 12164 10548 12216 10600
rect 13360 10548 13412 10600
rect 11612 10480 11664 10532
rect 14372 10480 14424 10532
rect 14832 10480 14884 10532
rect 12440 10412 12492 10464
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 6571 10310 6623 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 11904 10310 11956 10362
rect 11968 10310 12020 10362
rect 1492 10251 1544 10260
rect 1492 10217 1501 10251
rect 1501 10217 1535 10251
rect 1535 10217 1544 10251
rect 1492 10208 1544 10217
rect 1768 10208 1820 10260
rect 7380 10208 7432 10260
rect 7840 10208 7892 10260
rect 8576 10208 8628 10260
rect 9864 10208 9916 10260
rect 2412 10140 2464 10192
rect 4068 10140 4120 10192
rect 2044 10072 2096 10124
rect 2596 10115 2648 10124
rect 2596 10081 2605 10115
rect 2605 10081 2639 10115
rect 2639 10081 2648 10115
rect 2596 10072 2648 10081
rect 3148 10115 3200 10124
rect 3148 10081 3157 10115
rect 3157 10081 3191 10115
rect 3191 10081 3200 10115
rect 3148 10072 3200 10081
rect 2964 10004 3016 10056
rect 7196 10072 7248 10124
rect 7380 10115 7432 10124
rect 7380 10081 7389 10115
rect 7389 10081 7423 10115
rect 7423 10081 7432 10115
rect 7380 10072 7432 10081
rect 7472 10115 7524 10124
rect 7472 10081 7481 10115
rect 7481 10081 7515 10115
rect 7515 10081 7524 10115
rect 9404 10140 9456 10192
rect 7472 10072 7524 10081
rect 6184 10004 6236 10056
rect 5632 9936 5684 9988
rect 6828 10004 6880 10056
rect 7656 10004 7708 10056
rect 8300 10072 8352 10124
rect 9956 10072 10008 10124
rect 10600 10140 10652 10192
rect 14832 10208 14884 10260
rect 15844 10208 15896 10260
rect 16212 10208 16264 10260
rect 11060 10183 11112 10192
rect 11060 10149 11069 10183
rect 11069 10149 11103 10183
rect 11103 10149 11112 10183
rect 11060 10140 11112 10149
rect 12440 10115 12492 10124
rect 8944 10004 8996 10056
rect 10324 10004 10376 10056
rect 5816 9868 5868 9920
rect 6000 9868 6052 9920
rect 6920 9936 6972 9988
rect 8300 9936 8352 9988
rect 9680 9936 9732 9988
rect 10140 9936 10192 9988
rect 10784 10004 10836 10056
rect 12440 10081 12449 10115
rect 12449 10081 12483 10115
rect 12483 10081 12492 10115
rect 12440 10072 12492 10081
rect 12900 10072 12952 10124
rect 13360 10072 13412 10124
rect 16304 10072 16356 10124
rect 15568 10047 15620 10056
rect 15568 10013 15577 10047
rect 15577 10013 15611 10047
rect 15611 10013 15620 10047
rect 15568 10004 15620 10013
rect 15936 9979 15988 9988
rect 15936 9945 15945 9979
rect 15945 9945 15979 9979
rect 15979 9945 15988 9979
rect 15936 9936 15988 9945
rect 6736 9868 6788 9920
rect 7104 9868 7156 9920
rect 8116 9868 8168 9920
rect 9772 9868 9824 9920
rect 10048 9911 10100 9920
rect 10048 9877 10057 9911
rect 10057 9877 10091 9911
rect 10091 9877 10100 9911
rect 10048 9868 10100 9877
rect 11336 9868 11388 9920
rect 12624 9911 12676 9920
rect 12624 9877 12633 9911
rect 12633 9877 12667 9911
rect 12667 9877 12676 9911
rect 12624 9868 12676 9877
rect 13084 9911 13136 9920
rect 13084 9877 13093 9911
rect 13093 9877 13127 9911
rect 13127 9877 13136 9911
rect 13084 9868 13136 9877
rect 3680 9766 3732 9818
rect 3744 9766 3796 9818
rect 3808 9766 3860 9818
rect 3872 9766 3924 9818
rect 9078 9766 9130 9818
rect 9142 9766 9194 9818
rect 9206 9766 9258 9818
rect 9270 9766 9322 9818
rect 14475 9766 14527 9818
rect 14539 9766 14591 9818
rect 14603 9766 14655 9818
rect 14667 9766 14719 9818
rect 4068 9664 4120 9716
rect 6736 9664 6788 9716
rect 10048 9664 10100 9716
rect 15568 9664 15620 9716
rect 15936 9664 15988 9716
rect 2596 9639 2648 9648
rect 2596 9605 2605 9639
rect 2605 9605 2639 9639
rect 2639 9605 2648 9639
rect 2596 9596 2648 9605
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 2412 9528 2464 9580
rect 12256 9596 12308 9648
rect 3516 9528 3568 9580
rect 2688 9460 2740 9512
rect 3240 9460 3292 9512
rect 3976 9528 4028 9580
rect 4804 9503 4856 9512
rect 1400 9367 1452 9376
rect 1400 9333 1409 9367
rect 1409 9333 1443 9367
rect 1443 9333 1452 9367
rect 1400 9324 1452 9333
rect 1860 9367 1912 9376
rect 1860 9333 1869 9367
rect 1869 9333 1903 9367
rect 1903 9333 1912 9367
rect 1860 9324 1912 9333
rect 2228 9392 2280 9444
rect 4804 9469 4813 9503
rect 4813 9469 4847 9503
rect 4847 9469 4856 9503
rect 4804 9460 4856 9469
rect 4988 9503 5040 9512
rect 4988 9469 4997 9503
rect 4997 9469 5031 9503
rect 5031 9469 5040 9503
rect 4988 9460 5040 9469
rect 7472 9528 7524 9580
rect 7748 9528 7800 9580
rect 7932 9460 7984 9512
rect 8116 9503 8168 9512
rect 8116 9469 8125 9503
rect 8125 9469 8159 9503
rect 8159 9469 8168 9503
rect 8116 9460 8168 9469
rect 8208 9503 8260 9512
rect 8208 9469 8217 9503
rect 8217 9469 8251 9503
rect 8251 9469 8260 9503
rect 9680 9528 9732 9580
rect 10140 9528 10192 9580
rect 10232 9528 10284 9580
rect 11060 9528 11112 9580
rect 12716 9571 12768 9580
rect 12716 9537 12725 9571
rect 12725 9537 12759 9571
rect 12759 9537 12768 9571
rect 12716 9528 12768 9537
rect 13084 9528 13136 9580
rect 8208 9460 8260 9469
rect 9588 9503 9640 9512
rect 5632 9392 5684 9444
rect 7012 9435 7064 9444
rect 7012 9401 7021 9435
rect 7021 9401 7055 9435
rect 7055 9401 7064 9435
rect 7012 9392 7064 9401
rect 7196 9435 7248 9444
rect 7196 9401 7205 9435
rect 7205 9401 7239 9435
rect 7239 9401 7248 9435
rect 7196 9392 7248 9401
rect 8024 9392 8076 9444
rect 9588 9469 9597 9503
rect 9597 9469 9631 9503
rect 9631 9469 9640 9503
rect 9588 9460 9640 9469
rect 9772 9460 9824 9512
rect 10784 9503 10836 9512
rect 10784 9469 10793 9503
rect 10793 9469 10827 9503
rect 10827 9469 10836 9503
rect 10784 9460 10836 9469
rect 10876 9460 10928 9512
rect 12624 9460 12676 9512
rect 13268 9460 13320 9512
rect 14740 9460 14792 9512
rect 15936 9460 15988 9512
rect 9496 9392 9548 9444
rect 3608 9324 3660 9376
rect 8576 9367 8628 9376
rect 8576 9333 8585 9367
rect 8585 9333 8619 9367
rect 8619 9333 8628 9367
rect 8576 9324 8628 9333
rect 9036 9324 9088 9376
rect 10324 9324 10376 9376
rect 11152 9367 11204 9376
rect 11152 9333 11161 9367
rect 11161 9333 11195 9367
rect 11195 9333 11204 9367
rect 11152 9324 11204 9333
rect 11612 9324 11664 9376
rect 13360 9367 13412 9376
rect 13360 9333 13369 9367
rect 13369 9333 13403 9367
rect 13403 9333 13412 9367
rect 13360 9324 13412 9333
rect 13728 9324 13780 9376
rect 15200 9367 15252 9376
rect 15200 9333 15209 9367
rect 15209 9333 15243 9367
rect 15243 9333 15252 9367
rect 15200 9324 15252 9333
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 6571 9222 6623 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 11904 9222 11956 9274
rect 11968 9222 12020 9274
rect 2228 9163 2280 9172
rect 2228 9129 2237 9163
rect 2237 9129 2271 9163
rect 2271 9129 2280 9163
rect 2228 9120 2280 9129
rect 3608 9120 3660 9172
rect 5816 9120 5868 9172
rect 7104 9120 7156 9172
rect 9496 9120 9548 9172
rect 12348 9163 12400 9172
rect 12348 9129 12357 9163
rect 12357 9129 12391 9163
rect 12391 9129 12400 9163
rect 12348 9120 12400 9129
rect 13268 9120 13320 9172
rect 14740 9163 14792 9172
rect 14740 9129 14749 9163
rect 14749 9129 14783 9163
rect 14783 9129 14792 9163
rect 14740 9120 14792 9129
rect 1860 9052 1912 9104
rect 5816 8984 5868 9036
rect 1400 8916 1452 8968
rect 2780 8959 2832 8968
rect 2780 8925 2789 8959
rect 2789 8925 2823 8959
rect 2823 8925 2832 8959
rect 3148 8959 3200 8968
rect 2780 8916 2832 8925
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 5080 8959 5132 8968
rect 5080 8925 5089 8959
rect 5089 8925 5123 8959
rect 5123 8925 5132 8959
rect 5080 8916 5132 8925
rect 5356 8916 5408 8968
rect 2504 8848 2556 8900
rect 6368 8984 6420 9036
rect 6736 9027 6788 9036
rect 6736 8993 6745 9027
rect 6745 8993 6779 9027
rect 6779 8993 6788 9027
rect 6736 8984 6788 8993
rect 6920 9027 6972 9036
rect 6920 8993 6929 9027
rect 6929 8993 6963 9027
rect 6963 8993 6972 9027
rect 6920 8984 6972 8993
rect 7104 8984 7156 9036
rect 8300 8984 8352 9036
rect 9404 8984 9456 9036
rect 9680 8984 9732 9036
rect 9956 9027 10008 9036
rect 9956 8993 9965 9027
rect 9965 8993 9999 9027
rect 9999 8993 10008 9027
rect 9956 8984 10008 8993
rect 7932 8916 7984 8968
rect 8024 8916 8076 8968
rect 6552 8891 6604 8900
rect 2596 8780 2648 8832
rect 4620 8823 4672 8832
rect 4620 8789 4629 8823
rect 4629 8789 4663 8823
rect 4663 8789 4672 8823
rect 4620 8780 4672 8789
rect 5448 8780 5500 8832
rect 6000 8823 6052 8832
rect 6000 8789 6009 8823
rect 6009 8789 6043 8823
rect 6043 8789 6052 8823
rect 6000 8780 6052 8789
rect 6552 8857 6561 8891
rect 6561 8857 6595 8891
rect 6595 8857 6604 8891
rect 6552 8848 6604 8857
rect 6736 8780 6788 8832
rect 7472 8823 7524 8832
rect 7472 8789 7481 8823
rect 7481 8789 7515 8823
rect 7515 8789 7524 8823
rect 7472 8780 7524 8789
rect 8024 8780 8076 8832
rect 8484 8916 8536 8968
rect 13544 9052 13596 9104
rect 13728 9095 13780 9104
rect 13728 9061 13737 9095
rect 13737 9061 13771 9095
rect 13771 9061 13780 9095
rect 13728 9052 13780 9061
rect 15844 9052 15896 9104
rect 12256 9027 12308 9036
rect 12256 8993 12265 9027
rect 12265 8993 12299 9027
rect 12299 8993 12308 9027
rect 12256 8984 12308 8993
rect 13268 9027 13320 9036
rect 13268 8993 13277 9027
rect 13277 8993 13311 9027
rect 13311 8993 13320 9027
rect 13268 8984 13320 8993
rect 15016 8984 15068 9036
rect 15568 8984 15620 9036
rect 11336 8959 11388 8968
rect 8668 8848 8720 8900
rect 9864 8891 9916 8900
rect 9864 8857 9873 8891
rect 9873 8857 9907 8891
rect 9907 8857 9916 8891
rect 9864 8848 9916 8857
rect 9772 8780 9824 8832
rect 10784 8848 10836 8900
rect 11336 8925 11345 8959
rect 11345 8925 11379 8959
rect 11379 8925 11388 8959
rect 11336 8916 11388 8925
rect 12716 8916 12768 8968
rect 12992 8916 13044 8968
rect 15936 8916 15988 8968
rect 14372 8848 14424 8900
rect 3680 8678 3732 8730
rect 3744 8678 3796 8730
rect 3808 8678 3860 8730
rect 3872 8678 3924 8730
rect 9078 8678 9130 8730
rect 9142 8678 9194 8730
rect 9206 8678 9258 8730
rect 9270 8678 9322 8730
rect 14475 8678 14527 8730
rect 14539 8678 14591 8730
rect 14603 8678 14655 8730
rect 14667 8678 14719 8730
rect 2596 8619 2648 8628
rect 2596 8585 2605 8619
rect 2605 8585 2639 8619
rect 2639 8585 2648 8619
rect 2596 8576 2648 8585
rect 5080 8576 5132 8628
rect 5816 8576 5868 8628
rect 7840 8576 7892 8628
rect 8024 8576 8076 8628
rect 4436 8440 4488 8492
rect 2688 8372 2740 8424
rect 3148 8415 3200 8424
rect 3148 8381 3157 8415
rect 3157 8381 3191 8415
rect 3191 8381 3200 8415
rect 3148 8372 3200 8381
rect 8300 8508 8352 8560
rect 9588 8508 9640 8560
rect 10508 8576 10560 8628
rect 13544 8576 13596 8628
rect 4988 8440 5040 8492
rect 5356 8440 5408 8492
rect 5632 8483 5684 8492
rect 5632 8449 5641 8483
rect 5641 8449 5675 8483
rect 5675 8449 5684 8483
rect 5632 8440 5684 8449
rect 5908 8440 5960 8492
rect 6552 8440 6604 8492
rect 7104 8440 7156 8492
rect 8116 8440 8168 8492
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 5540 8372 5592 8381
rect 6000 8372 6052 8424
rect 7012 8372 7064 8424
rect 7288 8372 7340 8424
rect 7472 8415 7524 8424
rect 7472 8381 7481 8415
rect 7481 8381 7515 8415
rect 7515 8381 7524 8415
rect 7472 8372 7524 8381
rect 7748 8415 7800 8424
rect 1400 8347 1452 8356
rect 1400 8313 1409 8347
rect 1409 8313 1443 8347
rect 1443 8313 1452 8347
rect 1400 8304 1452 8313
rect 2136 8304 2188 8356
rect 6368 8304 6420 8356
rect 6920 8304 6972 8356
rect 7748 8381 7757 8415
rect 7757 8381 7791 8415
rect 7791 8381 7800 8415
rect 7748 8372 7800 8381
rect 7840 8372 7892 8424
rect 9404 8440 9456 8492
rect 9772 8440 9824 8492
rect 8760 8415 8812 8424
rect 8760 8381 8769 8415
rect 8769 8381 8803 8415
rect 8803 8381 8812 8415
rect 8760 8372 8812 8381
rect 9680 8372 9732 8424
rect 11244 8508 11296 8560
rect 11428 8508 11480 8560
rect 10324 8483 10376 8492
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 12992 8483 13044 8492
rect 10324 8440 10376 8449
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 14280 8440 14332 8492
rect 8208 8304 8260 8356
rect 4252 8236 4304 8288
rect 6000 8236 6052 8288
rect 7932 8279 7984 8288
rect 7932 8245 7941 8279
rect 7941 8245 7975 8279
rect 7975 8245 7984 8279
rect 7932 8236 7984 8245
rect 8024 8236 8076 8288
rect 9864 8304 9916 8356
rect 10048 8304 10100 8356
rect 10232 8236 10284 8288
rect 13728 8372 13780 8424
rect 14832 8415 14884 8424
rect 14832 8381 14841 8415
rect 14841 8381 14875 8415
rect 14875 8381 14884 8415
rect 14832 8372 14884 8381
rect 15292 8415 15344 8424
rect 15292 8381 15301 8415
rect 15301 8381 15335 8415
rect 15335 8381 15344 8415
rect 15292 8372 15344 8381
rect 13912 8347 13964 8356
rect 12808 8279 12860 8288
rect 12808 8245 12817 8279
rect 12817 8245 12851 8279
rect 12851 8245 12860 8279
rect 12808 8236 12860 8245
rect 13912 8313 13921 8347
rect 13921 8313 13955 8347
rect 13955 8313 13964 8347
rect 13912 8304 13964 8313
rect 15844 8304 15896 8356
rect 15108 8236 15160 8288
rect 15660 8279 15712 8288
rect 15660 8245 15669 8279
rect 15669 8245 15703 8279
rect 15703 8245 15712 8279
rect 15660 8236 15712 8245
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 6571 8134 6623 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 11904 8134 11956 8186
rect 11968 8134 12020 8186
rect 2596 8032 2648 8084
rect 2780 8032 2832 8084
rect 5724 8032 5776 8084
rect 7196 8032 7248 8084
rect 2228 7964 2280 8016
rect 2504 8007 2556 8016
rect 2504 7973 2513 8007
rect 2513 7973 2547 8007
rect 2547 7973 2556 8007
rect 2504 7964 2556 7973
rect 6184 7964 6236 8016
rect 1492 7896 1544 7948
rect 2688 7896 2740 7948
rect 4160 7896 4212 7948
rect 5540 7896 5592 7948
rect 5816 7896 5868 7948
rect 7104 7939 7156 7948
rect 7104 7905 7113 7939
rect 7113 7905 7147 7939
rect 7147 7905 7156 7939
rect 7104 7896 7156 7905
rect 7380 7964 7432 8016
rect 8668 7964 8720 8016
rect 12348 8032 12400 8084
rect 12808 8032 12860 8084
rect 14372 8032 14424 8084
rect 15200 8032 15252 8084
rect 5356 7828 5408 7880
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 1952 7760 2004 7812
rect 2228 7760 2280 7812
rect 7472 7828 7524 7880
rect 10232 7896 10284 7948
rect 11152 7939 11204 7948
rect 7932 7828 7984 7880
rect 11152 7905 11161 7939
rect 11161 7905 11195 7939
rect 11195 7905 11204 7939
rect 11152 7896 11204 7905
rect 11336 7896 11388 7948
rect 11520 7896 11572 7948
rect 10416 7828 10468 7880
rect 12716 7896 12768 7948
rect 13176 7939 13228 7948
rect 13176 7905 13185 7939
rect 13185 7905 13219 7939
rect 13219 7905 13228 7939
rect 13176 7896 13228 7905
rect 14924 7896 14976 7948
rect 15660 7964 15712 8016
rect 15292 7939 15344 7948
rect 15292 7905 15323 7939
rect 15323 7905 15344 7939
rect 15292 7896 15344 7905
rect 15844 7939 15896 7948
rect 15844 7905 15853 7939
rect 15853 7905 15887 7939
rect 15887 7905 15896 7939
rect 15844 7896 15896 7905
rect 17040 7896 17092 7948
rect 15016 7828 15068 7880
rect 4344 7735 4396 7744
rect 4344 7701 4353 7735
rect 4353 7701 4387 7735
rect 4387 7701 4396 7735
rect 4344 7692 4396 7701
rect 6736 7692 6788 7744
rect 6920 7735 6972 7744
rect 6920 7701 6929 7735
rect 6929 7701 6963 7735
rect 6963 7701 6972 7735
rect 6920 7692 6972 7701
rect 7748 7735 7800 7744
rect 7748 7701 7757 7735
rect 7757 7701 7791 7735
rect 7791 7701 7800 7735
rect 7748 7692 7800 7701
rect 9588 7692 9640 7744
rect 9864 7760 9916 7812
rect 9956 7692 10008 7744
rect 10048 7692 10100 7744
rect 13728 7735 13780 7744
rect 13728 7701 13737 7735
rect 13737 7701 13771 7735
rect 13771 7701 13780 7735
rect 13728 7692 13780 7701
rect 3680 7590 3732 7642
rect 3744 7590 3796 7642
rect 3808 7590 3860 7642
rect 3872 7590 3924 7642
rect 9078 7590 9130 7642
rect 9142 7590 9194 7642
rect 9206 7590 9258 7642
rect 9270 7590 9322 7642
rect 14475 7590 14527 7642
rect 14539 7590 14591 7642
rect 14603 7590 14655 7642
rect 14667 7590 14719 7642
rect 2688 7488 2740 7540
rect 5908 7488 5960 7540
rect 8668 7488 8720 7540
rect 9588 7488 9640 7540
rect 10140 7488 10192 7540
rect 12256 7488 12308 7540
rect 13176 7488 13228 7540
rect 15108 7488 15160 7540
rect 4252 7420 4304 7472
rect 7196 7420 7248 7472
rect 2872 7284 2924 7336
rect 3056 7284 3108 7336
rect 5540 7352 5592 7404
rect 10048 7420 10100 7472
rect 12164 7463 12216 7472
rect 12164 7429 12173 7463
rect 12173 7429 12207 7463
rect 12207 7429 12216 7463
rect 12164 7420 12216 7429
rect 15016 7463 15068 7472
rect 15016 7429 15025 7463
rect 15025 7429 15059 7463
rect 15059 7429 15068 7463
rect 15016 7420 15068 7429
rect 7748 7352 7800 7404
rect 4712 7284 4764 7336
rect 5632 7284 5684 7336
rect 5908 7284 5960 7336
rect 7380 7284 7432 7336
rect 8300 7327 8352 7336
rect 8300 7293 8309 7327
rect 8309 7293 8343 7327
rect 8343 7293 8352 7327
rect 8300 7284 8352 7293
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 8944 7284 8996 7336
rect 2688 7216 2740 7268
rect 3332 7216 3384 7268
rect 4160 7259 4212 7268
rect 4160 7225 4169 7259
rect 4169 7225 4203 7259
rect 4203 7225 4212 7259
rect 4160 7216 4212 7225
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 2504 7148 2556 7200
rect 5724 7216 5776 7268
rect 9680 7216 9732 7268
rect 8208 7148 8260 7200
rect 8576 7148 8628 7200
rect 9864 7259 9916 7268
rect 9864 7225 9873 7259
rect 9873 7225 9907 7259
rect 9907 7225 9916 7259
rect 10048 7259 10100 7268
rect 9864 7216 9916 7225
rect 10048 7225 10057 7259
rect 10057 7225 10091 7259
rect 10091 7225 10100 7259
rect 10048 7216 10100 7225
rect 10968 7284 11020 7336
rect 12992 7352 13044 7404
rect 15660 7284 15712 7336
rect 16396 7327 16448 7336
rect 16396 7293 16405 7327
rect 16405 7293 16439 7327
rect 16439 7293 16448 7327
rect 16396 7284 16448 7293
rect 12532 7216 12584 7268
rect 12808 7216 12860 7268
rect 10324 7148 10376 7200
rect 11060 7191 11112 7200
rect 11060 7157 11069 7191
rect 11069 7157 11103 7191
rect 11103 7157 11112 7191
rect 11060 7148 11112 7157
rect 14924 7216 14976 7268
rect 13636 7191 13688 7200
rect 13636 7157 13645 7191
rect 13645 7157 13679 7191
rect 13679 7157 13688 7191
rect 13636 7148 13688 7157
rect 14188 7148 14240 7200
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 6571 7046 6623 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 11904 7046 11956 7098
rect 11968 7046 12020 7098
rect 1584 6944 1636 6996
rect 5448 6944 5500 6996
rect 8208 6987 8260 6996
rect 8208 6953 8217 6987
rect 8217 6953 8251 6987
rect 8251 6953 8260 6987
rect 8208 6944 8260 6953
rect 8300 6944 8352 6996
rect 8944 6944 8996 6996
rect 10324 6944 10376 6996
rect 12808 6944 12860 6996
rect 13636 6944 13688 6996
rect 13728 6944 13780 6996
rect 15844 6944 15896 6996
rect 3056 6808 3108 6860
rect 4620 6808 4672 6860
rect 5908 6851 5960 6860
rect 2504 6740 2556 6792
rect 4068 6740 4120 6792
rect 4252 6783 4304 6792
rect 4252 6749 4261 6783
rect 4261 6749 4295 6783
rect 4295 6749 4304 6783
rect 4252 6740 4304 6749
rect 5908 6817 5917 6851
rect 5917 6817 5951 6851
rect 5951 6817 5960 6851
rect 5908 6808 5960 6817
rect 6000 6851 6052 6860
rect 6000 6817 6009 6851
rect 6009 6817 6043 6851
rect 6043 6817 6052 6851
rect 6000 6808 6052 6817
rect 6920 6876 6972 6928
rect 8484 6876 8536 6928
rect 7564 6808 7616 6860
rect 9680 6851 9732 6860
rect 9680 6817 9689 6851
rect 9689 6817 9723 6851
rect 9723 6817 9732 6851
rect 9680 6808 9732 6817
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 1952 6672 2004 6724
rect 4344 6715 4396 6724
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 3332 6647 3384 6656
rect 3332 6613 3341 6647
rect 3341 6613 3375 6647
rect 3375 6613 3384 6647
rect 3332 6604 3384 6613
rect 4344 6681 4353 6715
rect 4353 6681 4387 6715
rect 4387 6681 4396 6715
rect 4344 6672 4396 6681
rect 4712 6672 4764 6724
rect 7012 6672 7064 6724
rect 8208 6740 8260 6792
rect 10876 6808 10928 6860
rect 10968 6808 11020 6860
rect 10600 6740 10652 6792
rect 12164 6876 12216 6928
rect 12716 6919 12768 6928
rect 12716 6885 12725 6919
rect 12725 6885 12759 6919
rect 12759 6885 12768 6919
rect 12716 6876 12768 6885
rect 8484 6672 8536 6724
rect 7288 6604 7340 6656
rect 8576 6647 8628 6656
rect 8576 6613 8585 6647
rect 8585 6613 8619 6647
rect 8619 6613 8628 6647
rect 8576 6604 8628 6613
rect 8852 6604 8904 6656
rect 10140 6604 10192 6656
rect 13176 6808 13228 6860
rect 13912 6808 13964 6860
rect 14832 6851 14884 6860
rect 14832 6817 14841 6851
rect 14841 6817 14875 6851
rect 14875 6817 14884 6851
rect 14832 6808 14884 6817
rect 15200 6808 15252 6860
rect 16212 6808 16264 6860
rect 15384 6672 15436 6724
rect 15292 6604 15344 6656
rect 3680 6502 3732 6554
rect 3744 6502 3796 6554
rect 3808 6502 3860 6554
rect 3872 6502 3924 6554
rect 9078 6502 9130 6554
rect 9142 6502 9194 6554
rect 9206 6502 9258 6554
rect 9270 6502 9322 6554
rect 14475 6502 14527 6554
rect 14539 6502 14591 6554
rect 14603 6502 14655 6554
rect 14667 6502 14719 6554
rect 4068 6400 4120 6452
rect 5448 6443 5500 6452
rect 5448 6409 5457 6443
rect 5457 6409 5491 6443
rect 5491 6409 5500 6443
rect 5448 6400 5500 6409
rect 4896 6332 4948 6384
rect 8208 6400 8260 6452
rect 8392 6443 8444 6452
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 8668 6400 8720 6452
rect 10416 6400 10468 6452
rect 10968 6400 11020 6452
rect 14188 6443 14240 6452
rect 14188 6409 14197 6443
rect 14197 6409 14231 6443
rect 14231 6409 14240 6443
rect 14188 6400 14240 6409
rect 16212 6443 16264 6452
rect 16212 6409 16221 6443
rect 16221 6409 16255 6443
rect 16255 6409 16264 6443
rect 16212 6400 16264 6409
rect 2504 6264 2556 6316
rect 1952 6239 2004 6248
rect 1952 6205 1961 6239
rect 1961 6205 1995 6239
rect 1995 6205 2004 6239
rect 1952 6196 2004 6205
rect 2688 6196 2740 6248
rect 4344 6264 4396 6316
rect 7380 6332 7432 6384
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 8024 6264 8076 6316
rect 4528 6196 4580 6248
rect 1952 6060 2004 6112
rect 4712 6196 4764 6248
rect 5632 6239 5684 6248
rect 5632 6205 5641 6239
rect 5641 6205 5675 6239
rect 5675 6205 5684 6239
rect 5632 6196 5684 6205
rect 6000 6196 6052 6248
rect 7748 6196 7800 6248
rect 10140 6332 10192 6384
rect 11060 6332 11112 6384
rect 12256 6332 12308 6384
rect 8576 6264 8628 6316
rect 8484 6239 8536 6248
rect 8484 6205 8493 6239
rect 8493 6205 8527 6239
rect 8527 6205 8536 6239
rect 8484 6196 8536 6205
rect 7380 6128 7432 6180
rect 9036 6196 9088 6248
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 10600 6196 10652 6248
rect 13728 6196 13780 6248
rect 14372 6239 14424 6248
rect 14372 6205 14381 6239
rect 14381 6205 14415 6239
rect 14415 6205 14424 6239
rect 14372 6196 14424 6205
rect 15384 6239 15436 6248
rect 15384 6205 15393 6239
rect 15393 6205 15427 6239
rect 15427 6205 15436 6239
rect 15384 6196 15436 6205
rect 16212 6239 16264 6248
rect 16212 6205 16221 6239
rect 16221 6205 16255 6239
rect 16255 6205 16264 6239
rect 16212 6196 16264 6205
rect 4252 6060 4304 6112
rect 6828 6103 6880 6112
rect 6828 6069 6837 6103
rect 6837 6069 6871 6103
rect 6871 6069 6880 6103
rect 6828 6060 6880 6069
rect 7288 6060 7340 6112
rect 8116 6103 8168 6112
rect 8116 6069 8125 6103
rect 8125 6069 8159 6103
rect 8159 6069 8168 6103
rect 8116 6060 8168 6069
rect 8484 6060 8536 6112
rect 10232 6128 10284 6180
rect 9864 6060 9916 6112
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 6571 5958 6623 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 11904 5958 11956 6010
rect 11968 5958 12020 6010
rect 2320 5856 2372 5908
rect 4804 5856 4856 5908
rect 6920 5856 6972 5908
rect 1584 5720 1636 5772
rect 2872 5720 2924 5772
rect 4620 5763 4672 5772
rect 4620 5729 4629 5763
rect 4629 5729 4663 5763
rect 4663 5729 4672 5763
rect 4620 5720 4672 5729
rect 4896 5788 4948 5840
rect 7656 5856 7708 5908
rect 11612 5856 11664 5908
rect 12532 5856 12584 5908
rect 5632 5720 5684 5772
rect 8208 5763 8260 5772
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 5724 5652 5776 5704
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 7748 5695 7800 5704
rect 7748 5661 7757 5695
rect 7757 5661 7791 5695
rect 7791 5661 7800 5695
rect 7748 5652 7800 5661
rect 8208 5729 8217 5763
rect 8217 5729 8251 5763
rect 8251 5729 8260 5763
rect 8208 5720 8260 5729
rect 10968 5720 11020 5772
rect 8484 5652 8536 5704
rect 10508 5695 10560 5704
rect 2780 5584 2832 5636
rect 7012 5584 7064 5636
rect 7564 5584 7616 5636
rect 10508 5661 10517 5695
rect 10517 5661 10551 5695
rect 10551 5661 10560 5695
rect 10508 5652 10560 5661
rect 12256 5788 12308 5840
rect 13360 5788 13412 5840
rect 11152 5763 11204 5772
rect 11152 5729 11161 5763
rect 11161 5729 11195 5763
rect 11195 5729 11204 5763
rect 11612 5763 11664 5772
rect 11152 5720 11204 5729
rect 11612 5729 11621 5763
rect 11621 5729 11655 5763
rect 11655 5729 11664 5763
rect 11612 5720 11664 5729
rect 12072 5720 12124 5772
rect 13820 5763 13872 5772
rect 13820 5729 13829 5763
rect 13829 5729 13863 5763
rect 13863 5729 13872 5763
rect 13820 5720 13872 5729
rect 15568 5788 15620 5840
rect 15384 5720 15436 5772
rect 15936 5652 15988 5704
rect 5908 5559 5960 5568
rect 5908 5525 5917 5559
rect 5917 5525 5951 5559
rect 5951 5525 5960 5559
rect 5908 5516 5960 5525
rect 7288 5559 7340 5568
rect 7288 5525 7297 5559
rect 7297 5525 7331 5559
rect 7331 5525 7340 5559
rect 7288 5516 7340 5525
rect 8392 5516 8444 5568
rect 9956 5516 10008 5568
rect 10140 5559 10192 5568
rect 10140 5525 10149 5559
rect 10149 5525 10183 5559
rect 10183 5525 10192 5559
rect 10140 5516 10192 5525
rect 12164 5559 12216 5568
rect 12164 5525 12173 5559
rect 12173 5525 12207 5559
rect 12207 5525 12216 5559
rect 12164 5516 12216 5525
rect 14372 5559 14424 5568
rect 14372 5525 14381 5559
rect 14381 5525 14415 5559
rect 14415 5525 14424 5559
rect 14372 5516 14424 5525
rect 14832 5516 14884 5568
rect 15476 5516 15528 5568
rect 3680 5414 3732 5466
rect 3744 5414 3796 5466
rect 3808 5414 3860 5466
rect 3872 5414 3924 5466
rect 9078 5414 9130 5466
rect 9142 5414 9194 5466
rect 9206 5414 9258 5466
rect 9270 5414 9322 5466
rect 14475 5414 14527 5466
rect 14539 5414 14591 5466
rect 14603 5414 14655 5466
rect 14667 5414 14719 5466
rect 2320 5355 2372 5364
rect 2320 5321 2329 5355
rect 2329 5321 2363 5355
rect 2363 5321 2372 5355
rect 2320 5312 2372 5321
rect 2780 5355 2832 5364
rect 2780 5321 2789 5355
rect 2789 5321 2823 5355
rect 2823 5321 2832 5355
rect 2780 5312 2832 5321
rect 7196 5312 7248 5364
rect 8208 5312 8260 5364
rect 10140 5312 10192 5364
rect 14372 5312 14424 5364
rect 11612 5244 11664 5296
rect 4804 5176 4856 5228
rect 6460 5176 6512 5228
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 8944 5176 8996 5228
rect 13084 5176 13136 5228
rect 15476 5219 15528 5228
rect 15476 5185 15485 5219
rect 15485 5185 15519 5219
rect 15519 5185 15528 5219
rect 15476 5176 15528 5185
rect 1584 5108 1636 5160
rect 2412 5108 2464 5160
rect 5264 5151 5316 5160
rect 5264 5117 5273 5151
rect 5273 5117 5307 5151
rect 5307 5117 5316 5151
rect 5264 5108 5316 5117
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 7380 5151 7432 5160
rect 7380 5117 7389 5151
rect 7389 5117 7423 5151
rect 7423 5117 7432 5151
rect 7380 5108 7432 5117
rect 8116 5108 8168 5160
rect 9772 5108 9824 5160
rect 5080 5083 5132 5092
rect 5080 5049 5089 5083
rect 5089 5049 5123 5083
rect 5123 5049 5132 5083
rect 5080 5040 5132 5049
rect 8024 5040 8076 5092
rect 10508 5108 10560 5160
rect 11244 5108 11296 5160
rect 12072 5108 12124 5160
rect 13360 5108 13412 5160
rect 14280 5108 14332 5160
rect 11152 5040 11204 5092
rect 14188 5083 14240 5092
rect 14188 5049 14197 5083
rect 14197 5049 14231 5083
rect 14231 5049 14240 5083
rect 14188 5040 14240 5049
rect 4160 4972 4212 5024
rect 7748 4972 7800 5024
rect 8576 5015 8628 5024
rect 8576 4981 8585 5015
rect 8585 4981 8619 5015
rect 8619 4981 8628 5015
rect 8576 4972 8628 4981
rect 8668 4972 8720 5024
rect 12072 5015 12124 5024
rect 12072 4981 12081 5015
rect 12081 4981 12115 5015
rect 12115 4981 12124 5015
rect 12072 4972 12124 4981
rect 14004 4972 14056 5024
rect 15384 5108 15436 5160
rect 15936 5108 15988 5160
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 6571 4870 6623 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 11904 4870 11956 4922
rect 11968 4870 12020 4922
rect 3516 4768 3568 4820
rect 9404 4811 9456 4820
rect 1952 4632 2004 4684
rect 2412 4632 2464 4684
rect 7380 4700 7432 4752
rect 9404 4777 9413 4811
rect 9413 4777 9447 4811
rect 9447 4777 9456 4811
rect 9404 4768 9456 4777
rect 10140 4768 10192 4820
rect 10784 4768 10836 4820
rect 11244 4743 11296 4752
rect 5540 4675 5592 4684
rect 2780 4607 2832 4616
rect 2780 4573 2789 4607
rect 2789 4573 2823 4607
rect 2823 4573 2832 4607
rect 5540 4641 5549 4675
rect 5549 4641 5583 4675
rect 5583 4641 5592 4675
rect 5540 4632 5592 4641
rect 5908 4632 5960 4684
rect 7472 4632 7524 4684
rect 8024 4675 8076 4684
rect 8024 4641 8033 4675
rect 8033 4641 8067 4675
rect 8067 4641 8076 4675
rect 8024 4632 8076 4641
rect 8576 4675 8628 4684
rect 8576 4641 8585 4675
rect 8585 4641 8619 4675
rect 8619 4641 8628 4675
rect 8576 4632 8628 4641
rect 11244 4709 11253 4743
rect 11253 4709 11287 4743
rect 11287 4709 11296 4743
rect 11244 4700 11296 4709
rect 12164 4768 12216 4820
rect 15292 4768 15344 4820
rect 15936 4768 15988 4820
rect 16212 4768 16264 4820
rect 2780 4564 2832 4573
rect 5080 4564 5132 4616
rect 11612 4632 11664 4684
rect 12072 4675 12124 4684
rect 12072 4641 12081 4675
rect 12081 4641 12115 4675
rect 12115 4641 12124 4675
rect 12072 4632 12124 4641
rect 12900 4607 12952 4616
rect 12900 4573 12909 4607
rect 12909 4573 12943 4607
rect 12943 4573 12952 4607
rect 12900 4564 12952 4573
rect 13084 4607 13136 4616
rect 13084 4573 13093 4607
rect 13093 4573 13127 4607
rect 13127 4573 13136 4607
rect 13084 4564 13136 4573
rect 14004 4632 14056 4684
rect 15752 4700 15804 4752
rect 13728 4564 13780 4616
rect 15476 4632 15528 4684
rect 14832 4607 14884 4616
rect 14832 4573 14841 4607
rect 14841 4573 14875 4607
rect 14875 4573 14884 4607
rect 14832 4564 14884 4573
rect 3148 4428 3200 4480
rect 7380 4471 7432 4480
rect 7380 4437 7389 4471
rect 7389 4437 7423 4471
rect 7423 4437 7432 4471
rect 7380 4428 7432 4437
rect 8024 4471 8076 4480
rect 8024 4437 8033 4471
rect 8033 4437 8067 4471
rect 8067 4437 8076 4471
rect 8024 4428 8076 4437
rect 10140 4471 10192 4480
rect 10140 4437 10149 4471
rect 10149 4437 10183 4471
rect 10183 4437 10192 4471
rect 10140 4428 10192 4437
rect 3680 4326 3732 4378
rect 3744 4326 3796 4378
rect 3808 4326 3860 4378
rect 3872 4326 3924 4378
rect 9078 4326 9130 4378
rect 9142 4326 9194 4378
rect 9206 4326 9258 4378
rect 9270 4326 9322 4378
rect 14475 4326 14527 4378
rect 14539 4326 14591 4378
rect 14603 4326 14655 4378
rect 14667 4326 14719 4378
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 2780 4088 2832 4140
rect 4436 4088 4488 4140
rect 5540 4088 5592 4140
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 7380 4156 7432 4208
rect 7932 4156 7984 4208
rect 9588 4156 9640 4208
rect 15016 4224 15068 4276
rect 16120 4224 16172 4276
rect 8576 4131 8628 4140
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 10140 4088 10192 4140
rect 11152 4131 11204 4140
rect 11152 4097 11161 4131
rect 11161 4097 11195 4131
rect 11195 4097 11204 4131
rect 11152 4088 11204 4097
rect 12900 4156 12952 4208
rect 2320 4020 2372 4072
rect 4160 4063 4212 4072
rect 4160 4029 4169 4063
rect 4169 4029 4203 4063
rect 4203 4029 4212 4063
rect 4160 4020 4212 4029
rect 4804 4020 4856 4072
rect 5908 4020 5960 4072
rect 8024 4063 8076 4072
rect 8024 4029 8033 4063
rect 8033 4029 8067 4063
rect 8067 4029 8076 4063
rect 8024 4020 8076 4029
rect 9588 4063 9640 4072
rect 9588 4029 9597 4063
rect 9597 4029 9631 4063
rect 9631 4029 9640 4063
rect 9588 4020 9640 4029
rect 10232 4063 10284 4072
rect 10232 4029 10241 4063
rect 10241 4029 10275 4063
rect 10275 4029 10284 4063
rect 10232 4020 10284 4029
rect 10324 4020 10376 4072
rect 13820 4088 13872 4140
rect 15016 4088 15068 4140
rect 3516 3952 3568 4004
rect 1768 3884 1820 3936
rect 8668 3952 8720 4004
rect 8760 3952 8812 4004
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 8024 3884 8076 3936
rect 9036 3884 9088 3936
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 10784 3952 10836 4004
rect 12992 3952 13044 4004
rect 13084 3952 13136 4004
rect 13912 4020 13964 4072
rect 15660 4020 15712 4072
rect 11152 3884 11204 3936
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 13636 3927 13688 3936
rect 12440 3884 12492 3893
rect 13636 3893 13645 3927
rect 13645 3893 13679 3927
rect 13679 3893 13688 3927
rect 13636 3884 13688 3893
rect 16396 3884 16448 3936
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 6571 3782 6623 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 11904 3782 11956 3834
rect 11968 3782 12020 3834
rect 1768 3723 1820 3732
rect 1768 3689 1777 3723
rect 1777 3689 1811 3723
rect 1811 3689 1820 3723
rect 1768 3680 1820 3689
rect 3148 3655 3200 3664
rect 3148 3621 3157 3655
rect 3157 3621 3191 3655
rect 3191 3621 3200 3655
rect 3148 3612 3200 3621
rect 2688 3544 2740 3596
rect 2780 3476 2832 3528
rect 2136 3408 2188 3460
rect 11152 3680 11204 3732
rect 11428 3723 11480 3732
rect 11428 3689 11437 3723
rect 11437 3689 11471 3723
rect 11471 3689 11480 3723
rect 11428 3680 11480 3689
rect 12440 3723 12492 3732
rect 12440 3689 12449 3723
rect 12449 3689 12483 3723
rect 12483 3689 12492 3723
rect 12440 3680 12492 3689
rect 12992 3680 13044 3732
rect 15660 3680 15712 3732
rect 3332 3655 3384 3664
rect 3332 3621 3341 3655
rect 3341 3621 3375 3655
rect 3375 3621 3384 3655
rect 3332 3612 3384 3621
rect 5632 3612 5684 3664
rect 6920 3612 6972 3664
rect 7472 3655 7524 3664
rect 7472 3621 7481 3655
rect 7481 3621 7515 3655
rect 7515 3621 7524 3655
rect 7472 3612 7524 3621
rect 7932 3612 7984 3664
rect 8392 3612 8444 3664
rect 6736 3544 6788 3596
rect 8208 3587 8260 3596
rect 8208 3553 8217 3587
rect 8217 3553 8251 3587
rect 8251 3553 8260 3587
rect 8208 3544 8260 3553
rect 9036 3544 9088 3596
rect 9496 3587 9548 3596
rect 9496 3553 9505 3587
rect 9505 3553 9539 3587
rect 9539 3553 9548 3587
rect 9496 3544 9548 3553
rect 10232 3612 10284 3664
rect 11336 3655 11388 3664
rect 11336 3621 11345 3655
rect 11345 3621 11379 3655
rect 11379 3621 11388 3655
rect 11336 3612 11388 3621
rect 6368 3519 6420 3528
rect 6368 3485 6377 3519
rect 6377 3485 6411 3519
rect 6411 3485 6420 3519
rect 6368 3476 6420 3485
rect 9772 3476 9824 3528
rect 14004 3612 14056 3664
rect 13176 3544 13228 3596
rect 11612 3519 11664 3528
rect 11612 3485 11621 3519
rect 11621 3485 11655 3519
rect 11655 3485 11664 3519
rect 11612 3476 11664 3485
rect 12992 3519 13044 3528
rect 12992 3485 13001 3519
rect 13001 3485 13035 3519
rect 13035 3485 13044 3519
rect 12992 3476 13044 3485
rect 1860 3340 1912 3392
rect 3516 3340 3568 3392
rect 7656 3340 7708 3392
rect 8668 3340 8720 3392
rect 10324 3340 10376 3392
rect 10968 3383 11020 3392
rect 10968 3349 10977 3383
rect 10977 3349 11011 3383
rect 11011 3349 11020 3383
rect 10968 3340 11020 3349
rect 12440 3408 12492 3460
rect 13728 3544 13780 3596
rect 15292 3544 15344 3596
rect 13912 3476 13964 3528
rect 15016 3476 15068 3528
rect 16396 3587 16448 3596
rect 14280 3408 14332 3460
rect 16396 3553 16405 3587
rect 16405 3553 16439 3587
rect 16439 3553 16448 3587
rect 16396 3544 16448 3553
rect 13820 3340 13872 3392
rect 3680 3238 3732 3290
rect 3744 3238 3796 3290
rect 3808 3238 3860 3290
rect 3872 3238 3924 3290
rect 9078 3238 9130 3290
rect 9142 3238 9194 3290
rect 9206 3238 9258 3290
rect 9270 3238 9322 3290
rect 14475 3238 14527 3290
rect 14539 3238 14591 3290
rect 14603 3238 14655 3290
rect 14667 3238 14719 3290
rect 5540 3136 5592 3188
rect 6092 3136 6144 3188
rect 6184 3136 6236 3188
rect 8668 3136 8720 3188
rect 9496 3136 9548 3188
rect 10784 3179 10836 3188
rect 10784 3145 10793 3179
rect 10793 3145 10827 3179
rect 10827 3145 10836 3179
rect 10784 3136 10836 3145
rect 13176 3179 13228 3188
rect 13176 3145 13185 3179
rect 13185 3145 13219 3179
rect 13219 3145 13228 3179
rect 13176 3136 13228 3145
rect 1584 3000 1636 3052
rect 4160 3000 4212 3052
rect 1860 2975 1912 2984
rect 1860 2941 1869 2975
rect 1869 2941 1903 2975
rect 1903 2941 1912 2975
rect 1860 2932 1912 2941
rect 8852 3043 8904 3052
rect 6184 2932 6236 2984
rect 6736 2932 6788 2984
rect 7472 2975 7524 2984
rect 7472 2941 7481 2975
rect 7481 2941 7515 2975
rect 7515 2941 7524 2975
rect 7472 2932 7524 2941
rect 8852 3009 8861 3043
rect 8861 3009 8895 3043
rect 8895 3009 8904 3043
rect 8852 3000 8904 3009
rect 8944 3000 8996 3052
rect 9956 3000 10008 3052
rect 10968 3000 11020 3052
rect 13636 3000 13688 3052
rect 14188 3000 14240 3052
rect 15016 3000 15068 3052
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 5080 2864 5132 2916
rect 2964 2796 3016 2848
rect 5816 2796 5868 2848
rect 7196 2796 7248 2848
rect 9772 2864 9824 2916
rect 9864 2864 9916 2916
rect 10140 2864 10192 2916
rect 13820 2932 13872 2984
rect 15660 2932 15712 2984
rect 7840 2796 7892 2848
rect 8208 2796 8260 2848
rect 12992 2796 13044 2848
rect 13912 2864 13964 2916
rect 13820 2796 13872 2848
rect 15292 2796 15344 2848
rect 16396 2839 16448 2848
rect 16396 2805 16405 2839
rect 16405 2805 16439 2839
rect 16439 2805 16448 2839
rect 16396 2796 16448 2805
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 6571 2694 6623 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 11904 2694 11956 2746
rect 11968 2694 12020 2746
rect 2228 2635 2280 2644
rect 2228 2601 2237 2635
rect 2237 2601 2271 2635
rect 2271 2601 2280 2635
rect 2228 2592 2280 2601
rect 1584 2567 1636 2576
rect 1584 2533 1593 2567
rect 1593 2533 1627 2567
rect 1627 2533 1636 2567
rect 1584 2524 1636 2533
rect 4252 2592 4304 2644
rect 5080 2635 5132 2644
rect 5080 2601 5089 2635
rect 5089 2601 5123 2635
rect 5123 2601 5132 2635
rect 5080 2592 5132 2601
rect 5632 2592 5684 2644
rect 6276 2592 6328 2644
rect 9772 2592 9824 2644
rect 13912 2635 13964 2644
rect 13912 2601 13921 2635
rect 13921 2601 13955 2635
rect 13955 2601 13964 2635
rect 13912 2592 13964 2601
rect 14924 2592 14976 2644
rect 15660 2635 15712 2644
rect 15660 2601 15669 2635
rect 15669 2601 15703 2635
rect 15703 2601 15712 2635
rect 15660 2592 15712 2601
rect 480 2388 532 2440
rect 3056 2456 3108 2508
rect 4804 2456 4856 2508
rect 7932 2524 7984 2576
rect 10784 2524 10836 2576
rect 11612 2524 11664 2576
rect 12808 2524 12860 2576
rect 14832 2524 14884 2576
rect 15108 2524 15160 2576
rect 16396 2567 16448 2576
rect 7840 2499 7892 2508
rect 7840 2465 7849 2499
rect 7849 2465 7883 2499
rect 7883 2465 7892 2499
rect 7840 2456 7892 2465
rect 8300 2456 8352 2508
rect 9496 2456 9548 2508
rect 10048 2456 10100 2508
rect 10140 2456 10192 2508
rect 10968 2499 11020 2508
rect 10968 2465 10977 2499
rect 10977 2465 11011 2499
rect 11011 2465 11020 2499
rect 10968 2456 11020 2465
rect 12440 2456 12492 2508
rect 13820 2499 13872 2508
rect 13820 2465 13829 2499
rect 13829 2465 13863 2499
rect 13863 2465 13872 2499
rect 13820 2456 13872 2465
rect 15752 2456 15804 2508
rect 16396 2533 16405 2567
rect 16405 2533 16439 2567
rect 16439 2533 16448 2567
rect 16396 2524 16448 2533
rect 6920 2388 6972 2440
rect 7196 2388 7248 2440
rect 7656 2388 7708 2440
rect 13084 2388 13136 2440
rect 1400 2363 1452 2372
rect 1400 2329 1409 2363
rect 1409 2329 1443 2363
rect 1443 2329 1452 2363
rect 1400 2320 1452 2329
rect 7748 2320 7800 2372
rect 16580 2363 16632 2372
rect 16580 2329 16589 2363
rect 16589 2329 16623 2363
rect 16623 2329 16632 2363
rect 16580 2320 16632 2329
rect 1308 2252 1360 2304
rect 3680 2150 3732 2202
rect 3744 2150 3796 2202
rect 3808 2150 3860 2202
rect 3872 2150 3924 2202
rect 9078 2150 9130 2202
rect 9142 2150 9194 2202
rect 9206 2150 9258 2202
rect 9270 2150 9322 2202
rect 14475 2150 14527 2202
rect 14539 2150 14591 2202
rect 14603 2150 14655 2202
rect 14667 2150 14719 2202
<< metal2 >>
rect 478 19804 534 20604
rect 1858 19804 1914 20604
rect 3238 19804 3294 20604
rect 4618 19804 4674 20604
rect 5998 19804 6054 20604
rect 7378 19804 7434 20604
rect 8758 19804 8814 20604
rect 10138 19804 10194 20604
rect 11518 19804 11574 20604
rect 12898 19804 12954 20604
rect 14278 19804 14334 20604
rect 15658 19804 15714 20604
rect 17038 19804 17094 20604
rect 492 15978 520 19804
rect 1490 18456 1546 18465
rect 1490 18391 1546 18400
rect 1504 17882 1532 18391
rect 1492 17876 1544 17882
rect 1492 17818 1544 17824
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 1780 17134 1808 17614
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 1676 17060 1728 17066
rect 1676 17002 1728 17008
rect 1688 16726 1716 17002
rect 1676 16720 1728 16726
rect 1676 16662 1728 16668
rect 1400 16584 1452 16590
rect 1400 16526 1452 16532
rect 480 15972 532 15978
rect 480 15914 532 15920
rect 1308 15972 1360 15978
rect 1308 15914 1360 15920
rect 480 2440 532 2446
rect 480 2382 532 2388
rect 492 800 520 2382
rect 1320 2310 1348 15914
rect 1412 14958 1440 16526
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15706 1716 15846
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1780 15570 1808 17070
rect 1872 16046 1900 19804
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1964 16726 1992 16934
rect 1952 16720 2004 16726
rect 1952 16662 2004 16668
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 1768 15564 1820 15570
rect 1768 15506 1820 15512
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1412 12986 1440 14894
rect 1780 14482 1808 15506
rect 2136 15360 2188 15366
rect 2136 15302 2188 15308
rect 2228 15360 2280 15366
rect 2228 15302 2280 15308
rect 2148 14890 2176 15302
rect 2240 15026 2268 15302
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 2136 14884 2188 14890
rect 2136 14826 2188 14832
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1780 13394 1808 14418
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1400 12980 1452 12986
rect 1400 12922 1452 12928
rect 1964 12434 1992 14350
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2240 12714 2268 13126
rect 2228 12708 2280 12714
rect 2228 12650 2280 12656
rect 1872 12406 1992 12434
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1490 10296 1546 10305
rect 1780 10266 1808 10406
rect 1490 10231 1492 10240
rect 1544 10231 1546 10240
rect 1768 10260 1820 10266
rect 1492 10202 1544 10208
rect 1768 10202 1820 10208
rect 1872 9466 1900 12406
rect 2332 12374 2360 18022
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 2872 17060 2924 17066
rect 2872 17002 2924 17008
rect 2884 16250 2912 17002
rect 2976 16726 3004 17206
rect 3056 17128 3108 17134
rect 3056 17070 3108 17076
rect 2964 16720 3016 16726
rect 2964 16662 3016 16668
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2872 15564 2924 15570
rect 2976 15552 3004 16662
rect 3068 16454 3096 17070
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 3146 16416 3202 16425
rect 3068 16046 3096 16390
rect 3146 16351 3202 16360
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 2924 15524 3004 15552
rect 2872 15506 2924 15512
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2792 15094 2820 15438
rect 2780 15088 2832 15094
rect 2780 15030 2832 15036
rect 2792 14618 2820 15030
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2884 14260 2912 15506
rect 2964 15428 3016 15434
rect 2964 15370 3016 15376
rect 2976 14618 3004 15370
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 3068 14482 3096 15982
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 2884 14232 3096 14260
rect 2596 14000 2648 14006
rect 2596 13942 2648 13948
rect 2320 12368 2372 12374
rect 2320 12310 2372 12316
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2056 11218 2084 12242
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 1964 10010 1992 10610
rect 2056 10130 2084 11154
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2148 10810 2176 11086
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2240 10713 2268 12038
rect 2320 11756 2372 11762
rect 2608 11744 2636 13942
rect 2964 13796 3016 13802
rect 2884 13756 2964 13784
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2792 13394 2820 13670
rect 2884 13530 2912 13756
rect 2964 13738 3016 13744
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 3068 13394 3096 14232
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 2964 13252 3016 13258
rect 2964 13194 3016 13200
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2700 12850 2728 13126
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2870 12336 2926 12345
rect 2870 12271 2926 12280
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2608 11716 2728 11744
rect 2320 11698 2372 11704
rect 2226 10704 2282 10713
rect 2226 10639 2282 10648
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 1964 9982 2084 10010
rect 2056 9586 2084 9982
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 1872 9438 1992 9466
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1412 8974 1440 9318
rect 1872 9110 1900 9318
rect 1860 9104 1912 9110
rect 1860 9046 1912 9052
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1412 8480 1440 8910
rect 1412 8452 1532 8480
rect 1400 8356 1452 8362
rect 1400 8298 1452 8304
rect 1412 8265 1440 8298
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1504 7954 1532 8452
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1964 7818 1992 9438
rect 2228 9444 2280 9450
rect 2228 9386 2280 9392
rect 2240 9178 2268 9386
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 1952 7812 2004 7818
rect 1952 7754 2004 7760
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 7002 1624 7142
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1952 6724 2004 6730
rect 1952 6666 2004 6672
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1596 5778 1624 6598
rect 1964 6254 1992 6666
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1596 5166 1624 5714
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 1964 4690 1992 6054
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 1398 4176 1454 4185
rect 1398 4111 1400 4120
rect 1452 4111 1454 4120
rect 1400 4082 1452 4088
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1780 3738 1808 3878
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 2148 3466 2176 8298
rect 2240 8022 2268 9114
rect 2228 8016 2280 8022
rect 2228 7958 2280 7964
rect 2228 7812 2280 7818
rect 2228 7754 2280 7760
rect 2136 3460 2188 3466
rect 2136 3402 2188 3408
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 1596 2582 1624 2994
rect 1872 2990 1900 3334
rect 1860 2984 1912 2990
rect 1860 2926 1912 2932
rect 2240 2650 2268 7754
rect 2332 6914 2360 11698
rect 2504 11620 2556 11626
rect 2504 11562 2556 11568
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2424 10470 2452 11494
rect 2516 11218 2544 11562
rect 2608 11354 2636 11562
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2424 10198 2452 10406
rect 2412 10192 2464 10198
rect 2412 10134 2464 10140
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2608 9654 2636 10066
rect 2596 9648 2648 9654
rect 2596 9590 2648 9596
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2424 7188 2452 9522
rect 2700 9518 2728 11716
rect 2792 10742 2820 12038
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2504 8900 2556 8906
rect 2504 8842 2556 8848
rect 2516 8022 2544 8842
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2608 8634 2636 8774
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2608 8090 2636 8570
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2596 8084 2648 8090
rect 2596 8026 2648 8032
rect 2504 8016 2556 8022
rect 2504 7958 2556 7964
rect 2700 7954 2728 8366
rect 2792 8090 2820 8910
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2700 7546 2728 7890
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2884 7342 2912 12271
rect 2976 10538 3004 13194
rect 3068 10606 3096 13330
rect 3160 12850 3188 16351
rect 3252 14074 3280 19804
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 3344 16658 3372 17138
rect 3436 17134 3464 17818
rect 3654 17436 3950 17456
rect 3710 17434 3734 17436
rect 3790 17434 3814 17436
rect 3870 17434 3894 17436
rect 3732 17382 3734 17434
rect 3796 17382 3808 17434
rect 3870 17382 3872 17434
rect 3710 17380 3734 17382
rect 3790 17380 3814 17382
rect 3870 17380 3894 17382
rect 3654 17360 3950 17380
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 3332 16652 3384 16658
rect 3332 16594 3384 16600
rect 3344 15502 3372 16594
rect 3436 16114 3464 17070
rect 3654 16348 3950 16368
rect 3710 16346 3734 16348
rect 3790 16346 3814 16348
rect 3870 16346 3894 16348
rect 3732 16294 3734 16346
rect 3796 16294 3808 16346
rect 3870 16294 3872 16346
rect 3710 16292 3734 16294
rect 3790 16292 3814 16294
rect 3870 16292 3894 16294
rect 3654 16272 3950 16292
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 4172 15706 4200 15914
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 3332 15496 3384 15502
rect 3384 15456 3556 15484
rect 3332 15438 3384 15444
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 3344 14550 3372 14758
rect 3332 14544 3384 14550
rect 3332 14486 3384 14492
rect 3422 14376 3478 14385
rect 3422 14311 3478 14320
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 3332 13728 3384 13734
rect 3332 13670 3384 13676
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3146 12336 3202 12345
rect 3146 12271 3148 12280
rect 3200 12271 3202 12280
rect 3148 12242 3200 12248
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 3160 10130 3188 10610
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2688 7268 2740 7274
rect 2688 7210 2740 7216
rect 2504 7200 2556 7206
rect 2424 7160 2504 7188
rect 2504 7142 2556 7148
rect 2332 6886 2452 6914
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2332 5370 2360 5850
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2332 4078 2360 5306
rect 2424 5166 2452 6886
rect 2516 6798 2544 7142
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2516 6322 2544 6734
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2700 6254 2728 7210
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2424 4690 2452 5102
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2320 4072 2372 4078
rect 2320 4014 2372 4020
rect 2700 3602 2728 6190
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2780 5636 2832 5642
rect 2780 5578 2832 5584
rect 2792 5370 2820 5578
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2792 4146 2820 4558
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 1584 2576 1636 2582
rect 1584 2518 1636 2524
rect 1400 2372 1452 2378
rect 1400 2314 1452 2320
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1412 800 1440 2314
rect 2792 800 2820 3470
rect 2884 2145 2912 5714
rect 2976 2854 3004 9998
rect 3252 9518 3280 12922
rect 3344 12782 3372 13670
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3344 12306 3372 12582
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3148 8968 3200 8974
rect 3146 8936 3148 8945
rect 3200 8936 3202 8945
rect 3146 8871 3202 8880
rect 3160 8430 3188 8871
rect 3436 8514 3464 14311
rect 3528 13954 3556 15456
rect 3654 15260 3950 15280
rect 3710 15258 3734 15260
rect 3790 15258 3814 15260
rect 3870 15258 3894 15260
rect 3732 15206 3734 15258
rect 3796 15206 3808 15258
rect 3870 15206 3872 15258
rect 3710 15204 3734 15206
rect 3790 15204 3814 15206
rect 3870 15204 3894 15206
rect 3654 15184 3950 15204
rect 3988 15026 4016 15506
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 3654 14172 3950 14192
rect 3710 14170 3734 14172
rect 3790 14170 3814 14172
rect 3870 14170 3894 14172
rect 3732 14118 3734 14170
rect 3796 14118 3808 14170
rect 3870 14118 3872 14170
rect 3710 14116 3734 14118
rect 3790 14116 3814 14118
rect 3870 14116 3894 14118
rect 3654 14096 3950 14116
rect 3528 13926 3648 13954
rect 3516 13864 3568 13870
rect 3620 13841 3648 13926
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 3516 13806 3568 13812
rect 3606 13832 3662 13841
rect 3528 13462 3556 13806
rect 3606 13767 3662 13776
rect 3516 13456 3568 13462
rect 3516 13398 3568 13404
rect 3528 12986 3556 13398
rect 3620 13326 3648 13767
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 3654 13084 3950 13104
rect 3710 13082 3734 13084
rect 3790 13082 3814 13084
rect 3870 13082 3894 13084
rect 3732 13030 3734 13082
rect 3796 13030 3808 13082
rect 3870 13030 3872 13082
rect 3710 13028 3734 13030
rect 3790 13028 3814 13030
rect 3870 13028 3894 13030
rect 3654 13008 3950 13028
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3528 9586 3556 12786
rect 3988 12442 4016 13874
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 4080 12170 4108 13806
rect 4172 13802 4200 14758
rect 4264 14414 4292 16050
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4356 14958 4384 15302
rect 4344 14952 4396 14958
rect 4344 14894 4396 14900
rect 4252 14408 4304 14414
rect 4252 14350 4304 14356
rect 4356 14006 4384 14037
rect 4344 14000 4396 14006
rect 4342 13968 4344 13977
rect 4396 13968 4398 13977
rect 4342 13903 4398 13912
rect 4356 13870 4384 13903
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 4160 13796 4212 13802
rect 4160 13738 4212 13744
rect 4632 13734 4660 19804
rect 6012 17814 6040 19804
rect 6353 17980 6649 18000
rect 6409 17978 6433 17980
rect 6489 17978 6513 17980
rect 6569 17978 6593 17980
rect 6431 17926 6433 17978
rect 6495 17926 6507 17978
rect 6569 17926 6571 17978
rect 6409 17924 6433 17926
rect 6489 17924 6513 17926
rect 6569 17924 6593 17926
rect 6353 17904 6649 17924
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 5264 17536 5316 17542
rect 5264 17478 5316 17484
rect 4816 15978 4844 17478
rect 5276 17202 5304 17478
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5368 17134 5396 17614
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 5552 16522 5580 17682
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 5632 17604 5684 17610
rect 5632 17546 5684 17552
rect 5540 16516 5592 16522
rect 5540 16458 5592 16464
rect 4804 15972 4856 15978
rect 4804 15914 4856 15920
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 4894 13832 4950 13841
rect 4894 13767 4950 13776
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4264 12442 4292 13466
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 4252 12436 4304 12442
rect 4356 12434 4384 13194
rect 4632 12782 4660 13330
rect 4816 12850 4844 13398
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4356 12406 4476 12434
rect 4252 12378 4304 12384
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 3654 11996 3950 12016
rect 3710 11994 3734 11996
rect 3790 11994 3814 11996
rect 3870 11994 3894 11996
rect 3732 11942 3734 11994
rect 3796 11942 3808 11994
rect 3870 11942 3872 11994
rect 3710 11940 3734 11942
rect 3790 11940 3814 11942
rect 3870 11940 3894 11942
rect 3654 11920 3950 11940
rect 3654 10908 3950 10928
rect 3710 10906 3734 10908
rect 3790 10906 3814 10908
rect 3870 10906 3894 10908
rect 3732 10854 3734 10906
rect 3796 10854 3808 10906
rect 3870 10854 3872 10906
rect 3710 10852 3734 10854
rect 3790 10852 3814 10854
rect 3870 10852 3894 10854
rect 3654 10832 3950 10852
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 3654 9820 3950 9840
rect 3710 9818 3734 9820
rect 3790 9818 3814 9820
rect 3870 9818 3894 9820
rect 3732 9766 3734 9818
rect 3796 9766 3808 9818
rect 3870 9766 3872 9818
rect 3710 9764 3734 9766
rect 3790 9764 3814 9766
rect 3870 9764 3894 9766
rect 3654 9744 3950 9764
rect 3988 9586 4016 10542
rect 4080 10198 4108 12106
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4264 11914 4292 12038
rect 4172 11898 4292 11914
rect 4160 11892 4292 11898
rect 4212 11886 4292 11892
rect 4160 11834 4212 11840
rect 4172 11694 4200 11834
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 4172 10810 4200 11222
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4080 9722 4108 10134
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 9178 3648 9318
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3654 8732 3950 8752
rect 3710 8730 3734 8732
rect 3790 8730 3814 8732
rect 3870 8730 3894 8732
rect 3732 8678 3734 8730
rect 3796 8678 3808 8730
rect 3870 8678 3872 8730
rect 3710 8676 3734 8678
rect 3790 8676 3814 8678
rect 3870 8676 3894 8678
rect 3654 8656 3950 8676
rect 3436 8486 3556 8514
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3068 6866 3096 7278
rect 3332 7268 3384 7274
rect 3332 7210 3384 7216
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 3344 6662 3372 7210
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3054 6216 3110 6225
rect 3054 6151 3110 6160
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 3068 2514 3096 6151
rect 3528 4826 3556 8486
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 3654 7644 3950 7664
rect 3710 7642 3734 7644
rect 3790 7642 3814 7644
rect 3870 7642 3894 7644
rect 3732 7590 3734 7642
rect 3796 7590 3808 7642
rect 3870 7590 3872 7642
rect 3710 7588 3734 7590
rect 3790 7588 3814 7590
rect 3870 7588 3894 7590
rect 3654 7568 3950 7588
rect 4172 7274 4200 7890
rect 4264 7478 4292 8230
rect 4356 8106 4384 10950
rect 4448 8498 4476 12406
rect 4724 12306 4752 12718
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4540 11762 4568 11834
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4632 11694 4660 12038
rect 4908 11898 4936 13767
rect 5000 12918 5028 14214
rect 5092 14074 5120 14758
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 5092 13394 5120 14010
rect 5184 13977 5212 14962
rect 5644 14958 5672 17546
rect 5736 17270 5764 17614
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 5724 17264 5776 17270
rect 5724 17206 5776 17212
rect 5736 16726 5764 17206
rect 6353 16892 6649 16912
rect 6409 16890 6433 16892
rect 6489 16890 6513 16892
rect 6569 16890 6593 16892
rect 6431 16838 6433 16890
rect 6495 16838 6507 16890
rect 6569 16838 6571 16890
rect 6409 16836 6433 16838
rect 6489 16836 6513 16838
rect 6569 16836 6593 16838
rect 6353 16816 6649 16836
rect 5724 16720 5776 16726
rect 5724 16662 5776 16668
rect 5736 16046 5764 16662
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6000 16516 6052 16522
rect 6000 16458 6052 16464
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5724 15632 5776 15638
rect 6012 15609 6040 16458
rect 6104 16114 6132 16526
rect 6932 16454 6960 17274
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6276 16108 6328 16114
rect 6276 16050 6328 16056
rect 6184 15972 6236 15978
rect 6184 15914 6236 15920
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 5724 15574 5776 15580
rect 5998 15600 6054 15609
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5276 14074 5304 14350
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5170 13968 5226 13977
rect 5170 13903 5226 13912
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 4988 12912 5040 12918
rect 4988 12854 5040 12860
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 4908 11801 4936 11834
rect 4894 11792 4950 11801
rect 4894 11727 4950 11736
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4540 10810 4568 11086
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4908 10674 4936 11494
rect 5000 11014 5028 12854
rect 5080 12776 5132 12782
rect 5184 12764 5212 13903
rect 5632 13796 5684 13802
rect 5632 13738 5684 13744
rect 5644 13326 5672 13738
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5644 12918 5672 13262
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5132 12736 5212 12764
rect 5080 12718 5132 12724
rect 5092 12238 5120 12718
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 5092 11762 5120 12174
rect 5368 11898 5396 12242
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5368 11626 5396 11834
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5552 10470 5580 10610
rect 5644 10606 5672 12106
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5644 9738 5672 9930
rect 5552 9710 5672 9738
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4356 8078 4476 8106
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 4356 6882 4384 7686
rect 4264 6854 4384 6882
rect 4264 6798 4292 6854
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 3654 6556 3950 6576
rect 3710 6554 3734 6556
rect 3790 6554 3814 6556
rect 3870 6554 3894 6556
rect 3732 6502 3734 6554
rect 3796 6502 3808 6554
rect 3870 6502 3872 6554
rect 3710 6500 3734 6502
rect 3790 6500 3814 6502
rect 3870 6500 3894 6502
rect 3654 6480 3950 6500
rect 4080 6458 4108 6734
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4356 6322 4384 6666
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 3654 5468 3950 5488
rect 3710 5466 3734 5468
rect 3790 5466 3814 5468
rect 3870 5466 3894 5468
rect 3732 5414 3734 5466
rect 3796 5414 3808 5466
rect 3870 5414 3872 5466
rect 3710 5412 3734 5414
rect 3790 5412 3814 5414
rect 3870 5412 3894 5414
rect 3654 5392 3950 5412
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3160 3670 3188 4422
rect 3654 4380 3950 4400
rect 3710 4378 3734 4380
rect 3790 4378 3814 4380
rect 3870 4378 3894 4380
rect 3732 4326 3734 4378
rect 3796 4326 3808 4378
rect 3870 4326 3872 4378
rect 3710 4324 3734 4326
rect 3790 4324 3814 4326
rect 3870 4324 3894 4326
rect 3654 4304 3950 4324
rect 4172 4078 4200 4966
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 3516 4004 3568 4010
rect 3516 3946 3568 3952
rect 3148 3664 3200 3670
rect 3332 3664 3384 3670
rect 3148 3606 3200 3612
rect 3330 3632 3332 3641
rect 3384 3632 3386 3641
rect 3330 3567 3386 3576
rect 3528 3398 3556 3946
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3654 3292 3950 3312
rect 3710 3290 3734 3292
rect 3790 3290 3814 3292
rect 3870 3290 3894 3292
rect 3732 3238 3734 3290
rect 3796 3238 3808 3290
rect 3870 3238 3872 3290
rect 3710 3236 3734 3238
rect 3790 3236 3814 3238
rect 3870 3236 3894 3238
rect 3654 3216 3950 3236
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 3654 2204 3950 2224
rect 3710 2202 3734 2204
rect 3790 2202 3814 2204
rect 3870 2202 3894 2204
rect 3732 2150 3734 2202
rect 3796 2150 3808 2202
rect 3870 2150 3872 2202
rect 3710 2148 3734 2150
rect 3790 2148 3814 2150
rect 3870 2148 3894 2150
rect 2870 2136 2926 2145
rect 3654 2128 3950 2148
rect 2870 2071 2926 2080
rect 4172 800 4200 2994
rect 4264 2650 4292 6054
rect 4448 4146 4476 8078
rect 4632 6866 4660 8774
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4528 6248 4580 6254
rect 4632 6236 4660 6802
rect 4724 6730 4752 7278
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 4724 6254 4752 6666
rect 4580 6208 4660 6236
rect 4712 6248 4764 6254
rect 4528 6190 4580 6196
rect 4712 6190 4764 6196
rect 4816 5914 4844 9454
rect 5000 8498 5028 9454
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5092 8634 5120 8910
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5368 8498 5396 8910
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5368 7886 5396 8434
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5460 7290 5488 8774
rect 5552 8430 5580 9710
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5644 8498 5672 9386
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5552 7410 5580 7890
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5644 7342 5672 8434
rect 5736 8090 5764 15574
rect 5998 15535 6000 15544
rect 6052 15535 6054 15544
rect 6000 15506 6052 15512
rect 6104 15450 6132 15846
rect 6196 15638 6224 15914
rect 6184 15632 6236 15638
rect 6184 15574 6236 15580
rect 6288 15502 6316 16050
rect 6353 15804 6649 15824
rect 6409 15802 6433 15804
rect 6489 15802 6513 15804
rect 6569 15802 6593 15804
rect 6431 15750 6433 15802
rect 6495 15750 6507 15802
rect 6569 15750 6571 15802
rect 6409 15748 6433 15750
rect 6489 15748 6513 15750
rect 6569 15748 6593 15750
rect 6353 15728 6649 15748
rect 6932 15570 6960 16390
rect 7392 16232 7420 19804
rect 8772 18086 8800 19804
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 8484 17740 8536 17746
rect 8484 17682 8536 17688
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 7668 17134 7696 17682
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 7852 17134 7880 17478
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7576 16726 7604 16934
rect 7564 16720 7616 16726
rect 7564 16662 7616 16668
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 7392 16204 7604 16232
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7300 15609 7328 15982
rect 7286 15600 7342 15609
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 7196 15564 7248 15570
rect 7286 15535 7342 15544
rect 7196 15506 7248 15512
rect 6012 15422 6132 15450
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 6736 15428 6788 15434
rect 5908 14000 5960 14006
rect 5908 13942 5960 13948
rect 5920 13394 5948 13942
rect 6012 13870 6040 15422
rect 6736 15370 6788 15376
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6092 14272 6144 14278
rect 6092 14214 6144 14220
rect 6000 13864 6052 13870
rect 5998 13832 6000 13841
rect 6052 13832 6054 13841
rect 6104 13802 6132 14214
rect 5998 13767 6054 13776
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 6104 13394 6132 13738
rect 5908 13388 5960 13394
rect 5908 13330 5960 13336
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 5920 13258 5948 13330
rect 5908 13252 5960 13258
rect 5908 13194 5960 13200
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5828 12345 5856 13126
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 5814 12336 5870 12345
rect 5814 12271 5870 12280
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5828 11937 5856 12038
rect 5814 11928 5870 11937
rect 5814 11863 5870 11872
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5828 11014 5856 11562
rect 5816 11008 5868 11014
rect 5816 10950 5868 10956
rect 5828 10606 5856 10950
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5828 10282 5856 10542
rect 5920 10470 5948 11630
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5828 10254 5948 10282
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 5828 9178 5856 9862
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5828 8634 5856 8978
rect 5920 8820 5948 10254
rect 6012 9926 6040 12786
rect 6104 12374 6132 13330
rect 6184 13252 6236 13258
rect 6184 13194 6236 13200
rect 6092 12368 6144 12374
rect 6092 12310 6144 12316
rect 6196 12102 6224 13194
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 6196 11898 6224 12038
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6288 11642 6316 15302
rect 6748 14958 6776 15370
rect 6932 14958 6960 15506
rect 7208 15162 7236 15506
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6353 14716 6649 14736
rect 6409 14714 6433 14716
rect 6489 14714 6513 14716
rect 6569 14714 6593 14716
rect 6431 14662 6433 14714
rect 6495 14662 6507 14714
rect 6569 14662 6571 14714
rect 6409 14660 6433 14662
rect 6489 14660 6513 14662
rect 6569 14660 6593 14662
rect 6353 14640 6649 14660
rect 7208 14414 7236 15098
rect 7300 15094 7328 15535
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7288 15088 7340 15094
rect 7288 15030 7340 15036
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7392 14278 7420 15438
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6353 13628 6649 13648
rect 6409 13626 6433 13628
rect 6489 13626 6513 13628
rect 6569 13626 6593 13628
rect 6431 13574 6433 13626
rect 6495 13574 6507 13626
rect 6569 13574 6571 13626
rect 6409 13572 6433 13574
rect 6489 13572 6513 13574
rect 6569 13572 6593 13574
rect 6353 13552 6649 13572
rect 6748 13394 6776 14010
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 7012 13796 7064 13802
rect 7064 13756 7144 13784
rect 7012 13738 7064 13744
rect 7116 13462 7144 13756
rect 7208 13530 7236 13874
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7104 13456 7156 13462
rect 7104 13398 7156 13404
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 6748 13190 6776 13330
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 7024 12986 7052 13330
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6353 12540 6649 12560
rect 6409 12538 6433 12540
rect 6489 12538 6513 12540
rect 6569 12538 6593 12540
rect 6431 12486 6433 12538
rect 6495 12486 6507 12538
rect 6569 12486 6571 12538
rect 6409 12484 6433 12486
rect 6489 12484 6513 12486
rect 6569 12484 6593 12486
rect 6353 12464 6649 12484
rect 6644 12368 6696 12374
rect 6550 12336 6606 12345
rect 6644 12310 6696 12316
rect 6550 12271 6552 12280
rect 6604 12271 6606 12280
rect 6552 12242 6604 12248
rect 6550 12200 6606 12209
rect 6368 12164 6420 12170
rect 6550 12135 6552 12144
rect 6368 12106 6420 12112
rect 6604 12135 6606 12144
rect 6552 12106 6604 12112
rect 6104 11614 6316 11642
rect 6380 11626 6408 12106
rect 6368 11620 6420 11626
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 6000 8832 6052 8838
rect 5920 8792 6000 8820
rect 6000 8774 6052 8780
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5828 8498 5948 8514
rect 5828 8492 5960 8498
rect 5828 8486 5908 8492
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5828 7954 5856 8486
rect 5908 8434 5960 8440
rect 6012 8430 6040 8774
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5632 7336 5684 7342
rect 5460 7262 5580 7290
rect 5632 7278 5684 7284
rect 5736 7274 5764 7822
rect 5920 7546 5948 7822
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5460 6458 5488 6938
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4618 5808 4674 5817
rect 4618 5743 4620 5752
rect 4672 5743 4674 5752
rect 4620 5714 4672 5720
rect 4816 5234 4844 5850
rect 4908 5846 4936 6326
rect 5552 6236 5580 7262
rect 5724 7268 5776 7274
rect 5724 7210 5776 7216
rect 5632 6248 5684 6254
rect 5552 6208 5632 6236
rect 5632 6190 5684 6196
rect 4896 5840 4948 5846
rect 4896 5782 4948 5788
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4816 4078 4844 5170
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4908 2774 4936 5782
rect 5644 5778 5672 6190
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5736 5710 5764 7210
rect 5920 6866 5948 7278
rect 6012 6866 6040 8230
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6012 6254 6040 6802
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5276 5166 5304 5646
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 5092 4622 5120 5034
rect 5920 4690 5948 5510
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 5552 4146 5580 4626
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5920 4078 5948 4626
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 4816 2746 4936 2774
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4816 2514 4844 2746
rect 5092 2650 5120 2858
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 5552 800 5580 3130
rect 5644 2650 5672 3606
rect 5814 3496 5870 3505
rect 5814 3431 5870 3440
rect 5828 2854 5856 3431
rect 6104 3194 6132 11614
rect 6368 11562 6420 11568
rect 6184 11552 6236 11558
rect 6656 11540 6684 12310
rect 6748 11801 6776 12718
rect 7024 12209 7052 12922
rect 7010 12200 7066 12209
rect 7010 12135 7066 12144
rect 7010 11928 7066 11937
rect 7010 11863 7066 11872
rect 6734 11792 6790 11801
rect 6734 11727 6790 11736
rect 6748 11694 6776 11727
rect 7024 11694 7052 11863
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 6656 11512 6776 11540
rect 6184 11494 6236 11500
rect 6196 10810 6224 11494
rect 6353 11452 6649 11472
rect 6409 11450 6433 11452
rect 6489 11450 6513 11452
rect 6569 11450 6593 11452
rect 6431 11398 6433 11450
rect 6495 11398 6507 11450
rect 6569 11398 6571 11450
rect 6409 11396 6433 11398
rect 6489 11396 6513 11398
rect 6569 11396 6593 11398
rect 6353 11376 6649 11396
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6196 10062 6224 10406
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6196 8022 6224 9998
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6196 2990 6224 3130
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 6288 2650 6316 10610
rect 6748 10606 6776 11512
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6353 10364 6649 10384
rect 6409 10362 6433 10364
rect 6489 10362 6513 10364
rect 6569 10362 6593 10364
rect 6431 10310 6433 10362
rect 6495 10310 6507 10362
rect 6569 10310 6571 10362
rect 6409 10308 6433 10310
rect 6489 10308 6513 10310
rect 6569 10308 6593 10310
rect 6353 10288 6649 10308
rect 6748 9926 6776 10542
rect 6840 10062 6868 10950
rect 7116 10810 7144 13398
rect 7380 13252 7432 13258
rect 7380 13194 7432 13200
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7208 12306 7236 13126
rect 7392 12782 7420 13194
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7484 12442 7512 12650
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7300 11694 7328 12378
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7392 11762 7420 12174
rect 7484 12170 7512 12378
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7208 11218 7236 11290
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7300 11082 7328 11630
rect 7392 11218 7420 11698
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6748 9722 6776 9862
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6353 9276 6649 9296
rect 6409 9274 6433 9276
rect 6489 9274 6513 9276
rect 6569 9274 6593 9276
rect 6431 9222 6433 9274
rect 6495 9222 6507 9274
rect 6569 9222 6571 9274
rect 6409 9220 6433 9222
rect 6489 9220 6513 9222
rect 6569 9220 6593 9222
rect 6353 9200 6649 9220
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6736 9036 6788 9042
rect 6840 9024 6868 9998
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6932 9042 6960 9930
rect 7116 9926 7144 10746
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7392 10130 7420 10202
rect 7484 10130 7512 11290
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7208 9450 7236 10066
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7024 9353 7052 9386
rect 7010 9344 7066 9353
rect 7010 9279 7066 9288
rect 6788 8996 6868 9024
rect 6920 9036 6972 9042
rect 6736 8978 6788 8984
rect 6920 8978 6972 8984
rect 6380 8362 6408 8978
rect 6552 8900 6604 8906
rect 6552 8842 6604 8848
rect 6564 8498 6592 8842
rect 6748 8838 6776 8978
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6932 8362 6960 8978
rect 7024 8430 7052 9279
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7116 9042 7144 9114
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6353 8188 6649 8208
rect 6409 8186 6433 8188
rect 6489 8186 6513 8188
rect 6569 8186 6593 8188
rect 6431 8134 6433 8186
rect 6495 8134 6507 8186
rect 6569 8134 6571 8186
rect 6409 8132 6433 8134
rect 6489 8132 6513 8134
rect 6569 8132 6593 8134
rect 6353 8112 6649 8132
rect 7116 7954 7144 8434
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6353 7100 6649 7120
rect 6409 7098 6433 7100
rect 6489 7098 6513 7100
rect 6569 7098 6593 7100
rect 6431 7046 6433 7098
rect 6495 7046 6507 7098
rect 6569 7046 6571 7098
rect 6409 7044 6433 7046
rect 6489 7044 6513 7046
rect 6569 7044 6593 7046
rect 6353 7024 6649 7044
rect 6353 6012 6649 6032
rect 6409 6010 6433 6012
rect 6489 6010 6513 6012
rect 6569 6010 6593 6012
rect 6431 5958 6433 6010
rect 6495 5958 6507 6010
rect 6569 5958 6571 6010
rect 6409 5956 6433 5958
rect 6489 5956 6513 5958
rect 6569 5956 6593 5958
rect 6353 5936 6649 5956
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6472 5234 6500 5646
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6353 4924 6649 4944
rect 6409 4922 6433 4924
rect 6489 4922 6513 4924
rect 6569 4922 6593 4924
rect 6431 4870 6433 4922
rect 6495 4870 6507 4922
rect 6569 4870 6571 4922
rect 6409 4868 6433 4870
rect 6489 4868 6513 4870
rect 6569 4868 6593 4870
rect 6353 4848 6649 4868
rect 6353 3836 6649 3856
rect 6409 3834 6433 3836
rect 6489 3834 6513 3836
rect 6569 3834 6593 3836
rect 6431 3782 6433 3834
rect 6495 3782 6507 3834
rect 6569 3782 6571 3834
rect 6409 3780 6433 3782
rect 6489 3780 6513 3782
rect 6569 3780 6593 3782
rect 6353 3760 6649 3780
rect 6748 3602 6776 7686
rect 6932 6934 6960 7686
rect 7208 7478 7236 8026
rect 7196 7472 7248 7478
rect 7196 7414 7248 7420
rect 7300 7324 7328 8366
rect 7392 8022 7420 10066
rect 7484 9586 7512 10066
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7484 8430 7512 8774
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7484 7886 7512 8366
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7380 7336 7432 7342
rect 7300 7296 7380 7324
rect 7380 7278 7432 7284
rect 6920 6928 6972 6934
rect 6920 6870 6972 6876
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6840 5166 6868 6054
rect 6932 5914 6960 6870
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7024 5642 7052 6666
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7300 6322 7328 6598
rect 7392 6390 7420 7278
rect 7576 6866 7604 16204
rect 8036 16046 8064 16390
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 8312 15570 8340 16186
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 7932 14884 7984 14890
rect 7932 14826 7984 14832
rect 8024 14884 8076 14890
rect 8024 14826 8076 14832
rect 7944 14074 7972 14826
rect 8036 14618 8064 14826
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 8024 14476 8076 14482
rect 8128 14464 8156 15438
rect 8404 14958 8432 17478
rect 8496 16046 8524 17682
rect 9052 17436 9348 17456
rect 9108 17434 9132 17436
rect 9188 17434 9212 17436
rect 9268 17434 9292 17436
rect 9130 17382 9132 17434
rect 9194 17382 9206 17434
rect 9268 17382 9270 17434
rect 9108 17380 9132 17382
rect 9188 17380 9212 17382
rect 9268 17380 9292 17382
rect 9052 17360 9348 17380
rect 9052 16348 9348 16368
rect 9108 16346 9132 16348
rect 9188 16346 9212 16348
rect 9268 16346 9292 16348
rect 9130 16294 9132 16346
rect 9194 16294 9206 16346
rect 9268 16294 9270 16346
rect 9108 16292 9132 16294
rect 9188 16292 9212 16294
rect 9268 16292 9292 16294
rect 9052 16272 9348 16292
rect 9600 16182 9628 17682
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9588 16176 9640 16182
rect 9588 16118 9640 16124
rect 9692 16114 9720 17478
rect 9784 16794 9812 17682
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9784 16250 9812 16730
rect 9876 16658 9904 17002
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8680 15502 8708 16050
rect 9692 15552 9720 16050
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9784 15706 9812 15982
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9692 15524 9812 15552
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8760 15428 8812 15434
rect 8760 15370 8812 15376
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 8772 15314 8800 15370
rect 8680 15286 8800 15314
rect 8392 14952 8444 14958
rect 8392 14894 8444 14900
rect 8392 14544 8444 14550
rect 8392 14486 8444 14492
rect 8076 14436 8156 14464
rect 8024 14418 8076 14424
rect 8128 14074 8156 14436
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8220 14006 8248 14418
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8404 13938 8432 14486
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7668 13462 7696 13670
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7668 12782 7696 13398
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7852 12986 7880 13262
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7944 12850 7972 13466
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8128 12918 8156 13262
rect 8116 12912 8168 12918
rect 8116 12854 8168 12860
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7852 12434 7880 12582
rect 7668 12406 7880 12434
rect 7668 12306 7696 12406
rect 7840 12368 7892 12374
rect 7840 12310 7892 12316
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 7668 10062 7696 12242
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7760 11286 7788 12038
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7852 10266 7880 12310
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8036 11150 8064 11494
rect 8128 11218 8156 12854
rect 8220 12306 8248 13330
rect 8496 12714 8524 14350
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 8208 12300 8260 12306
rect 8260 12260 8340 12288
rect 8208 12242 8260 12248
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 8312 10130 8340 12260
rect 8496 11694 8524 12650
rect 8680 12442 8708 15286
rect 9052 15260 9348 15280
rect 9108 15258 9132 15260
rect 9188 15258 9212 15260
rect 9268 15258 9292 15260
rect 9130 15206 9132 15258
rect 9194 15206 9206 15258
rect 9268 15206 9270 15258
rect 9108 15204 9132 15206
rect 9188 15204 9212 15206
rect 9268 15204 9292 15206
rect 9052 15184 9348 15204
rect 9692 14958 9720 15370
rect 9784 15026 9812 15524
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 8772 14618 8800 14894
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8772 13938 8800 14554
rect 9876 14414 9904 16594
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 9968 15638 9996 16526
rect 10152 16454 10180 19804
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 10416 17332 10468 17338
rect 10416 17274 10468 17280
rect 10428 17218 10456 17274
rect 10428 17190 10640 17218
rect 10428 17134 10456 17190
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10520 16658 10548 17070
rect 10508 16652 10560 16658
rect 10508 16594 10560 16600
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10232 16516 10284 16522
rect 10232 16458 10284 16464
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10244 15638 10272 16458
rect 10428 15706 10456 16526
rect 10612 15706 10640 17190
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10692 15972 10744 15978
rect 10692 15914 10744 15920
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 9968 15162 9996 15574
rect 10704 15366 10732 15914
rect 10888 15858 10916 17070
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10980 16046 11008 16594
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10888 15830 11008 15858
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9968 14482 9996 14962
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10244 14482 10272 14758
rect 10336 14618 10364 14894
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9052 14172 9348 14192
rect 9108 14170 9132 14172
rect 9188 14170 9212 14172
rect 9268 14170 9292 14172
rect 9130 14118 9132 14170
rect 9194 14118 9206 14170
rect 9268 14118 9270 14170
rect 9108 14116 9132 14118
rect 9188 14116 9212 14118
rect 9268 14116 9292 14118
rect 9052 14096 9348 14116
rect 9784 14074 9812 14214
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 9784 13734 9812 14010
rect 10244 13802 10272 14418
rect 10704 13938 10732 14894
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10232 13796 10284 13802
rect 10232 13738 10284 13744
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 10704 13530 10732 13874
rect 10888 13852 10916 15642
rect 10980 15094 11008 15830
rect 11072 15094 11100 17478
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 11164 16726 11192 17002
rect 11348 16726 11376 17478
rect 11152 16720 11204 16726
rect 11152 16662 11204 16668
rect 11336 16720 11388 16726
rect 11336 16662 11388 16668
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11256 16182 11284 16594
rect 11440 16250 11468 16594
rect 11532 16538 11560 19804
rect 11750 17980 12046 18000
rect 11806 17978 11830 17980
rect 11886 17978 11910 17980
rect 11966 17978 11990 17980
rect 11828 17926 11830 17978
rect 11892 17926 11904 17978
rect 11966 17926 11968 17978
rect 11806 17924 11830 17926
rect 11886 17924 11910 17926
rect 11966 17924 11990 17926
rect 11750 17904 12046 17924
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 11750 16892 12046 16912
rect 11806 16890 11830 16892
rect 11886 16890 11910 16892
rect 11966 16890 11990 16892
rect 11828 16838 11830 16890
rect 11892 16838 11904 16890
rect 11966 16838 11968 16890
rect 11806 16836 11830 16838
rect 11886 16836 11910 16838
rect 11966 16836 11990 16838
rect 11750 16816 12046 16836
rect 12268 16794 12296 16934
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12164 16584 12216 16590
rect 11532 16510 11652 16538
rect 12164 16526 12216 16532
rect 11520 16448 11572 16454
rect 11520 16390 11572 16396
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 11244 16176 11296 16182
rect 11244 16118 11296 16124
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 10980 14940 11008 15030
rect 10980 14912 11100 14940
rect 10968 14544 11020 14550
rect 10968 14486 11020 14492
rect 10980 14074 11008 14486
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 11072 14006 11100 14912
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11060 14000 11112 14006
rect 11164 13988 11192 14214
rect 11112 13960 11192 13988
rect 11060 13942 11112 13948
rect 10968 13864 11020 13870
rect 10888 13824 10968 13852
rect 10968 13806 11020 13812
rect 10980 13530 11008 13806
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 9052 13084 9348 13104
rect 9108 13082 9132 13084
rect 9188 13082 9212 13084
rect 9268 13082 9292 13084
rect 9130 13030 9132 13082
rect 9194 13030 9206 13082
rect 9268 13030 9270 13082
rect 9108 13028 9132 13030
rect 9188 13028 9212 13030
rect 9268 13028 9292 13030
rect 9052 13008 9348 13028
rect 10888 12850 10916 13466
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 9508 12306 9536 12582
rect 10796 12306 10824 12718
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 9052 11996 9348 12016
rect 9108 11994 9132 11996
rect 9188 11994 9212 11996
rect 9268 11994 9292 11996
rect 9130 11942 9132 11994
rect 9194 11942 9206 11994
rect 9268 11942 9270 11994
rect 9108 11940 9132 11942
rect 9188 11940 9212 11942
rect 9268 11940 9292 11942
rect 9052 11920 9348 11940
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8496 11286 8524 11630
rect 8760 11620 8812 11626
rect 8760 11562 8812 11568
rect 8772 11354 8800 11562
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8484 11280 8536 11286
rect 8484 11222 8536 11228
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9968 11150 9996 11222
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9052 10908 9348 10928
rect 9108 10906 9132 10908
rect 9188 10906 9212 10908
rect 9268 10906 9292 10908
rect 9130 10854 9132 10906
rect 9194 10854 9206 10906
rect 9268 10854 9270 10906
rect 9108 10852 9132 10854
rect 9188 10852 9212 10854
rect 9268 10852 9292 10854
rect 9052 10832 9348 10852
rect 9876 10810 9904 11086
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 8666 10704 8722 10713
rect 8666 10639 8668 10648
rect 8720 10639 8722 10648
rect 8760 10668 8812 10674
rect 8668 10610 8720 10616
rect 8760 10610 8812 10616
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8588 10266 8616 10406
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7760 8430 7788 9522
rect 8128 9518 8156 9862
rect 7932 9512 7984 9518
rect 7930 9480 7932 9489
rect 8116 9512 8168 9518
rect 7984 9480 7986 9489
rect 8116 9454 8168 9460
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 7930 9415 7986 9424
rect 8024 9444 8076 9450
rect 8024 9386 8076 9392
rect 8036 8974 8064 9386
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7852 8430 7880 8570
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7944 8294 7972 8910
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 8634 8064 8774
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8128 8498 8156 9454
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8220 8362 8248 9454
rect 8312 9042 8340 9930
rect 8576 9376 8628 9382
rect 8628 9336 8708 9364
rect 8576 9318 8628 9324
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8312 8566 8340 8978
rect 8484 8968 8536 8974
rect 8482 8936 8484 8945
rect 8536 8936 8538 8945
rect 8680 8906 8708 9336
rect 8482 8871 8538 8880
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 7944 7886 7972 8230
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7760 7410 7788 7686
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 8036 6798 8064 8230
rect 8312 7342 8340 8502
rect 8680 8022 8708 8842
rect 8772 8430 8800 10610
rect 10244 10606 10272 11494
rect 10888 11354 10916 12786
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10888 10606 10916 11290
rect 10980 10674 11008 13466
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11072 12986 11100 13126
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 11164 10606 11192 13960
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9404 10192 9456 10198
rect 9404 10134 9456 10140
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 8680 7546 8708 7958
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8300 7336 8352 7342
rect 8576 7336 8628 7342
rect 8300 7278 8352 7284
rect 8404 7296 8576 7324
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8220 7002 8248 7142
rect 8312 7002 8340 7278
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7392 6186 7420 6326
rect 8036 6322 8064 6734
rect 8220 6458 8248 6734
rect 8404 6458 8432 7296
rect 8576 7278 8628 7284
rect 8588 7206 8616 7278
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8484 6928 8536 6934
rect 8484 6870 8536 6876
rect 8496 6730 8524 6870
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 7300 5574 7328 6054
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7668 5817 7696 5850
rect 7654 5808 7710 5817
rect 7654 5743 7710 5752
rect 7760 5710 7788 6190
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6840 4146 6868 5102
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 7208 3942 7236 5306
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7392 4758 7420 5102
rect 7380 4752 7432 4758
rect 7380 4694 7432 4700
rect 7392 4570 7420 4694
rect 7472 4684 7524 4690
rect 7576 4672 7604 5578
rect 8036 5234 8064 6258
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 8128 5166 8156 6054
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8220 5370 8248 5714
rect 8404 5574 8432 6394
rect 8588 6322 8616 6598
rect 8680 6458 8708 7482
rect 8956 7342 8984 9998
rect 9052 9820 9348 9840
rect 9108 9818 9132 9820
rect 9188 9818 9212 9820
rect 9268 9818 9292 9820
rect 9130 9766 9132 9818
rect 9194 9766 9206 9818
rect 9268 9766 9270 9818
rect 9108 9764 9132 9766
rect 9188 9764 9212 9766
rect 9268 9764 9292 9766
rect 9052 9744 9348 9764
rect 9036 9376 9088 9382
rect 9034 9344 9036 9353
rect 9088 9344 9090 9353
rect 9034 9279 9090 9288
rect 9416 9042 9444 10134
rect 9692 9994 9720 10406
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9692 9586 9720 9930
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9508 9178 9536 9386
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9052 8732 9348 8752
rect 9108 8730 9132 8732
rect 9188 8730 9212 8732
rect 9268 8730 9292 8732
rect 9130 8678 9132 8730
rect 9194 8678 9206 8730
rect 9268 8678 9270 8730
rect 9108 8676 9132 8678
rect 9188 8676 9212 8678
rect 9268 8676 9292 8678
rect 9052 8656 9348 8676
rect 9600 8566 9628 9454
rect 9692 9042 9720 9522
rect 9784 9518 9812 9862
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9876 8906 9904 10202
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9968 9042 9996 10066
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 10060 9722 10088 9862
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9772 8832 9824 8838
rect 9824 8780 9904 8786
rect 9772 8774 9904 8780
rect 9784 8758 9904 8774
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9052 7644 9348 7664
rect 9108 7642 9132 7644
rect 9188 7642 9212 7644
rect 9268 7642 9292 7644
rect 9130 7590 9132 7642
rect 9194 7590 9206 7642
rect 9268 7590 9270 7642
rect 9108 7588 9132 7590
rect 9188 7588 9212 7590
rect 9268 7588 9292 7590
rect 9052 7568 9348 7588
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8496 6118 8524 6190
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8496 5710 8524 6054
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7524 4644 7604 4672
rect 7472 4626 7524 4632
rect 7392 4542 7512 4570
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7392 4214 7420 4422
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 6918 3768 6974 3777
rect 6918 3703 6974 3712
rect 6932 3670 6960 3703
rect 7484 3670 7512 4542
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6368 3528 6420 3534
rect 6366 3496 6368 3505
rect 6420 3496 6422 3505
rect 6366 3431 6422 3440
rect 6748 2990 6776 3538
rect 7484 2990 7512 3606
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 6353 2748 6649 2768
rect 6409 2746 6433 2748
rect 6489 2746 6513 2748
rect 6569 2746 6593 2748
rect 6431 2694 6433 2746
rect 6495 2694 6507 2746
rect 6569 2694 6571 2746
rect 6409 2692 6433 2694
rect 6489 2692 6513 2694
rect 6569 2692 6593 2694
rect 6353 2672 6649 2692
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 7208 2446 7236 2790
rect 7668 2446 7696 3334
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 6932 800 6960 2382
rect 7760 2378 7788 4966
rect 8036 4690 8064 5034
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8588 4690 8616 4966
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 7944 3670 7972 4150
rect 8036 4078 8064 4422
rect 8588 4146 8616 4626
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 8036 3942 8064 4014
rect 8680 4010 8708 4966
rect 8668 4004 8720 4010
rect 8668 3946 8720 3952
rect 8760 4004 8812 4010
rect 8760 3946 8812 3952
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 8772 3777 8800 3946
rect 8758 3768 8814 3777
rect 8758 3703 8814 3712
rect 7932 3664 7984 3670
rect 8392 3664 8444 3670
rect 7932 3606 7984 3612
rect 8390 3632 8392 3641
rect 8444 3632 8446 3641
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7852 2514 7880 2790
rect 7944 2582 7972 3606
rect 8208 3596 8260 3602
rect 8390 3567 8446 3576
rect 8208 3538 8260 3544
rect 8220 2854 8248 3538
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8680 3194 8708 3334
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 8864 3058 8892 6598
rect 8956 6236 8984 6938
rect 9052 6556 9348 6576
rect 9108 6554 9132 6556
rect 9188 6554 9212 6556
rect 9268 6554 9292 6556
rect 9130 6502 9132 6554
rect 9194 6502 9206 6554
rect 9268 6502 9270 6554
rect 9108 6500 9132 6502
rect 9188 6500 9212 6502
rect 9268 6500 9292 6502
rect 9052 6480 9348 6500
rect 9036 6248 9088 6254
rect 8956 6208 9036 6236
rect 9036 6190 9088 6196
rect 9052 5468 9348 5488
rect 9108 5466 9132 5468
rect 9188 5466 9212 5468
rect 9268 5466 9292 5468
rect 9130 5414 9132 5466
rect 9194 5414 9206 5466
rect 9268 5414 9270 5466
rect 9108 5412 9132 5414
rect 9188 5412 9212 5414
rect 9268 5412 9292 5414
rect 9052 5392 9348 5412
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8956 3058 8984 5170
rect 9416 4826 9444 8434
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9600 7546 9628 7686
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9692 7274 9720 8366
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9052 4380 9348 4400
rect 9108 4378 9132 4380
rect 9188 4378 9212 4380
rect 9268 4378 9292 4380
rect 9130 4326 9132 4378
rect 9194 4326 9206 4378
rect 9268 4326 9270 4378
rect 9108 4324 9132 4326
rect 9188 4324 9212 4326
rect 9268 4324 9292 4326
rect 9052 4304 9348 4324
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9600 4078 9628 4150
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9048 3602 9076 3878
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9052 3292 9348 3312
rect 9108 3290 9132 3292
rect 9188 3290 9212 3292
rect 9268 3290 9292 3292
rect 9130 3238 9132 3290
rect 9194 3238 9206 3290
rect 9268 3238 9270 3290
rect 9108 3236 9132 3238
rect 9188 3236 9212 3238
rect 9268 3236 9292 3238
rect 9052 3216 9348 3236
rect 9508 3194 9536 3538
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 7932 2576 7984 2582
rect 7932 2518 7984 2524
rect 9508 2514 9536 3130
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 8312 800 8340 2450
rect 9052 2204 9348 2224
rect 9108 2202 9132 2204
rect 9188 2202 9212 2204
rect 9268 2202 9292 2204
rect 9130 2150 9132 2202
rect 9194 2150 9206 2202
rect 9268 2150 9270 2202
rect 9108 2148 9132 2150
rect 9188 2148 9212 2150
rect 9268 2148 9292 2150
rect 9052 2128 9348 2148
rect 9692 800 9720 6802
rect 9784 5166 9812 8434
rect 9876 8362 9904 8758
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 9876 7274 9904 7754
rect 9968 7750 9996 8978
rect 10060 8362 10088 9658
rect 10152 9586 10180 9930
rect 10244 9586 10272 10542
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10612 10198 10640 10474
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9968 7154 9996 7686
rect 10060 7478 10088 7686
rect 10152 7546 10180 9522
rect 10244 8294 10272 9522
rect 10336 9382 10364 9998
rect 10796 9518 10824 9998
rect 11072 9586 11100 10134
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 10784 9512 10836 9518
rect 10876 9512 10928 9518
rect 10784 9454 10836 9460
rect 10874 9480 10876 9489
rect 10928 9480 10930 9489
rect 11256 9466 11284 15846
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11348 14006 11376 14350
rect 11336 14000 11388 14006
rect 11336 13942 11388 13948
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11348 12986 11376 13262
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11348 12374 11376 12922
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 10874 9415 10930 9424
rect 11072 9438 11284 9466
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10336 8498 10364 9318
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10244 7954 10272 8230
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10244 7834 10272 7890
rect 10416 7880 10468 7886
rect 10244 7828 10416 7834
rect 10244 7822 10468 7828
rect 10244 7806 10456 7822
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 10060 7274 10088 7414
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 9968 7126 10088 7154
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9784 2922 9812 3470
rect 9876 2922 9904 6054
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9968 3058 9996 5510
rect 10060 4026 10088 7126
rect 10152 6662 10180 7482
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10152 6390 10180 6598
rect 10140 6384 10192 6390
rect 10140 6326 10192 6332
rect 10244 6186 10272 7806
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10336 7002 10364 7142
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10428 6254 10456 6394
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 10520 5710 10548 8570
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10612 6254 10640 6734
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10152 5370 10180 5510
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10152 4826 10180 5306
rect 10520 5166 10548 5646
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10796 4826 10824 8842
rect 11072 7426 11100 9438
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11164 7954 11192 9318
rect 11348 8974 11376 9862
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11244 8560 11296 8566
rect 11244 8502 11296 8508
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 10888 7398 11100 7426
rect 10888 6866 10916 7398
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10980 6866 11008 7278
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10980 6458 11008 6802
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 11072 6390 11100 7142
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11256 6202 11284 8502
rect 11348 7954 11376 8910
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11256 6174 11376 6202
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 10980 5658 11008 5714
rect 10980 5630 11100 5658
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10152 4146 10180 4422
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10232 4072 10284 4078
rect 10060 3998 10180 4026
rect 10232 4014 10284 4020
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 9864 2916 9916 2922
rect 9864 2858 9916 2864
rect 9784 2650 9812 2858
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 10060 2514 10088 3878
rect 10152 2922 10180 3998
rect 10244 3670 10272 4014
rect 10232 3664 10284 3670
rect 10232 3606 10284 3612
rect 10140 2916 10192 2922
rect 10140 2858 10192 2864
rect 10244 2774 10272 3606
rect 10336 3398 10364 4014
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10796 3194 10824 3946
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10152 2746 10272 2774
rect 10152 2514 10180 2746
rect 10796 2582 10824 3130
rect 10980 3058 11008 3334
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 10980 2514 11008 2994
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 11072 800 11100 5630
rect 11164 5098 11192 5714
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11164 4146 11192 5034
rect 11256 4758 11284 5102
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11164 3738 11192 3878
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11348 3670 11376 6174
rect 11440 3738 11468 8502
rect 11532 7954 11560 16390
rect 11624 15638 11652 16510
rect 11750 15804 12046 15824
rect 11806 15802 11830 15804
rect 11886 15802 11910 15804
rect 11966 15802 11990 15804
rect 11828 15750 11830 15802
rect 11892 15750 11904 15802
rect 11966 15750 11968 15802
rect 11806 15748 11830 15750
rect 11886 15748 11910 15750
rect 11966 15748 11990 15750
rect 11750 15728 12046 15748
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 12176 15570 12204 16526
rect 12452 16522 12480 17614
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12544 17338 12572 17478
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12348 16516 12400 16522
rect 12348 16458 12400 16464
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 11750 14716 12046 14736
rect 11806 14714 11830 14716
rect 11886 14714 11910 14716
rect 11966 14714 11990 14716
rect 11828 14662 11830 14714
rect 11892 14662 11904 14714
rect 11966 14662 11968 14714
rect 11806 14660 11830 14662
rect 11886 14660 11910 14662
rect 11966 14660 11990 14662
rect 11750 14640 12046 14660
rect 12360 14414 12388 16458
rect 12728 16250 12756 16594
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12716 15972 12768 15978
rect 12716 15914 12768 15920
rect 12728 15706 12756 15914
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12440 15564 12492 15570
rect 12820 15552 12848 16594
rect 12492 15524 12848 15552
rect 12440 15506 12492 15512
rect 12440 14884 12492 14890
rect 12440 14826 12492 14832
rect 12452 14618 12480 14826
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12544 14550 12572 15524
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12532 14544 12584 14550
rect 12532 14486 12584 14492
rect 12636 14482 12664 14894
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 11750 13628 12046 13648
rect 11806 13626 11830 13628
rect 11886 13626 11910 13628
rect 11966 13626 11990 13628
rect 11828 13574 11830 13626
rect 11892 13574 11904 13626
rect 11966 13574 11968 13626
rect 11806 13572 11830 13574
rect 11886 13572 11910 13574
rect 11966 13572 11990 13574
rect 11750 13552 12046 13572
rect 12360 13394 12388 14350
rect 12452 13734 12480 14418
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12636 13938 12664 14214
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12452 13462 12480 13670
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 11624 12306 11652 13330
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11808 12714 11836 13126
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 11796 12708 11848 12714
rect 11796 12650 11848 12656
rect 11750 12540 12046 12560
rect 11806 12538 11830 12540
rect 11886 12538 11910 12540
rect 11966 12538 11990 12540
rect 11828 12486 11830 12538
rect 11892 12486 11904 12538
rect 11966 12486 11968 12538
rect 11806 12484 11830 12486
rect 11886 12484 11910 12486
rect 11966 12484 11990 12486
rect 11750 12464 12046 12484
rect 12084 12306 12112 12718
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 11624 11354 11652 12242
rect 12176 11694 12204 13330
rect 12256 12776 12308 12782
rect 12256 12718 12308 12724
rect 12268 12442 12296 12718
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 12544 11898 12572 13738
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12728 12306 12756 12582
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12820 12170 12848 13262
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 11750 11452 12046 11472
rect 11806 11450 11830 11452
rect 11886 11450 11910 11452
rect 11966 11450 11990 11452
rect 11828 11398 11830 11450
rect 11892 11398 11904 11450
rect 11966 11398 11968 11450
rect 11806 11396 11830 11398
rect 11886 11396 11910 11398
rect 11966 11396 11990 11398
rect 11750 11376 12046 11396
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11624 10538 11652 11290
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 12084 10810 12112 11222
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 12176 10606 12204 11630
rect 12636 11150 12664 12038
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12820 10810 12848 11222
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 11612 10532 11664 10538
rect 11612 10474 11664 10480
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 11750 10364 12046 10384
rect 11806 10362 11830 10364
rect 11886 10362 11910 10364
rect 11966 10362 11990 10364
rect 11828 10310 11830 10362
rect 11892 10310 11904 10362
rect 11966 10310 11968 10362
rect 11806 10308 11830 10310
rect 11886 10308 11910 10310
rect 11966 10308 11990 10310
rect 11750 10288 12046 10308
rect 12452 10130 12480 10406
rect 12912 10130 12940 19804
rect 14292 17814 14320 19804
rect 15672 17882 15700 19804
rect 16394 19136 16450 19145
rect 16394 19071 16450 19080
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 14280 17808 14332 17814
rect 14280 17750 14332 17756
rect 14924 17808 14976 17814
rect 14924 17750 14976 17756
rect 14832 17740 14884 17746
rect 14832 17682 14884 17688
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 13096 16794 13124 17614
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13188 17066 13216 17478
rect 14449 17436 14745 17456
rect 14505 17434 14529 17436
rect 14585 17434 14609 17436
rect 14665 17434 14689 17436
rect 14527 17382 14529 17434
rect 14591 17382 14603 17434
rect 14665 17382 14667 17434
rect 14505 17380 14529 17382
rect 14585 17380 14609 17382
rect 14665 17380 14689 17382
rect 14449 17360 14745 17380
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 13176 17060 13228 17066
rect 13176 17002 13228 17008
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 13096 15638 13124 16730
rect 14384 16590 14412 17070
rect 14844 16998 14872 17682
rect 14832 16992 14884 16998
rect 14832 16934 14884 16940
rect 14936 16810 14964 17750
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 15028 17202 15056 17478
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15120 17066 15148 17546
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 14844 16782 14964 16810
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 13188 15570 13216 16186
rect 13464 15978 13492 16390
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 13096 14482 13124 15438
rect 13188 14822 13216 15506
rect 13280 15162 13308 15506
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 13648 15026 13676 15302
rect 13832 15094 13860 15506
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 13924 14958 13952 16050
rect 14384 15910 14412 16526
rect 14449 16348 14745 16368
rect 14505 16346 14529 16348
rect 14585 16346 14609 16348
rect 14665 16346 14689 16348
rect 14527 16294 14529 16346
rect 14591 16294 14603 16346
rect 14665 16294 14667 16346
rect 14505 16292 14529 16294
rect 14585 16292 14609 16294
rect 14665 16292 14689 16294
rect 14449 16272 14745 16292
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14384 15502 14412 15846
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13188 14618 13216 14758
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 13096 13530 13124 14418
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 13188 13462 13216 14418
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14108 14074 14136 14350
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13188 12782 13216 13126
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 13004 11762 13032 12718
rect 13188 12306 13216 12718
rect 13280 12374 13308 13330
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13268 12368 13320 12374
rect 13268 12310 13320 12316
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 13096 11694 13124 12038
rect 13280 11830 13308 12310
rect 13648 12102 13676 12786
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13740 11898 13768 12650
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13832 11830 13860 12922
rect 14108 12782 14136 14010
rect 14096 12776 14148 12782
rect 14016 12736 14096 12764
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 13832 11694 13860 11766
rect 14016 11762 14044 12736
rect 14096 12718 14148 12724
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 14108 10674 14136 12582
rect 14292 12306 14320 14418
rect 14384 13870 14412 15438
rect 14449 15260 14745 15280
rect 14505 15258 14529 15260
rect 14585 15258 14609 15260
rect 14665 15258 14689 15260
rect 14527 15206 14529 15258
rect 14591 15206 14603 15258
rect 14665 15206 14667 15258
rect 14505 15204 14529 15206
rect 14585 15204 14609 15206
rect 14665 15204 14689 15206
rect 14449 15184 14745 15204
rect 14844 15144 14872 16782
rect 15396 16590 15424 16934
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 14752 15116 14872 15144
rect 14924 15156 14976 15162
rect 14752 14346 14780 15116
rect 14924 15098 14976 15104
rect 14936 14958 14964 15098
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 14832 14544 14884 14550
rect 14832 14486 14884 14492
rect 14740 14340 14792 14346
rect 14740 14282 14792 14288
rect 14449 14172 14745 14192
rect 14505 14170 14529 14172
rect 14585 14170 14609 14172
rect 14665 14170 14689 14172
rect 14527 14118 14529 14170
rect 14591 14118 14603 14170
rect 14665 14118 14667 14170
rect 14505 14116 14529 14118
rect 14585 14116 14609 14118
rect 14665 14116 14689 14118
rect 14449 14096 14745 14116
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14292 12170 14320 12242
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14292 11694 14320 12106
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14384 11218 14412 13806
rect 14844 13258 14872 14486
rect 14936 14362 14964 14894
rect 15028 14482 15056 15914
rect 15212 15638 15240 15982
rect 15580 15638 15608 17614
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 15764 17105 15792 17478
rect 15750 17096 15806 17105
rect 15750 17031 15806 17040
rect 15200 15632 15252 15638
rect 15200 15574 15252 15580
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15120 14822 15148 14894
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 14936 14334 15056 14362
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14936 13938 14964 14214
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 15028 13530 15056 14334
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 14832 13252 14884 13258
rect 14832 13194 14884 13200
rect 14449 13084 14745 13104
rect 14505 13082 14529 13084
rect 14585 13082 14609 13084
rect 14665 13082 14689 13084
rect 14527 13030 14529 13082
rect 14591 13030 14603 13082
rect 14665 13030 14667 13082
rect 14505 13028 14529 13030
rect 14585 13028 14609 13030
rect 14665 13028 14689 13030
rect 14449 13008 14745 13028
rect 14844 12986 14872 13194
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 15120 12442 15148 14758
rect 15856 14482 15884 14758
rect 15948 14618 15976 14894
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15844 14476 15896 14482
rect 15844 14418 15896 14424
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15580 12782 15608 13262
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15396 12374 15424 12718
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15384 12368 15436 12374
rect 15384 12310 15436 12316
rect 15488 12306 15516 12650
rect 15672 12306 15700 14418
rect 15752 13456 15804 13462
rect 15752 13398 15804 13404
rect 15764 12782 15792 13398
rect 15856 13394 15884 14418
rect 15948 14074 15976 14554
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 14449 11996 14745 12016
rect 14505 11994 14529 11996
rect 14585 11994 14609 11996
rect 14665 11994 14689 11996
rect 14527 11942 14529 11994
rect 14591 11942 14603 11994
rect 14665 11942 14667 11994
rect 14505 11940 14529 11942
rect 14585 11940 14609 11942
rect 14665 11940 14689 11942
rect 14449 11920 14745 11940
rect 15120 11286 15148 12038
rect 15488 11762 15516 12242
rect 15764 11898 15792 12718
rect 15936 12368 15988 12374
rect 15936 12310 15988 12316
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15108 11280 15160 11286
rect 15108 11222 15160 11228
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14384 11082 14412 11154
rect 14372 11076 14424 11082
rect 14372 11018 14424 11024
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 13372 10130 13400 10542
rect 14384 10538 14412 11018
rect 14922 10976 14978 10985
rect 14449 10908 14745 10928
rect 14922 10911 14978 10920
rect 14505 10906 14529 10908
rect 14585 10906 14609 10908
rect 14665 10906 14689 10908
rect 14527 10854 14529 10906
rect 14591 10854 14603 10906
rect 14665 10854 14667 10906
rect 14505 10852 14529 10854
rect 14585 10852 14609 10854
rect 14665 10852 14689 10854
rect 14449 10832 14745 10852
rect 14372 10532 14424 10538
rect 14372 10474 14424 10480
rect 14832 10532 14884 10538
rect 14832 10474 14884 10480
rect 14844 10266 14872 10474
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11624 5914 11652 9318
rect 11750 9276 12046 9296
rect 11806 9274 11830 9276
rect 11886 9274 11910 9276
rect 11966 9274 11990 9276
rect 11828 9222 11830 9274
rect 11892 9222 11904 9274
rect 11966 9222 11968 9274
rect 11806 9220 11830 9222
rect 11886 9220 11910 9222
rect 11966 9220 11990 9222
rect 11750 9200 12046 9220
rect 12268 9042 12296 9590
rect 12636 9518 12664 9862
rect 13096 9586 13124 9862
rect 14449 9820 14745 9840
rect 14505 9818 14529 9820
rect 14585 9818 14609 9820
rect 14665 9818 14689 9820
rect 14527 9766 14529 9818
rect 14591 9766 14603 9818
rect 14665 9766 14667 9818
rect 14505 9764 14529 9766
rect 14585 9764 14609 9766
rect 14665 9764 14689 9766
rect 14449 9744 14745 9764
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 11750 8188 12046 8208
rect 11806 8186 11830 8188
rect 11886 8186 11910 8188
rect 11966 8186 11990 8188
rect 11828 8134 11830 8186
rect 11892 8134 11904 8186
rect 11966 8134 11968 8186
rect 11806 8132 11830 8134
rect 11886 8132 11910 8134
rect 11966 8132 11990 8134
rect 11750 8112 12046 8132
rect 12360 8090 12388 9114
rect 12728 8974 12756 9522
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 13280 9178 13308 9454
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13280 9042 13308 9114
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 13004 8498 13032 8910
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12820 8090 12848 8230
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12164 7472 12216 7478
rect 12164 7414 12216 7420
rect 11750 7100 12046 7120
rect 11806 7098 11830 7100
rect 11886 7098 11910 7100
rect 11966 7098 11990 7100
rect 11828 7046 11830 7098
rect 11892 7046 11904 7098
rect 11966 7046 11968 7098
rect 11806 7044 11830 7046
rect 11886 7044 11910 7046
rect 11966 7044 11990 7046
rect 11750 7024 12046 7044
rect 12176 6934 12204 7414
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 12268 6390 12296 7482
rect 12532 7268 12584 7274
rect 12532 7210 12584 7216
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 11750 6012 12046 6032
rect 11806 6010 11830 6012
rect 11886 6010 11910 6012
rect 11966 6010 11990 6012
rect 11828 5958 11830 6010
rect 11892 5958 11904 6010
rect 11966 5958 11968 6010
rect 11806 5956 11830 5958
rect 11886 5956 11910 5958
rect 11966 5956 11990 5958
rect 11750 5936 12046 5956
rect 12544 5914 12572 7210
rect 12728 6934 12756 7890
rect 13004 7410 13032 8434
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13188 7546 13216 7890
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 12820 7002 12848 7210
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 12256 5840 12308 5846
rect 12176 5788 12256 5794
rect 12176 5782 12308 5788
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 12176 5766 12296 5782
rect 11624 5302 11652 5714
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 11624 4690 11652 5238
rect 12084 5166 12112 5714
rect 12176 5574 12204 5766
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 11750 4924 12046 4944
rect 11806 4922 11830 4924
rect 11886 4922 11910 4924
rect 11966 4922 11990 4924
rect 11828 4870 11830 4922
rect 11892 4870 11904 4922
rect 11966 4870 11968 4922
rect 11806 4868 11830 4870
rect 11886 4868 11910 4870
rect 11966 4868 11990 4870
rect 11750 4848 12046 4868
rect 12084 4690 12112 4966
rect 12176 4826 12204 5510
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 11750 3836 12046 3856
rect 11806 3834 11830 3836
rect 11886 3834 11910 3836
rect 11966 3834 11990 3836
rect 11828 3782 11830 3834
rect 11892 3782 11904 3834
rect 11966 3782 11968 3834
rect 11806 3780 11830 3782
rect 11886 3780 11910 3782
rect 11966 3780 11990 3782
rect 11750 3760 12046 3780
rect 12452 3738 12480 3878
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11624 2582 11652 3470
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12452 2990 12480 3402
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 11750 2748 12046 2768
rect 11806 2746 11830 2748
rect 11886 2746 11910 2748
rect 11966 2746 11990 2748
rect 11828 2694 11830 2746
rect 11892 2694 11904 2746
rect 11966 2694 11968 2746
rect 11806 2692 11830 2694
rect 11886 2692 11910 2694
rect 11966 2692 11990 2694
rect 11750 2672 12046 2692
rect 12820 2582 12848 6938
rect 13188 6866 13216 7482
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 13372 5846 13400 9318
rect 13740 9110 13768 9318
rect 14752 9178 14780 9454
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13728 9104 13780 9110
rect 13728 9046 13780 9052
rect 13556 8634 13584 9046
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13740 8430 13768 9046
rect 14830 8936 14886 8945
rect 14372 8900 14424 8906
rect 14830 8871 14886 8880
rect 14372 8842 14424 8848
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13648 7002 13676 7142
rect 13740 7002 13768 7686
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13740 6254 13768 6938
rect 13924 6866 13952 8298
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 14200 6458 14228 7142
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 13096 4622 13124 5170
rect 13372 5166 13400 5782
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 12912 4214 12940 4558
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 13096 4010 13124 4558
rect 12992 4004 13044 4010
rect 12992 3946 13044 3952
rect 13084 4004 13136 4010
rect 13084 3946 13136 3952
rect 13004 3738 13032 3946
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13004 2854 13032 3470
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12452 800 12480 2450
rect 13096 2446 13124 3946
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 13188 3194 13216 3538
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13648 3058 13676 3878
rect 13740 3602 13768 4558
rect 13832 4146 13860 5714
rect 14292 5250 14320 8434
rect 14384 8090 14412 8842
rect 14449 8732 14745 8752
rect 14505 8730 14529 8732
rect 14585 8730 14609 8732
rect 14665 8730 14689 8732
rect 14527 8678 14529 8730
rect 14591 8678 14603 8730
rect 14665 8678 14667 8730
rect 14505 8676 14529 8678
rect 14585 8676 14609 8678
rect 14665 8676 14689 8678
rect 14449 8656 14745 8676
rect 14844 8430 14872 8871
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14936 7954 14964 10911
rect 15856 10418 15884 11834
rect 15948 11694 15976 12310
rect 16040 11778 16068 17682
rect 16120 17604 16172 17610
rect 16120 17546 16172 17552
rect 16132 11898 16160 17546
rect 16212 14884 16264 14890
rect 16212 14826 16264 14832
rect 16224 14618 16252 14826
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16224 12986 16252 13738
rect 16316 13530 16344 14418
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16040 11750 16160 11778
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 15948 11558 15976 11630
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15948 11354 15976 11494
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 16040 10674 16068 11630
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 15764 10390 15884 10418
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15580 9722 15608 9998
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 15028 7886 15056 8978
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14449 7644 14745 7664
rect 14505 7642 14529 7644
rect 14585 7642 14609 7644
rect 14665 7642 14689 7644
rect 14527 7590 14529 7642
rect 14591 7590 14603 7642
rect 14665 7590 14667 7642
rect 14505 7588 14529 7590
rect 14585 7588 14609 7590
rect 14665 7588 14689 7590
rect 14449 7568 14745 7588
rect 15028 7478 15056 7822
rect 15120 7546 15148 8230
rect 15212 8090 15240 9318
rect 15580 9042 15608 9658
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15304 7954 15332 8366
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15672 8022 15700 8230
rect 15660 8016 15712 8022
rect 15660 7958 15712 7964
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 15672 7342 15700 7958
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 14924 7268 14976 7274
rect 14924 7210 14976 7216
rect 14370 6896 14426 6905
rect 14370 6831 14426 6840
rect 14832 6860 14884 6866
rect 14384 6254 14412 6831
rect 14832 6802 14884 6808
rect 14449 6556 14745 6576
rect 14505 6554 14529 6556
rect 14585 6554 14609 6556
rect 14665 6554 14689 6556
rect 14527 6502 14529 6554
rect 14591 6502 14603 6554
rect 14665 6502 14667 6554
rect 14505 6500 14529 6502
rect 14585 6500 14609 6502
rect 14665 6500 14689 6502
rect 14449 6480 14745 6500
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14844 5574 14872 6802
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 14384 5370 14412 5510
rect 14449 5468 14745 5488
rect 14505 5466 14529 5468
rect 14585 5466 14609 5468
rect 14665 5466 14689 5468
rect 14527 5414 14529 5466
rect 14591 5414 14603 5466
rect 14665 5414 14667 5466
rect 14505 5412 14529 5414
rect 14585 5412 14609 5414
rect 14665 5412 14689 5414
rect 14449 5392 14745 5412
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14292 5222 14412 5250
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14188 5092 14240 5098
rect 14188 5034 14240 5040
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 14016 4690 14044 4966
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13912 4072 13964 4078
rect 13912 4014 13964 4020
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13924 3534 13952 4014
rect 14016 3670 14044 4626
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 13832 2990 13860 3334
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13924 2922 13952 3470
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 13820 2848 13872 2854
rect 14016 2802 14044 3606
rect 14200 3058 14228 5034
rect 14292 3466 14320 5102
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 14384 2825 14412 5222
rect 14832 4616 14884 4622
rect 14832 4558 14884 4564
rect 14449 4380 14745 4400
rect 14505 4378 14529 4380
rect 14585 4378 14609 4380
rect 14665 4378 14689 4380
rect 14527 4326 14529 4378
rect 14591 4326 14603 4378
rect 14665 4326 14667 4378
rect 14505 4324 14529 4326
rect 14585 4324 14609 4326
rect 14665 4324 14689 4326
rect 14449 4304 14745 4324
rect 14449 3292 14745 3312
rect 14505 3290 14529 3292
rect 14585 3290 14609 3292
rect 14665 3290 14689 3292
rect 14527 3238 14529 3290
rect 14591 3238 14603 3290
rect 14665 3238 14667 3290
rect 14505 3236 14529 3238
rect 14585 3236 14609 3238
rect 14665 3236 14689 3238
rect 14449 3216 14745 3236
rect 13872 2796 14044 2802
rect 13820 2790 14044 2796
rect 13832 2774 14044 2790
rect 14370 2816 14426 2825
rect 13924 2650 13952 2774
rect 14370 2751 14426 2760
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 14844 2582 14872 4558
rect 14936 2650 14964 7210
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15106 4856 15162 4865
rect 15106 4791 15162 4800
rect 15016 4276 15068 4282
rect 15016 4218 15068 4224
rect 15028 4146 15056 4218
rect 15016 4140 15068 4146
rect 15016 4082 15068 4088
rect 15028 3534 15056 4082
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 15028 3058 15056 3470
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 15120 2582 15148 4791
rect 14832 2576 14884 2582
rect 14832 2518 14884 2524
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13832 800 13860 2450
rect 14449 2204 14745 2224
rect 14505 2202 14529 2204
rect 14585 2202 14609 2204
rect 14665 2202 14689 2204
rect 14527 2150 14529 2202
rect 14591 2150 14603 2202
rect 14665 2150 14667 2202
rect 14505 2148 14529 2150
rect 14585 2148 14609 2150
rect 14665 2148 14689 2150
rect 14449 2128 14745 2148
rect 15212 800 15240 6802
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15304 4826 15332 6598
rect 15396 6254 15424 6666
rect 15384 6248 15436 6254
rect 15384 6190 15436 6196
rect 15396 5778 15424 6190
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15396 5166 15424 5714
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15488 5234 15516 5510
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15488 4690 15516 5170
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15304 2854 15332 3538
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15580 2774 15608 5782
rect 15764 4758 15792 10390
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15856 9110 15884 10202
rect 15936 9988 15988 9994
rect 15936 9930 15988 9936
rect 15948 9722 15976 9930
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 15856 8362 15884 9046
rect 15948 8974 15976 9454
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15844 8356 15896 8362
rect 15844 8298 15896 8304
rect 15948 8242 15976 8910
rect 15856 8214 15976 8242
rect 15856 7954 15884 8214
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15856 7002 15884 7890
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15948 5166 15976 5646
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 15948 4826 15976 5102
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 15752 4752 15804 4758
rect 15752 4694 15804 4700
rect 16132 4282 16160 11750
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16224 10266 16252 11154
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16316 10130 16344 12718
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16408 7342 16436 19071
rect 17052 17814 17080 19804
rect 17040 17808 17092 17814
rect 17040 17750 17092 17756
rect 16488 16448 16540 16454
rect 16488 16390 16540 16396
rect 16500 16182 16528 16390
rect 16488 16176 16540 16182
rect 16488 16118 16540 16124
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16592 15706 16620 15982
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 17038 15056 17094 15065
rect 17038 14991 17094 15000
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16500 13394 16528 14350
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16578 13016 16634 13025
rect 16578 12951 16634 12960
rect 16592 12306 16620 12951
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 17052 7954 17080 14991
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16224 6458 16252 6802
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16212 6248 16264 6254
rect 16212 6190 16264 6196
rect 16224 4826 16252 6190
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15672 3738 15700 4014
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15672 2990 15700 3674
rect 16408 3602 16436 3878
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 16396 2848 16448 2854
rect 16396 2790 16448 2796
rect 15580 2746 15700 2774
rect 15672 2650 15700 2746
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 16408 2582 16436 2790
rect 16396 2576 16448 2582
rect 16396 2518 16448 2524
rect 15752 2508 15804 2514
rect 15752 2450 15804 2456
rect 478 0 534 800
rect 1398 0 1454 800
rect 2778 0 2834 800
rect 4158 0 4214 800
rect 5538 0 5594 800
rect 6918 0 6974 800
rect 8298 0 8354 800
rect 9678 0 9734 800
rect 11058 0 11114 800
rect 12438 0 12494 800
rect 13818 0 13874 800
rect 15198 0 15254 800
rect 15764 785 15792 2450
rect 16580 2372 16632 2378
rect 16580 2314 16632 2320
rect 16592 800 16620 2314
rect 15750 776 15806 785
rect 15750 711 15806 720
rect 16578 0 16634 800
<< via2 >>
rect 1490 18400 1546 18456
rect 1490 10260 1546 10296
rect 1490 10240 1492 10260
rect 1492 10240 1544 10260
rect 1544 10240 1546 10260
rect 3146 16360 3202 16416
rect 2870 12280 2926 12336
rect 2226 10648 2282 10704
rect 1398 8200 1454 8256
rect 1398 4140 1454 4176
rect 1398 4120 1400 4140
rect 1400 4120 1452 4140
rect 1452 4120 1454 4140
rect 3654 17434 3710 17436
rect 3734 17434 3790 17436
rect 3814 17434 3870 17436
rect 3894 17434 3950 17436
rect 3654 17382 3680 17434
rect 3680 17382 3710 17434
rect 3734 17382 3744 17434
rect 3744 17382 3790 17434
rect 3814 17382 3860 17434
rect 3860 17382 3870 17434
rect 3894 17382 3924 17434
rect 3924 17382 3950 17434
rect 3654 17380 3710 17382
rect 3734 17380 3790 17382
rect 3814 17380 3870 17382
rect 3894 17380 3950 17382
rect 3654 16346 3710 16348
rect 3734 16346 3790 16348
rect 3814 16346 3870 16348
rect 3894 16346 3950 16348
rect 3654 16294 3680 16346
rect 3680 16294 3710 16346
rect 3734 16294 3744 16346
rect 3744 16294 3790 16346
rect 3814 16294 3860 16346
rect 3860 16294 3870 16346
rect 3894 16294 3924 16346
rect 3924 16294 3950 16346
rect 3654 16292 3710 16294
rect 3734 16292 3790 16294
rect 3814 16292 3870 16294
rect 3894 16292 3950 16294
rect 3422 14320 3478 14376
rect 3146 12300 3202 12336
rect 3146 12280 3148 12300
rect 3148 12280 3200 12300
rect 3200 12280 3202 12300
rect 3146 8916 3148 8936
rect 3148 8916 3200 8936
rect 3200 8916 3202 8936
rect 3146 8880 3202 8916
rect 3654 15258 3710 15260
rect 3734 15258 3790 15260
rect 3814 15258 3870 15260
rect 3894 15258 3950 15260
rect 3654 15206 3680 15258
rect 3680 15206 3710 15258
rect 3734 15206 3744 15258
rect 3744 15206 3790 15258
rect 3814 15206 3860 15258
rect 3860 15206 3870 15258
rect 3894 15206 3924 15258
rect 3924 15206 3950 15258
rect 3654 15204 3710 15206
rect 3734 15204 3790 15206
rect 3814 15204 3870 15206
rect 3894 15204 3950 15206
rect 3654 14170 3710 14172
rect 3734 14170 3790 14172
rect 3814 14170 3870 14172
rect 3894 14170 3950 14172
rect 3654 14118 3680 14170
rect 3680 14118 3710 14170
rect 3734 14118 3744 14170
rect 3744 14118 3790 14170
rect 3814 14118 3860 14170
rect 3860 14118 3870 14170
rect 3894 14118 3924 14170
rect 3924 14118 3950 14170
rect 3654 14116 3710 14118
rect 3734 14116 3790 14118
rect 3814 14116 3870 14118
rect 3894 14116 3950 14118
rect 3606 13776 3662 13832
rect 3654 13082 3710 13084
rect 3734 13082 3790 13084
rect 3814 13082 3870 13084
rect 3894 13082 3950 13084
rect 3654 13030 3680 13082
rect 3680 13030 3710 13082
rect 3734 13030 3744 13082
rect 3744 13030 3790 13082
rect 3814 13030 3860 13082
rect 3860 13030 3870 13082
rect 3894 13030 3924 13082
rect 3924 13030 3950 13082
rect 3654 13028 3710 13030
rect 3734 13028 3790 13030
rect 3814 13028 3870 13030
rect 3894 13028 3950 13030
rect 4342 13948 4344 13968
rect 4344 13948 4396 13968
rect 4396 13948 4398 13968
rect 4342 13912 4398 13948
rect 6353 17978 6409 17980
rect 6433 17978 6489 17980
rect 6513 17978 6569 17980
rect 6593 17978 6649 17980
rect 6353 17926 6379 17978
rect 6379 17926 6409 17978
rect 6433 17926 6443 17978
rect 6443 17926 6489 17978
rect 6513 17926 6559 17978
rect 6559 17926 6569 17978
rect 6593 17926 6623 17978
rect 6623 17926 6649 17978
rect 6353 17924 6409 17926
rect 6433 17924 6489 17926
rect 6513 17924 6569 17926
rect 6593 17924 6649 17926
rect 4894 13776 4950 13832
rect 3654 11994 3710 11996
rect 3734 11994 3790 11996
rect 3814 11994 3870 11996
rect 3894 11994 3950 11996
rect 3654 11942 3680 11994
rect 3680 11942 3710 11994
rect 3734 11942 3744 11994
rect 3744 11942 3790 11994
rect 3814 11942 3860 11994
rect 3860 11942 3870 11994
rect 3894 11942 3924 11994
rect 3924 11942 3950 11994
rect 3654 11940 3710 11942
rect 3734 11940 3790 11942
rect 3814 11940 3870 11942
rect 3894 11940 3950 11942
rect 3654 10906 3710 10908
rect 3734 10906 3790 10908
rect 3814 10906 3870 10908
rect 3894 10906 3950 10908
rect 3654 10854 3680 10906
rect 3680 10854 3710 10906
rect 3734 10854 3744 10906
rect 3744 10854 3790 10906
rect 3814 10854 3860 10906
rect 3860 10854 3870 10906
rect 3894 10854 3924 10906
rect 3924 10854 3950 10906
rect 3654 10852 3710 10854
rect 3734 10852 3790 10854
rect 3814 10852 3870 10854
rect 3894 10852 3950 10854
rect 3654 9818 3710 9820
rect 3734 9818 3790 9820
rect 3814 9818 3870 9820
rect 3894 9818 3950 9820
rect 3654 9766 3680 9818
rect 3680 9766 3710 9818
rect 3734 9766 3744 9818
rect 3744 9766 3790 9818
rect 3814 9766 3860 9818
rect 3860 9766 3870 9818
rect 3894 9766 3924 9818
rect 3924 9766 3950 9818
rect 3654 9764 3710 9766
rect 3734 9764 3790 9766
rect 3814 9764 3870 9766
rect 3894 9764 3950 9766
rect 3654 8730 3710 8732
rect 3734 8730 3790 8732
rect 3814 8730 3870 8732
rect 3894 8730 3950 8732
rect 3654 8678 3680 8730
rect 3680 8678 3710 8730
rect 3734 8678 3744 8730
rect 3744 8678 3790 8730
rect 3814 8678 3860 8730
rect 3860 8678 3870 8730
rect 3894 8678 3924 8730
rect 3924 8678 3950 8730
rect 3654 8676 3710 8678
rect 3734 8676 3790 8678
rect 3814 8676 3870 8678
rect 3894 8676 3950 8678
rect 3054 6160 3110 6216
rect 3654 7642 3710 7644
rect 3734 7642 3790 7644
rect 3814 7642 3870 7644
rect 3894 7642 3950 7644
rect 3654 7590 3680 7642
rect 3680 7590 3710 7642
rect 3734 7590 3744 7642
rect 3744 7590 3790 7642
rect 3814 7590 3860 7642
rect 3860 7590 3870 7642
rect 3894 7590 3924 7642
rect 3924 7590 3950 7642
rect 3654 7588 3710 7590
rect 3734 7588 3790 7590
rect 3814 7588 3870 7590
rect 3894 7588 3950 7590
rect 6353 16890 6409 16892
rect 6433 16890 6489 16892
rect 6513 16890 6569 16892
rect 6593 16890 6649 16892
rect 6353 16838 6379 16890
rect 6379 16838 6409 16890
rect 6433 16838 6443 16890
rect 6443 16838 6489 16890
rect 6513 16838 6559 16890
rect 6559 16838 6569 16890
rect 6593 16838 6623 16890
rect 6623 16838 6649 16890
rect 6353 16836 6409 16838
rect 6433 16836 6489 16838
rect 6513 16836 6569 16838
rect 6593 16836 6649 16838
rect 5170 13912 5226 13968
rect 4894 11736 4950 11792
rect 3654 6554 3710 6556
rect 3734 6554 3790 6556
rect 3814 6554 3870 6556
rect 3894 6554 3950 6556
rect 3654 6502 3680 6554
rect 3680 6502 3710 6554
rect 3734 6502 3744 6554
rect 3744 6502 3790 6554
rect 3814 6502 3860 6554
rect 3860 6502 3870 6554
rect 3894 6502 3924 6554
rect 3924 6502 3950 6554
rect 3654 6500 3710 6502
rect 3734 6500 3790 6502
rect 3814 6500 3870 6502
rect 3894 6500 3950 6502
rect 3654 5466 3710 5468
rect 3734 5466 3790 5468
rect 3814 5466 3870 5468
rect 3894 5466 3950 5468
rect 3654 5414 3680 5466
rect 3680 5414 3710 5466
rect 3734 5414 3744 5466
rect 3744 5414 3790 5466
rect 3814 5414 3860 5466
rect 3860 5414 3870 5466
rect 3894 5414 3924 5466
rect 3924 5414 3950 5466
rect 3654 5412 3710 5414
rect 3734 5412 3790 5414
rect 3814 5412 3870 5414
rect 3894 5412 3950 5414
rect 3654 4378 3710 4380
rect 3734 4378 3790 4380
rect 3814 4378 3870 4380
rect 3894 4378 3950 4380
rect 3654 4326 3680 4378
rect 3680 4326 3710 4378
rect 3734 4326 3744 4378
rect 3744 4326 3790 4378
rect 3814 4326 3860 4378
rect 3860 4326 3870 4378
rect 3894 4326 3924 4378
rect 3924 4326 3950 4378
rect 3654 4324 3710 4326
rect 3734 4324 3790 4326
rect 3814 4324 3870 4326
rect 3894 4324 3950 4326
rect 3330 3612 3332 3632
rect 3332 3612 3384 3632
rect 3384 3612 3386 3632
rect 3330 3576 3386 3612
rect 3654 3290 3710 3292
rect 3734 3290 3790 3292
rect 3814 3290 3870 3292
rect 3894 3290 3950 3292
rect 3654 3238 3680 3290
rect 3680 3238 3710 3290
rect 3734 3238 3744 3290
rect 3744 3238 3790 3290
rect 3814 3238 3860 3290
rect 3860 3238 3870 3290
rect 3894 3238 3924 3290
rect 3924 3238 3950 3290
rect 3654 3236 3710 3238
rect 3734 3236 3790 3238
rect 3814 3236 3870 3238
rect 3894 3236 3950 3238
rect 3654 2202 3710 2204
rect 3734 2202 3790 2204
rect 3814 2202 3870 2204
rect 3894 2202 3950 2204
rect 3654 2150 3680 2202
rect 3680 2150 3710 2202
rect 3734 2150 3744 2202
rect 3744 2150 3790 2202
rect 3814 2150 3860 2202
rect 3860 2150 3870 2202
rect 3894 2150 3924 2202
rect 3924 2150 3950 2202
rect 3654 2148 3710 2150
rect 3734 2148 3790 2150
rect 3814 2148 3870 2150
rect 3894 2148 3950 2150
rect 2870 2080 2926 2136
rect 5998 15564 6054 15600
rect 5998 15544 6000 15564
rect 6000 15544 6052 15564
rect 6052 15544 6054 15564
rect 6353 15802 6409 15804
rect 6433 15802 6489 15804
rect 6513 15802 6569 15804
rect 6593 15802 6649 15804
rect 6353 15750 6379 15802
rect 6379 15750 6409 15802
rect 6433 15750 6443 15802
rect 6443 15750 6489 15802
rect 6513 15750 6559 15802
rect 6559 15750 6569 15802
rect 6593 15750 6623 15802
rect 6623 15750 6649 15802
rect 6353 15748 6409 15750
rect 6433 15748 6489 15750
rect 6513 15748 6569 15750
rect 6593 15748 6649 15750
rect 7286 15544 7342 15600
rect 5998 13812 6000 13832
rect 6000 13812 6052 13832
rect 6052 13812 6054 13832
rect 5998 13776 6054 13812
rect 5814 12280 5870 12336
rect 5814 11872 5870 11928
rect 6353 14714 6409 14716
rect 6433 14714 6489 14716
rect 6513 14714 6569 14716
rect 6593 14714 6649 14716
rect 6353 14662 6379 14714
rect 6379 14662 6409 14714
rect 6433 14662 6443 14714
rect 6443 14662 6489 14714
rect 6513 14662 6559 14714
rect 6559 14662 6569 14714
rect 6593 14662 6623 14714
rect 6623 14662 6649 14714
rect 6353 14660 6409 14662
rect 6433 14660 6489 14662
rect 6513 14660 6569 14662
rect 6593 14660 6649 14662
rect 6353 13626 6409 13628
rect 6433 13626 6489 13628
rect 6513 13626 6569 13628
rect 6593 13626 6649 13628
rect 6353 13574 6379 13626
rect 6379 13574 6409 13626
rect 6433 13574 6443 13626
rect 6443 13574 6489 13626
rect 6513 13574 6559 13626
rect 6559 13574 6569 13626
rect 6593 13574 6623 13626
rect 6623 13574 6649 13626
rect 6353 13572 6409 13574
rect 6433 13572 6489 13574
rect 6513 13572 6569 13574
rect 6593 13572 6649 13574
rect 6353 12538 6409 12540
rect 6433 12538 6489 12540
rect 6513 12538 6569 12540
rect 6593 12538 6649 12540
rect 6353 12486 6379 12538
rect 6379 12486 6409 12538
rect 6433 12486 6443 12538
rect 6443 12486 6489 12538
rect 6513 12486 6559 12538
rect 6559 12486 6569 12538
rect 6593 12486 6623 12538
rect 6623 12486 6649 12538
rect 6353 12484 6409 12486
rect 6433 12484 6489 12486
rect 6513 12484 6569 12486
rect 6593 12484 6649 12486
rect 6550 12300 6606 12336
rect 6550 12280 6552 12300
rect 6552 12280 6604 12300
rect 6604 12280 6606 12300
rect 6550 12164 6606 12200
rect 6550 12144 6552 12164
rect 6552 12144 6604 12164
rect 6604 12144 6606 12164
rect 4618 5772 4674 5808
rect 4618 5752 4620 5772
rect 4620 5752 4672 5772
rect 4672 5752 4674 5772
rect 5814 3440 5870 3496
rect 7010 12144 7066 12200
rect 7010 11872 7066 11928
rect 6734 11736 6790 11792
rect 6353 11450 6409 11452
rect 6433 11450 6489 11452
rect 6513 11450 6569 11452
rect 6593 11450 6649 11452
rect 6353 11398 6379 11450
rect 6379 11398 6409 11450
rect 6433 11398 6443 11450
rect 6443 11398 6489 11450
rect 6513 11398 6559 11450
rect 6559 11398 6569 11450
rect 6593 11398 6623 11450
rect 6623 11398 6649 11450
rect 6353 11396 6409 11398
rect 6433 11396 6489 11398
rect 6513 11396 6569 11398
rect 6593 11396 6649 11398
rect 6353 10362 6409 10364
rect 6433 10362 6489 10364
rect 6513 10362 6569 10364
rect 6593 10362 6649 10364
rect 6353 10310 6379 10362
rect 6379 10310 6409 10362
rect 6433 10310 6443 10362
rect 6443 10310 6489 10362
rect 6513 10310 6559 10362
rect 6559 10310 6569 10362
rect 6593 10310 6623 10362
rect 6623 10310 6649 10362
rect 6353 10308 6409 10310
rect 6433 10308 6489 10310
rect 6513 10308 6569 10310
rect 6593 10308 6649 10310
rect 6353 9274 6409 9276
rect 6433 9274 6489 9276
rect 6513 9274 6569 9276
rect 6593 9274 6649 9276
rect 6353 9222 6379 9274
rect 6379 9222 6409 9274
rect 6433 9222 6443 9274
rect 6443 9222 6489 9274
rect 6513 9222 6559 9274
rect 6559 9222 6569 9274
rect 6593 9222 6623 9274
rect 6623 9222 6649 9274
rect 6353 9220 6409 9222
rect 6433 9220 6489 9222
rect 6513 9220 6569 9222
rect 6593 9220 6649 9222
rect 7010 9288 7066 9344
rect 6353 8186 6409 8188
rect 6433 8186 6489 8188
rect 6513 8186 6569 8188
rect 6593 8186 6649 8188
rect 6353 8134 6379 8186
rect 6379 8134 6409 8186
rect 6433 8134 6443 8186
rect 6443 8134 6489 8186
rect 6513 8134 6559 8186
rect 6559 8134 6569 8186
rect 6593 8134 6623 8186
rect 6623 8134 6649 8186
rect 6353 8132 6409 8134
rect 6433 8132 6489 8134
rect 6513 8132 6569 8134
rect 6593 8132 6649 8134
rect 6353 7098 6409 7100
rect 6433 7098 6489 7100
rect 6513 7098 6569 7100
rect 6593 7098 6649 7100
rect 6353 7046 6379 7098
rect 6379 7046 6409 7098
rect 6433 7046 6443 7098
rect 6443 7046 6489 7098
rect 6513 7046 6559 7098
rect 6559 7046 6569 7098
rect 6593 7046 6623 7098
rect 6623 7046 6649 7098
rect 6353 7044 6409 7046
rect 6433 7044 6489 7046
rect 6513 7044 6569 7046
rect 6593 7044 6649 7046
rect 6353 6010 6409 6012
rect 6433 6010 6489 6012
rect 6513 6010 6569 6012
rect 6593 6010 6649 6012
rect 6353 5958 6379 6010
rect 6379 5958 6409 6010
rect 6433 5958 6443 6010
rect 6443 5958 6489 6010
rect 6513 5958 6559 6010
rect 6559 5958 6569 6010
rect 6593 5958 6623 6010
rect 6623 5958 6649 6010
rect 6353 5956 6409 5958
rect 6433 5956 6489 5958
rect 6513 5956 6569 5958
rect 6593 5956 6649 5958
rect 6353 4922 6409 4924
rect 6433 4922 6489 4924
rect 6513 4922 6569 4924
rect 6593 4922 6649 4924
rect 6353 4870 6379 4922
rect 6379 4870 6409 4922
rect 6433 4870 6443 4922
rect 6443 4870 6489 4922
rect 6513 4870 6559 4922
rect 6559 4870 6569 4922
rect 6593 4870 6623 4922
rect 6623 4870 6649 4922
rect 6353 4868 6409 4870
rect 6433 4868 6489 4870
rect 6513 4868 6569 4870
rect 6593 4868 6649 4870
rect 6353 3834 6409 3836
rect 6433 3834 6489 3836
rect 6513 3834 6569 3836
rect 6593 3834 6649 3836
rect 6353 3782 6379 3834
rect 6379 3782 6409 3834
rect 6433 3782 6443 3834
rect 6443 3782 6489 3834
rect 6513 3782 6559 3834
rect 6559 3782 6569 3834
rect 6593 3782 6623 3834
rect 6623 3782 6649 3834
rect 6353 3780 6409 3782
rect 6433 3780 6489 3782
rect 6513 3780 6569 3782
rect 6593 3780 6649 3782
rect 9052 17434 9108 17436
rect 9132 17434 9188 17436
rect 9212 17434 9268 17436
rect 9292 17434 9348 17436
rect 9052 17382 9078 17434
rect 9078 17382 9108 17434
rect 9132 17382 9142 17434
rect 9142 17382 9188 17434
rect 9212 17382 9258 17434
rect 9258 17382 9268 17434
rect 9292 17382 9322 17434
rect 9322 17382 9348 17434
rect 9052 17380 9108 17382
rect 9132 17380 9188 17382
rect 9212 17380 9268 17382
rect 9292 17380 9348 17382
rect 9052 16346 9108 16348
rect 9132 16346 9188 16348
rect 9212 16346 9268 16348
rect 9292 16346 9348 16348
rect 9052 16294 9078 16346
rect 9078 16294 9108 16346
rect 9132 16294 9142 16346
rect 9142 16294 9188 16346
rect 9212 16294 9258 16346
rect 9258 16294 9268 16346
rect 9292 16294 9322 16346
rect 9322 16294 9348 16346
rect 9052 16292 9108 16294
rect 9132 16292 9188 16294
rect 9212 16292 9268 16294
rect 9292 16292 9348 16294
rect 9052 15258 9108 15260
rect 9132 15258 9188 15260
rect 9212 15258 9268 15260
rect 9292 15258 9348 15260
rect 9052 15206 9078 15258
rect 9078 15206 9108 15258
rect 9132 15206 9142 15258
rect 9142 15206 9188 15258
rect 9212 15206 9258 15258
rect 9258 15206 9268 15258
rect 9292 15206 9322 15258
rect 9322 15206 9348 15258
rect 9052 15204 9108 15206
rect 9132 15204 9188 15206
rect 9212 15204 9268 15206
rect 9292 15204 9348 15206
rect 9052 14170 9108 14172
rect 9132 14170 9188 14172
rect 9212 14170 9268 14172
rect 9292 14170 9348 14172
rect 9052 14118 9078 14170
rect 9078 14118 9108 14170
rect 9132 14118 9142 14170
rect 9142 14118 9188 14170
rect 9212 14118 9258 14170
rect 9258 14118 9268 14170
rect 9292 14118 9322 14170
rect 9322 14118 9348 14170
rect 9052 14116 9108 14118
rect 9132 14116 9188 14118
rect 9212 14116 9268 14118
rect 9292 14116 9348 14118
rect 11750 17978 11806 17980
rect 11830 17978 11886 17980
rect 11910 17978 11966 17980
rect 11990 17978 12046 17980
rect 11750 17926 11776 17978
rect 11776 17926 11806 17978
rect 11830 17926 11840 17978
rect 11840 17926 11886 17978
rect 11910 17926 11956 17978
rect 11956 17926 11966 17978
rect 11990 17926 12020 17978
rect 12020 17926 12046 17978
rect 11750 17924 11806 17926
rect 11830 17924 11886 17926
rect 11910 17924 11966 17926
rect 11990 17924 12046 17926
rect 11750 16890 11806 16892
rect 11830 16890 11886 16892
rect 11910 16890 11966 16892
rect 11990 16890 12046 16892
rect 11750 16838 11776 16890
rect 11776 16838 11806 16890
rect 11830 16838 11840 16890
rect 11840 16838 11886 16890
rect 11910 16838 11956 16890
rect 11956 16838 11966 16890
rect 11990 16838 12020 16890
rect 12020 16838 12046 16890
rect 11750 16836 11806 16838
rect 11830 16836 11886 16838
rect 11910 16836 11966 16838
rect 11990 16836 12046 16838
rect 9052 13082 9108 13084
rect 9132 13082 9188 13084
rect 9212 13082 9268 13084
rect 9292 13082 9348 13084
rect 9052 13030 9078 13082
rect 9078 13030 9108 13082
rect 9132 13030 9142 13082
rect 9142 13030 9188 13082
rect 9212 13030 9258 13082
rect 9258 13030 9268 13082
rect 9292 13030 9322 13082
rect 9322 13030 9348 13082
rect 9052 13028 9108 13030
rect 9132 13028 9188 13030
rect 9212 13028 9268 13030
rect 9292 13028 9348 13030
rect 9052 11994 9108 11996
rect 9132 11994 9188 11996
rect 9212 11994 9268 11996
rect 9292 11994 9348 11996
rect 9052 11942 9078 11994
rect 9078 11942 9108 11994
rect 9132 11942 9142 11994
rect 9142 11942 9188 11994
rect 9212 11942 9258 11994
rect 9258 11942 9268 11994
rect 9292 11942 9322 11994
rect 9322 11942 9348 11994
rect 9052 11940 9108 11942
rect 9132 11940 9188 11942
rect 9212 11940 9268 11942
rect 9292 11940 9348 11942
rect 9052 10906 9108 10908
rect 9132 10906 9188 10908
rect 9212 10906 9268 10908
rect 9292 10906 9348 10908
rect 9052 10854 9078 10906
rect 9078 10854 9108 10906
rect 9132 10854 9142 10906
rect 9142 10854 9188 10906
rect 9212 10854 9258 10906
rect 9258 10854 9268 10906
rect 9292 10854 9322 10906
rect 9322 10854 9348 10906
rect 9052 10852 9108 10854
rect 9132 10852 9188 10854
rect 9212 10852 9268 10854
rect 9292 10852 9348 10854
rect 8666 10668 8722 10704
rect 8666 10648 8668 10668
rect 8668 10648 8720 10668
rect 8720 10648 8722 10668
rect 7930 9460 7932 9480
rect 7932 9460 7984 9480
rect 7984 9460 7986 9480
rect 7930 9424 7986 9460
rect 8482 8916 8484 8936
rect 8484 8916 8536 8936
rect 8536 8916 8538 8936
rect 8482 8880 8538 8916
rect 7654 5752 7710 5808
rect 9052 9818 9108 9820
rect 9132 9818 9188 9820
rect 9212 9818 9268 9820
rect 9292 9818 9348 9820
rect 9052 9766 9078 9818
rect 9078 9766 9108 9818
rect 9132 9766 9142 9818
rect 9142 9766 9188 9818
rect 9212 9766 9258 9818
rect 9258 9766 9268 9818
rect 9292 9766 9322 9818
rect 9322 9766 9348 9818
rect 9052 9764 9108 9766
rect 9132 9764 9188 9766
rect 9212 9764 9268 9766
rect 9292 9764 9348 9766
rect 9034 9324 9036 9344
rect 9036 9324 9088 9344
rect 9088 9324 9090 9344
rect 9034 9288 9090 9324
rect 9052 8730 9108 8732
rect 9132 8730 9188 8732
rect 9212 8730 9268 8732
rect 9292 8730 9348 8732
rect 9052 8678 9078 8730
rect 9078 8678 9108 8730
rect 9132 8678 9142 8730
rect 9142 8678 9188 8730
rect 9212 8678 9258 8730
rect 9258 8678 9268 8730
rect 9292 8678 9322 8730
rect 9322 8678 9348 8730
rect 9052 8676 9108 8678
rect 9132 8676 9188 8678
rect 9212 8676 9268 8678
rect 9292 8676 9348 8678
rect 9052 7642 9108 7644
rect 9132 7642 9188 7644
rect 9212 7642 9268 7644
rect 9292 7642 9348 7644
rect 9052 7590 9078 7642
rect 9078 7590 9108 7642
rect 9132 7590 9142 7642
rect 9142 7590 9188 7642
rect 9212 7590 9258 7642
rect 9258 7590 9268 7642
rect 9292 7590 9322 7642
rect 9322 7590 9348 7642
rect 9052 7588 9108 7590
rect 9132 7588 9188 7590
rect 9212 7588 9268 7590
rect 9292 7588 9348 7590
rect 6918 3712 6974 3768
rect 6366 3476 6368 3496
rect 6368 3476 6420 3496
rect 6420 3476 6422 3496
rect 6366 3440 6422 3476
rect 6353 2746 6409 2748
rect 6433 2746 6489 2748
rect 6513 2746 6569 2748
rect 6593 2746 6649 2748
rect 6353 2694 6379 2746
rect 6379 2694 6409 2746
rect 6433 2694 6443 2746
rect 6443 2694 6489 2746
rect 6513 2694 6559 2746
rect 6559 2694 6569 2746
rect 6593 2694 6623 2746
rect 6623 2694 6649 2746
rect 6353 2692 6409 2694
rect 6433 2692 6489 2694
rect 6513 2692 6569 2694
rect 6593 2692 6649 2694
rect 8758 3712 8814 3768
rect 8390 3612 8392 3632
rect 8392 3612 8444 3632
rect 8444 3612 8446 3632
rect 8390 3576 8446 3612
rect 9052 6554 9108 6556
rect 9132 6554 9188 6556
rect 9212 6554 9268 6556
rect 9292 6554 9348 6556
rect 9052 6502 9078 6554
rect 9078 6502 9108 6554
rect 9132 6502 9142 6554
rect 9142 6502 9188 6554
rect 9212 6502 9258 6554
rect 9258 6502 9268 6554
rect 9292 6502 9322 6554
rect 9322 6502 9348 6554
rect 9052 6500 9108 6502
rect 9132 6500 9188 6502
rect 9212 6500 9268 6502
rect 9292 6500 9348 6502
rect 9052 5466 9108 5468
rect 9132 5466 9188 5468
rect 9212 5466 9268 5468
rect 9292 5466 9348 5468
rect 9052 5414 9078 5466
rect 9078 5414 9108 5466
rect 9132 5414 9142 5466
rect 9142 5414 9188 5466
rect 9212 5414 9258 5466
rect 9258 5414 9268 5466
rect 9292 5414 9322 5466
rect 9322 5414 9348 5466
rect 9052 5412 9108 5414
rect 9132 5412 9188 5414
rect 9212 5412 9268 5414
rect 9292 5412 9348 5414
rect 9052 4378 9108 4380
rect 9132 4378 9188 4380
rect 9212 4378 9268 4380
rect 9292 4378 9348 4380
rect 9052 4326 9078 4378
rect 9078 4326 9108 4378
rect 9132 4326 9142 4378
rect 9142 4326 9188 4378
rect 9212 4326 9258 4378
rect 9258 4326 9268 4378
rect 9292 4326 9322 4378
rect 9322 4326 9348 4378
rect 9052 4324 9108 4326
rect 9132 4324 9188 4326
rect 9212 4324 9268 4326
rect 9292 4324 9348 4326
rect 9052 3290 9108 3292
rect 9132 3290 9188 3292
rect 9212 3290 9268 3292
rect 9292 3290 9348 3292
rect 9052 3238 9078 3290
rect 9078 3238 9108 3290
rect 9132 3238 9142 3290
rect 9142 3238 9188 3290
rect 9212 3238 9258 3290
rect 9258 3238 9268 3290
rect 9292 3238 9322 3290
rect 9322 3238 9348 3290
rect 9052 3236 9108 3238
rect 9132 3236 9188 3238
rect 9212 3236 9268 3238
rect 9292 3236 9348 3238
rect 9052 2202 9108 2204
rect 9132 2202 9188 2204
rect 9212 2202 9268 2204
rect 9292 2202 9348 2204
rect 9052 2150 9078 2202
rect 9078 2150 9108 2202
rect 9132 2150 9142 2202
rect 9142 2150 9188 2202
rect 9212 2150 9258 2202
rect 9258 2150 9268 2202
rect 9292 2150 9322 2202
rect 9322 2150 9348 2202
rect 9052 2148 9108 2150
rect 9132 2148 9188 2150
rect 9212 2148 9268 2150
rect 9292 2148 9348 2150
rect 10874 9460 10876 9480
rect 10876 9460 10928 9480
rect 10928 9460 10930 9480
rect 10874 9424 10930 9460
rect 11750 15802 11806 15804
rect 11830 15802 11886 15804
rect 11910 15802 11966 15804
rect 11990 15802 12046 15804
rect 11750 15750 11776 15802
rect 11776 15750 11806 15802
rect 11830 15750 11840 15802
rect 11840 15750 11886 15802
rect 11910 15750 11956 15802
rect 11956 15750 11966 15802
rect 11990 15750 12020 15802
rect 12020 15750 12046 15802
rect 11750 15748 11806 15750
rect 11830 15748 11886 15750
rect 11910 15748 11966 15750
rect 11990 15748 12046 15750
rect 11750 14714 11806 14716
rect 11830 14714 11886 14716
rect 11910 14714 11966 14716
rect 11990 14714 12046 14716
rect 11750 14662 11776 14714
rect 11776 14662 11806 14714
rect 11830 14662 11840 14714
rect 11840 14662 11886 14714
rect 11910 14662 11956 14714
rect 11956 14662 11966 14714
rect 11990 14662 12020 14714
rect 12020 14662 12046 14714
rect 11750 14660 11806 14662
rect 11830 14660 11886 14662
rect 11910 14660 11966 14662
rect 11990 14660 12046 14662
rect 11750 13626 11806 13628
rect 11830 13626 11886 13628
rect 11910 13626 11966 13628
rect 11990 13626 12046 13628
rect 11750 13574 11776 13626
rect 11776 13574 11806 13626
rect 11830 13574 11840 13626
rect 11840 13574 11886 13626
rect 11910 13574 11956 13626
rect 11956 13574 11966 13626
rect 11990 13574 12020 13626
rect 12020 13574 12046 13626
rect 11750 13572 11806 13574
rect 11830 13572 11886 13574
rect 11910 13572 11966 13574
rect 11990 13572 12046 13574
rect 11750 12538 11806 12540
rect 11830 12538 11886 12540
rect 11910 12538 11966 12540
rect 11990 12538 12046 12540
rect 11750 12486 11776 12538
rect 11776 12486 11806 12538
rect 11830 12486 11840 12538
rect 11840 12486 11886 12538
rect 11910 12486 11956 12538
rect 11956 12486 11966 12538
rect 11990 12486 12020 12538
rect 12020 12486 12046 12538
rect 11750 12484 11806 12486
rect 11830 12484 11886 12486
rect 11910 12484 11966 12486
rect 11990 12484 12046 12486
rect 11750 11450 11806 11452
rect 11830 11450 11886 11452
rect 11910 11450 11966 11452
rect 11990 11450 12046 11452
rect 11750 11398 11776 11450
rect 11776 11398 11806 11450
rect 11830 11398 11840 11450
rect 11840 11398 11886 11450
rect 11910 11398 11956 11450
rect 11956 11398 11966 11450
rect 11990 11398 12020 11450
rect 12020 11398 12046 11450
rect 11750 11396 11806 11398
rect 11830 11396 11886 11398
rect 11910 11396 11966 11398
rect 11990 11396 12046 11398
rect 11750 10362 11806 10364
rect 11830 10362 11886 10364
rect 11910 10362 11966 10364
rect 11990 10362 12046 10364
rect 11750 10310 11776 10362
rect 11776 10310 11806 10362
rect 11830 10310 11840 10362
rect 11840 10310 11886 10362
rect 11910 10310 11956 10362
rect 11956 10310 11966 10362
rect 11990 10310 12020 10362
rect 12020 10310 12046 10362
rect 11750 10308 11806 10310
rect 11830 10308 11886 10310
rect 11910 10308 11966 10310
rect 11990 10308 12046 10310
rect 16394 19080 16450 19136
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14609 17434 14665 17436
rect 14689 17434 14745 17436
rect 14449 17382 14475 17434
rect 14475 17382 14505 17434
rect 14529 17382 14539 17434
rect 14539 17382 14585 17434
rect 14609 17382 14655 17434
rect 14655 17382 14665 17434
rect 14689 17382 14719 17434
rect 14719 17382 14745 17434
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14609 17380 14665 17382
rect 14689 17380 14745 17382
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14609 16346 14665 16348
rect 14689 16346 14745 16348
rect 14449 16294 14475 16346
rect 14475 16294 14505 16346
rect 14529 16294 14539 16346
rect 14539 16294 14585 16346
rect 14609 16294 14655 16346
rect 14655 16294 14665 16346
rect 14689 16294 14719 16346
rect 14719 16294 14745 16346
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14609 16292 14665 16294
rect 14689 16292 14745 16294
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14609 15258 14665 15260
rect 14689 15258 14745 15260
rect 14449 15206 14475 15258
rect 14475 15206 14505 15258
rect 14529 15206 14539 15258
rect 14539 15206 14585 15258
rect 14609 15206 14655 15258
rect 14655 15206 14665 15258
rect 14689 15206 14719 15258
rect 14719 15206 14745 15258
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 14609 15204 14665 15206
rect 14689 15204 14745 15206
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14609 14170 14665 14172
rect 14689 14170 14745 14172
rect 14449 14118 14475 14170
rect 14475 14118 14505 14170
rect 14529 14118 14539 14170
rect 14539 14118 14585 14170
rect 14609 14118 14655 14170
rect 14655 14118 14665 14170
rect 14689 14118 14719 14170
rect 14719 14118 14745 14170
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14609 14116 14665 14118
rect 14689 14116 14745 14118
rect 15750 17040 15806 17096
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14609 13082 14665 13084
rect 14689 13082 14745 13084
rect 14449 13030 14475 13082
rect 14475 13030 14505 13082
rect 14529 13030 14539 13082
rect 14539 13030 14585 13082
rect 14609 13030 14655 13082
rect 14655 13030 14665 13082
rect 14689 13030 14719 13082
rect 14719 13030 14745 13082
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14609 13028 14665 13030
rect 14689 13028 14745 13030
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14609 11994 14665 11996
rect 14689 11994 14745 11996
rect 14449 11942 14475 11994
rect 14475 11942 14505 11994
rect 14529 11942 14539 11994
rect 14539 11942 14585 11994
rect 14609 11942 14655 11994
rect 14655 11942 14665 11994
rect 14689 11942 14719 11994
rect 14719 11942 14745 11994
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14609 11940 14665 11942
rect 14689 11940 14745 11942
rect 14922 10920 14978 10976
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14609 10906 14665 10908
rect 14689 10906 14745 10908
rect 14449 10854 14475 10906
rect 14475 10854 14505 10906
rect 14529 10854 14539 10906
rect 14539 10854 14585 10906
rect 14609 10854 14655 10906
rect 14655 10854 14665 10906
rect 14689 10854 14719 10906
rect 14719 10854 14745 10906
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14609 10852 14665 10854
rect 14689 10852 14745 10854
rect 11750 9274 11806 9276
rect 11830 9274 11886 9276
rect 11910 9274 11966 9276
rect 11990 9274 12046 9276
rect 11750 9222 11776 9274
rect 11776 9222 11806 9274
rect 11830 9222 11840 9274
rect 11840 9222 11886 9274
rect 11910 9222 11956 9274
rect 11956 9222 11966 9274
rect 11990 9222 12020 9274
rect 12020 9222 12046 9274
rect 11750 9220 11806 9222
rect 11830 9220 11886 9222
rect 11910 9220 11966 9222
rect 11990 9220 12046 9222
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14609 9818 14665 9820
rect 14689 9818 14745 9820
rect 14449 9766 14475 9818
rect 14475 9766 14505 9818
rect 14529 9766 14539 9818
rect 14539 9766 14585 9818
rect 14609 9766 14655 9818
rect 14655 9766 14665 9818
rect 14689 9766 14719 9818
rect 14719 9766 14745 9818
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14609 9764 14665 9766
rect 14689 9764 14745 9766
rect 11750 8186 11806 8188
rect 11830 8186 11886 8188
rect 11910 8186 11966 8188
rect 11990 8186 12046 8188
rect 11750 8134 11776 8186
rect 11776 8134 11806 8186
rect 11830 8134 11840 8186
rect 11840 8134 11886 8186
rect 11910 8134 11956 8186
rect 11956 8134 11966 8186
rect 11990 8134 12020 8186
rect 12020 8134 12046 8186
rect 11750 8132 11806 8134
rect 11830 8132 11886 8134
rect 11910 8132 11966 8134
rect 11990 8132 12046 8134
rect 11750 7098 11806 7100
rect 11830 7098 11886 7100
rect 11910 7098 11966 7100
rect 11990 7098 12046 7100
rect 11750 7046 11776 7098
rect 11776 7046 11806 7098
rect 11830 7046 11840 7098
rect 11840 7046 11886 7098
rect 11910 7046 11956 7098
rect 11956 7046 11966 7098
rect 11990 7046 12020 7098
rect 12020 7046 12046 7098
rect 11750 7044 11806 7046
rect 11830 7044 11886 7046
rect 11910 7044 11966 7046
rect 11990 7044 12046 7046
rect 11750 6010 11806 6012
rect 11830 6010 11886 6012
rect 11910 6010 11966 6012
rect 11990 6010 12046 6012
rect 11750 5958 11776 6010
rect 11776 5958 11806 6010
rect 11830 5958 11840 6010
rect 11840 5958 11886 6010
rect 11910 5958 11956 6010
rect 11956 5958 11966 6010
rect 11990 5958 12020 6010
rect 12020 5958 12046 6010
rect 11750 5956 11806 5958
rect 11830 5956 11886 5958
rect 11910 5956 11966 5958
rect 11990 5956 12046 5958
rect 11750 4922 11806 4924
rect 11830 4922 11886 4924
rect 11910 4922 11966 4924
rect 11990 4922 12046 4924
rect 11750 4870 11776 4922
rect 11776 4870 11806 4922
rect 11830 4870 11840 4922
rect 11840 4870 11886 4922
rect 11910 4870 11956 4922
rect 11956 4870 11966 4922
rect 11990 4870 12020 4922
rect 12020 4870 12046 4922
rect 11750 4868 11806 4870
rect 11830 4868 11886 4870
rect 11910 4868 11966 4870
rect 11990 4868 12046 4870
rect 11750 3834 11806 3836
rect 11830 3834 11886 3836
rect 11910 3834 11966 3836
rect 11990 3834 12046 3836
rect 11750 3782 11776 3834
rect 11776 3782 11806 3834
rect 11830 3782 11840 3834
rect 11840 3782 11886 3834
rect 11910 3782 11956 3834
rect 11956 3782 11966 3834
rect 11990 3782 12020 3834
rect 12020 3782 12046 3834
rect 11750 3780 11806 3782
rect 11830 3780 11886 3782
rect 11910 3780 11966 3782
rect 11990 3780 12046 3782
rect 11750 2746 11806 2748
rect 11830 2746 11886 2748
rect 11910 2746 11966 2748
rect 11990 2746 12046 2748
rect 11750 2694 11776 2746
rect 11776 2694 11806 2746
rect 11830 2694 11840 2746
rect 11840 2694 11886 2746
rect 11910 2694 11956 2746
rect 11956 2694 11966 2746
rect 11990 2694 12020 2746
rect 12020 2694 12046 2746
rect 11750 2692 11806 2694
rect 11830 2692 11886 2694
rect 11910 2692 11966 2694
rect 11990 2692 12046 2694
rect 14830 8880 14886 8936
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14609 8730 14665 8732
rect 14689 8730 14745 8732
rect 14449 8678 14475 8730
rect 14475 8678 14505 8730
rect 14529 8678 14539 8730
rect 14539 8678 14585 8730
rect 14609 8678 14655 8730
rect 14655 8678 14665 8730
rect 14689 8678 14719 8730
rect 14719 8678 14745 8730
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14609 8676 14665 8678
rect 14689 8676 14745 8678
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14609 7642 14665 7644
rect 14689 7642 14745 7644
rect 14449 7590 14475 7642
rect 14475 7590 14505 7642
rect 14529 7590 14539 7642
rect 14539 7590 14585 7642
rect 14609 7590 14655 7642
rect 14655 7590 14665 7642
rect 14689 7590 14719 7642
rect 14719 7590 14745 7642
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14609 7588 14665 7590
rect 14689 7588 14745 7590
rect 14370 6840 14426 6896
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14609 6554 14665 6556
rect 14689 6554 14745 6556
rect 14449 6502 14475 6554
rect 14475 6502 14505 6554
rect 14529 6502 14539 6554
rect 14539 6502 14585 6554
rect 14609 6502 14655 6554
rect 14655 6502 14665 6554
rect 14689 6502 14719 6554
rect 14719 6502 14745 6554
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14609 6500 14665 6502
rect 14689 6500 14745 6502
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14609 5466 14665 5468
rect 14689 5466 14745 5468
rect 14449 5414 14475 5466
rect 14475 5414 14505 5466
rect 14529 5414 14539 5466
rect 14539 5414 14585 5466
rect 14609 5414 14655 5466
rect 14655 5414 14665 5466
rect 14689 5414 14719 5466
rect 14719 5414 14745 5466
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 14609 5412 14665 5414
rect 14689 5412 14745 5414
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14609 4378 14665 4380
rect 14689 4378 14745 4380
rect 14449 4326 14475 4378
rect 14475 4326 14505 4378
rect 14529 4326 14539 4378
rect 14539 4326 14585 4378
rect 14609 4326 14655 4378
rect 14655 4326 14665 4378
rect 14689 4326 14719 4378
rect 14719 4326 14745 4378
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14609 4324 14665 4326
rect 14689 4324 14745 4326
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14609 3290 14665 3292
rect 14689 3290 14745 3292
rect 14449 3238 14475 3290
rect 14475 3238 14505 3290
rect 14529 3238 14539 3290
rect 14539 3238 14585 3290
rect 14609 3238 14655 3290
rect 14655 3238 14665 3290
rect 14689 3238 14719 3290
rect 14719 3238 14745 3290
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14609 3236 14665 3238
rect 14689 3236 14745 3238
rect 14370 2760 14426 2816
rect 15106 4800 15162 4856
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14609 2202 14665 2204
rect 14689 2202 14745 2204
rect 14449 2150 14475 2202
rect 14475 2150 14505 2202
rect 14529 2150 14539 2202
rect 14539 2150 14585 2202
rect 14609 2150 14655 2202
rect 14655 2150 14665 2202
rect 14689 2150 14719 2202
rect 14719 2150 14745 2202
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
rect 14609 2148 14665 2150
rect 14689 2148 14745 2150
rect 17038 15000 17094 15056
rect 16578 12960 16634 13016
rect 15750 720 15806 776
<< metal3 >>
rect 16389 19138 16455 19141
rect 17660 19138 18460 19168
rect 16389 19136 18460 19138
rect 16389 19080 16394 19136
rect 16450 19080 18460 19136
rect 16389 19078 18460 19080
rect 16389 19075 16455 19078
rect 17660 19048 18460 19078
rect 0 18458 800 18488
rect 1485 18458 1551 18461
rect 0 18456 1551 18458
rect 0 18400 1490 18456
rect 1546 18400 1551 18456
rect 0 18398 1551 18400
rect 0 18368 800 18398
rect 1485 18395 1551 18398
rect 6341 17984 6661 17985
rect 6341 17920 6349 17984
rect 6413 17920 6429 17984
rect 6493 17920 6509 17984
rect 6573 17920 6589 17984
rect 6653 17920 6661 17984
rect 6341 17919 6661 17920
rect 11738 17984 12058 17985
rect 11738 17920 11746 17984
rect 11810 17920 11826 17984
rect 11890 17920 11906 17984
rect 11970 17920 11986 17984
rect 12050 17920 12058 17984
rect 11738 17919 12058 17920
rect 3642 17440 3962 17441
rect 3642 17376 3650 17440
rect 3714 17376 3730 17440
rect 3794 17376 3810 17440
rect 3874 17376 3890 17440
rect 3954 17376 3962 17440
rect 3642 17375 3962 17376
rect 9040 17440 9360 17441
rect 9040 17376 9048 17440
rect 9112 17376 9128 17440
rect 9192 17376 9208 17440
rect 9272 17376 9288 17440
rect 9352 17376 9360 17440
rect 9040 17375 9360 17376
rect 14437 17440 14757 17441
rect 14437 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14605 17440
rect 14669 17376 14685 17440
rect 14749 17376 14757 17440
rect 14437 17375 14757 17376
rect 15745 17098 15811 17101
rect 17660 17098 18460 17128
rect 15745 17096 18460 17098
rect 15745 17040 15750 17096
rect 15806 17040 18460 17096
rect 15745 17038 18460 17040
rect 15745 17035 15811 17038
rect 17660 17008 18460 17038
rect 6341 16896 6661 16897
rect 6341 16832 6349 16896
rect 6413 16832 6429 16896
rect 6493 16832 6509 16896
rect 6573 16832 6589 16896
rect 6653 16832 6661 16896
rect 6341 16831 6661 16832
rect 11738 16896 12058 16897
rect 11738 16832 11746 16896
rect 11810 16832 11826 16896
rect 11890 16832 11906 16896
rect 11970 16832 11986 16896
rect 12050 16832 12058 16896
rect 11738 16831 12058 16832
rect 0 16418 800 16448
rect 3141 16418 3207 16421
rect 0 16416 3207 16418
rect 0 16360 3146 16416
rect 3202 16360 3207 16416
rect 0 16358 3207 16360
rect 0 16328 800 16358
rect 3141 16355 3207 16358
rect 3642 16352 3962 16353
rect 3642 16288 3650 16352
rect 3714 16288 3730 16352
rect 3794 16288 3810 16352
rect 3874 16288 3890 16352
rect 3954 16288 3962 16352
rect 3642 16287 3962 16288
rect 9040 16352 9360 16353
rect 9040 16288 9048 16352
rect 9112 16288 9128 16352
rect 9192 16288 9208 16352
rect 9272 16288 9288 16352
rect 9352 16288 9360 16352
rect 9040 16287 9360 16288
rect 14437 16352 14757 16353
rect 14437 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14605 16352
rect 14669 16288 14685 16352
rect 14749 16288 14757 16352
rect 14437 16287 14757 16288
rect 6341 15808 6661 15809
rect 6341 15744 6349 15808
rect 6413 15744 6429 15808
rect 6493 15744 6509 15808
rect 6573 15744 6589 15808
rect 6653 15744 6661 15808
rect 6341 15743 6661 15744
rect 11738 15808 12058 15809
rect 11738 15744 11746 15808
rect 11810 15744 11826 15808
rect 11890 15744 11906 15808
rect 11970 15744 11986 15808
rect 12050 15744 12058 15808
rect 11738 15743 12058 15744
rect 5993 15602 6059 15605
rect 7281 15602 7347 15605
rect 5993 15600 7347 15602
rect 5993 15544 5998 15600
rect 6054 15544 7286 15600
rect 7342 15544 7347 15600
rect 5993 15542 7347 15544
rect 5993 15539 6059 15542
rect 7281 15539 7347 15542
rect 3642 15264 3962 15265
rect 3642 15200 3650 15264
rect 3714 15200 3730 15264
rect 3794 15200 3810 15264
rect 3874 15200 3890 15264
rect 3954 15200 3962 15264
rect 3642 15199 3962 15200
rect 9040 15264 9360 15265
rect 9040 15200 9048 15264
rect 9112 15200 9128 15264
rect 9192 15200 9208 15264
rect 9272 15200 9288 15264
rect 9352 15200 9360 15264
rect 9040 15199 9360 15200
rect 14437 15264 14757 15265
rect 14437 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14605 15264
rect 14669 15200 14685 15264
rect 14749 15200 14757 15264
rect 14437 15199 14757 15200
rect 17033 15058 17099 15061
rect 17660 15058 18460 15088
rect 17033 15056 18460 15058
rect 17033 15000 17038 15056
rect 17094 15000 18460 15056
rect 17033 14998 18460 15000
rect 17033 14995 17099 14998
rect 17660 14968 18460 14998
rect 6341 14720 6661 14721
rect 6341 14656 6349 14720
rect 6413 14656 6429 14720
rect 6493 14656 6509 14720
rect 6573 14656 6589 14720
rect 6653 14656 6661 14720
rect 6341 14655 6661 14656
rect 11738 14720 12058 14721
rect 11738 14656 11746 14720
rect 11810 14656 11826 14720
rect 11890 14656 11906 14720
rect 11970 14656 11986 14720
rect 12050 14656 12058 14720
rect 11738 14655 12058 14656
rect 0 14378 800 14408
rect 3417 14378 3483 14381
rect 0 14376 3483 14378
rect 0 14320 3422 14376
rect 3478 14320 3483 14376
rect 0 14318 3483 14320
rect 0 14288 800 14318
rect 3417 14315 3483 14318
rect 3642 14176 3962 14177
rect 3642 14112 3650 14176
rect 3714 14112 3730 14176
rect 3794 14112 3810 14176
rect 3874 14112 3890 14176
rect 3954 14112 3962 14176
rect 3642 14111 3962 14112
rect 9040 14176 9360 14177
rect 9040 14112 9048 14176
rect 9112 14112 9128 14176
rect 9192 14112 9208 14176
rect 9272 14112 9288 14176
rect 9352 14112 9360 14176
rect 9040 14111 9360 14112
rect 14437 14176 14757 14177
rect 14437 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14605 14176
rect 14669 14112 14685 14176
rect 14749 14112 14757 14176
rect 14437 14111 14757 14112
rect 4337 13970 4403 13973
rect 5165 13970 5231 13973
rect 4337 13968 5231 13970
rect 4337 13912 4342 13968
rect 4398 13912 5170 13968
rect 5226 13912 5231 13968
rect 4337 13910 5231 13912
rect 4337 13907 4403 13910
rect 5165 13907 5231 13910
rect 3601 13834 3667 13837
rect 4889 13834 4955 13837
rect 5993 13834 6059 13837
rect 3601 13832 6059 13834
rect 3601 13776 3606 13832
rect 3662 13776 4894 13832
rect 4950 13776 5998 13832
rect 6054 13776 6059 13832
rect 3601 13774 6059 13776
rect 3601 13771 3667 13774
rect 4889 13771 4955 13774
rect 5993 13771 6059 13774
rect 6341 13632 6661 13633
rect 6341 13568 6349 13632
rect 6413 13568 6429 13632
rect 6493 13568 6509 13632
rect 6573 13568 6589 13632
rect 6653 13568 6661 13632
rect 6341 13567 6661 13568
rect 11738 13632 12058 13633
rect 11738 13568 11746 13632
rect 11810 13568 11826 13632
rect 11890 13568 11906 13632
rect 11970 13568 11986 13632
rect 12050 13568 12058 13632
rect 11738 13567 12058 13568
rect 3642 13088 3962 13089
rect 3642 13024 3650 13088
rect 3714 13024 3730 13088
rect 3794 13024 3810 13088
rect 3874 13024 3890 13088
rect 3954 13024 3962 13088
rect 3642 13023 3962 13024
rect 9040 13088 9360 13089
rect 9040 13024 9048 13088
rect 9112 13024 9128 13088
rect 9192 13024 9208 13088
rect 9272 13024 9288 13088
rect 9352 13024 9360 13088
rect 9040 13023 9360 13024
rect 14437 13088 14757 13089
rect 14437 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14605 13088
rect 14669 13024 14685 13088
rect 14749 13024 14757 13088
rect 14437 13023 14757 13024
rect 16573 13018 16639 13021
rect 17660 13018 18460 13048
rect 16573 13016 18460 13018
rect 16573 12960 16578 13016
rect 16634 12960 18460 13016
rect 16573 12958 18460 12960
rect 16573 12955 16639 12958
rect 17660 12928 18460 12958
rect 6341 12544 6661 12545
rect 6341 12480 6349 12544
rect 6413 12480 6429 12544
rect 6493 12480 6509 12544
rect 6573 12480 6589 12544
rect 6653 12480 6661 12544
rect 6341 12479 6661 12480
rect 11738 12544 12058 12545
rect 11738 12480 11746 12544
rect 11810 12480 11826 12544
rect 11890 12480 11906 12544
rect 11970 12480 11986 12544
rect 12050 12480 12058 12544
rect 11738 12479 12058 12480
rect 0 12338 800 12368
rect 2865 12338 2931 12341
rect 0 12336 2931 12338
rect 0 12280 2870 12336
rect 2926 12280 2931 12336
rect 0 12278 2931 12280
rect 0 12248 800 12278
rect 2865 12275 2931 12278
rect 3141 12338 3207 12341
rect 5809 12338 5875 12341
rect 6545 12338 6611 12341
rect 3141 12336 6611 12338
rect 3141 12280 3146 12336
rect 3202 12280 5814 12336
rect 5870 12280 6550 12336
rect 6606 12280 6611 12336
rect 3141 12278 6611 12280
rect 3141 12275 3207 12278
rect 5809 12275 5875 12278
rect 6545 12275 6611 12278
rect 6545 12202 6611 12205
rect 7005 12202 7071 12205
rect 6545 12200 7071 12202
rect 6545 12144 6550 12200
rect 6606 12144 7010 12200
rect 7066 12144 7071 12200
rect 6545 12142 7071 12144
rect 6545 12139 6611 12142
rect 7005 12139 7071 12142
rect 3642 12000 3962 12001
rect 3642 11936 3650 12000
rect 3714 11936 3730 12000
rect 3794 11936 3810 12000
rect 3874 11936 3890 12000
rect 3954 11936 3962 12000
rect 3642 11935 3962 11936
rect 9040 12000 9360 12001
rect 9040 11936 9048 12000
rect 9112 11936 9128 12000
rect 9192 11936 9208 12000
rect 9272 11936 9288 12000
rect 9352 11936 9360 12000
rect 9040 11935 9360 11936
rect 14437 12000 14757 12001
rect 14437 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14605 12000
rect 14669 11936 14685 12000
rect 14749 11936 14757 12000
rect 14437 11935 14757 11936
rect 5809 11930 5875 11933
rect 7005 11930 7071 11933
rect 5809 11928 7071 11930
rect 5809 11872 5814 11928
rect 5870 11872 7010 11928
rect 7066 11872 7071 11928
rect 5809 11870 7071 11872
rect 5809 11867 5875 11870
rect 7005 11867 7071 11870
rect 4889 11794 4955 11797
rect 6729 11794 6795 11797
rect 4889 11792 6795 11794
rect 4889 11736 4894 11792
rect 4950 11736 6734 11792
rect 6790 11736 6795 11792
rect 4889 11734 6795 11736
rect 4889 11731 4955 11734
rect 6729 11731 6795 11734
rect 6341 11456 6661 11457
rect 6341 11392 6349 11456
rect 6413 11392 6429 11456
rect 6493 11392 6509 11456
rect 6573 11392 6589 11456
rect 6653 11392 6661 11456
rect 6341 11391 6661 11392
rect 11738 11456 12058 11457
rect 11738 11392 11746 11456
rect 11810 11392 11826 11456
rect 11890 11392 11906 11456
rect 11970 11392 11986 11456
rect 12050 11392 12058 11456
rect 11738 11391 12058 11392
rect 14917 10978 14983 10981
rect 17660 10978 18460 11008
rect 14917 10976 18460 10978
rect 14917 10920 14922 10976
rect 14978 10920 18460 10976
rect 14917 10918 18460 10920
rect 14917 10915 14983 10918
rect 3642 10912 3962 10913
rect 3642 10848 3650 10912
rect 3714 10848 3730 10912
rect 3794 10848 3810 10912
rect 3874 10848 3890 10912
rect 3954 10848 3962 10912
rect 3642 10847 3962 10848
rect 9040 10912 9360 10913
rect 9040 10848 9048 10912
rect 9112 10848 9128 10912
rect 9192 10848 9208 10912
rect 9272 10848 9288 10912
rect 9352 10848 9360 10912
rect 9040 10847 9360 10848
rect 14437 10912 14757 10913
rect 14437 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14605 10912
rect 14669 10848 14685 10912
rect 14749 10848 14757 10912
rect 17660 10888 18460 10918
rect 14437 10847 14757 10848
rect 2221 10706 2287 10709
rect 8661 10706 8727 10709
rect 2221 10704 8727 10706
rect 2221 10648 2226 10704
rect 2282 10648 8666 10704
rect 8722 10648 8727 10704
rect 2221 10646 8727 10648
rect 2221 10643 2287 10646
rect 8661 10643 8727 10646
rect 6341 10368 6661 10369
rect 0 10298 800 10328
rect 6341 10304 6349 10368
rect 6413 10304 6429 10368
rect 6493 10304 6509 10368
rect 6573 10304 6589 10368
rect 6653 10304 6661 10368
rect 6341 10303 6661 10304
rect 11738 10368 12058 10369
rect 11738 10304 11746 10368
rect 11810 10304 11826 10368
rect 11890 10304 11906 10368
rect 11970 10304 11986 10368
rect 12050 10304 12058 10368
rect 11738 10303 12058 10304
rect 1485 10298 1551 10301
rect 0 10296 1551 10298
rect 0 10240 1490 10296
rect 1546 10240 1551 10296
rect 0 10238 1551 10240
rect 0 10208 800 10238
rect 1485 10235 1551 10238
rect 3642 9824 3962 9825
rect 3642 9760 3650 9824
rect 3714 9760 3730 9824
rect 3794 9760 3810 9824
rect 3874 9760 3890 9824
rect 3954 9760 3962 9824
rect 3642 9759 3962 9760
rect 9040 9824 9360 9825
rect 9040 9760 9048 9824
rect 9112 9760 9128 9824
rect 9192 9760 9208 9824
rect 9272 9760 9288 9824
rect 9352 9760 9360 9824
rect 9040 9759 9360 9760
rect 14437 9824 14757 9825
rect 14437 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14605 9824
rect 14669 9760 14685 9824
rect 14749 9760 14757 9824
rect 14437 9759 14757 9760
rect 7925 9482 7991 9485
rect 10869 9482 10935 9485
rect 7925 9480 10935 9482
rect 7925 9424 7930 9480
rect 7986 9424 10874 9480
rect 10930 9424 10935 9480
rect 7925 9422 10935 9424
rect 7925 9419 7991 9422
rect 10869 9419 10935 9422
rect 7005 9346 7071 9349
rect 9029 9346 9095 9349
rect 7005 9344 9095 9346
rect 7005 9288 7010 9344
rect 7066 9288 9034 9344
rect 9090 9288 9095 9344
rect 7005 9286 9095 9288
rect 7005 9283 7071 9286
rect 9029 9283 9095 9286
rect 6341 9280 6661 9281
rect 6341 9216 6349 9280
rect 6413 9216 6429 9280
rect 6493 9216 6509 9280
rect 6573 9216 6589 9280
rect 6653 9216 6661 9280
rect 6341 9215 6661 9216
rect 11738 9280 12058 9281
rect 11738 9216 11746 9280
rect 11810 9216 11826 9280
rect 11890 9216 11906 9280
rect 11970 9216 11986 9280
rect 12050 9216 12058 9280
rect 11738 9215 12058 9216
rect 3141 8938 3207 8941
rect 8477 8938 8543 8941
rect 3141 8936 8543 8938
rect 3141 8880 3146 8936
rect 3202 8880 8482 8936
rect 8538 8880 8543 8936
rect 3141 8878 8543 8880
rect 3141 8875 3207 8878
rect 8477 8875 8543 8878
rect 14825 8938 14891 8941
rect 17660 8938 18460 8968
rect 14825 8936 18460 8938
rect 14825 8880 14830 8936
rect 14886 8880 18460 8936
rect 14825 8878 18460 8880
rect 14825 8875 14891 8878
rect 17660 8848 18460 8878
rect 3642 8736 3962 8737
rect 3642 8672 3650 8736
rect 3714 8672 3730 8736
rect 3794 8672 3810 8736
rect 3874 8672 3890 8736
rect 3954 8672 3962 8736
rect 3642 8671 3962 8672
rect 9040 8736 9360 8737
rect 9040 8672 9048 8736
rect 9112 8672 9128 8736
rect 9192 8672 9208 8736
rect 9272 8672 9288 8736
rect 9352 8672 9360 8736
rect 9040 8671 9360 8672
rect 14437 8736 14757 8737
rect 14437 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14605 8736
rect 14669 8672 14685 8736
rect 14749 8672 14757 8736
rect 14437 8671 14757 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 6341 8192 6661 8193
rect 6341 8128 6349 8192
rect 6413 8128 6429 8192
rect 6493 8128 6509 8192
rect 6573 8128 6589 8192
rect 6653 8128 6661 8192
rect 6341 8127 6661 8128
rect 11738 8192 12058 8193
rect 11738 8128 11746 8192
rect 11810 8128 11826 8192
rect 11890 8128 11906 8192
rect 11970 8128 11986 8192
rect 12050 8128 12058 8192
rect 11738 8127 12058 8128
rect 3642 7648 3962 7649
rect 3642 7584 3650 7648
rect 3714 7584 3730 7648
rect 3794 7584 3810 7648
rect 3874 7584 3890 7648
rect 3954 7584 3962 7648
rect 3642 7583 3962 7584
rect 9040 7648 9360 7649
rect 9040 7584 9048 7648
rect 9112 7584 9128 7648
rect 9192 7584 9208 7648
rect 9272 7584 9288 7648
rect 9352 7584 9360 7648
rect 9040 7583 9360 7584
rect 14437 7648 14757 7649
rect 14437 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14605 7648
rect 14669 7584 14685 7648
rect 14749 7584 14757 7648
rect 14437 7583 14757 7584
rect 6341 7104 6661 7105
rect 6341 7040 6349 7104
rect 6413 7040 6429 7104
rect 6493 7040 6509 7104
rect 6573 7040 6589 7104
rect 6653 7040 6661 7104
rect 6341 7039 6661 7040
rect 11738 7104 12058 7105
rect 11738 7040 11746 7104
rect 11810 7040 11826 7104
rect 11890 7040 11906 7104
rect 11970 7040 11986 7104
rect 12050 7040 12058 7104
rect 11738 7039 12058 7040
rect 14365 6898 14431 6901
rect 17660 6898 18460 6928
rect 14365 6896 18460 6898
rect 14365 6840 14370 6896
rect 14426 6840 18460 6896
rect 14365 6838 18460 6840
rect 14365 6835 14431 6838
rect 17660 6808 18460 6838
rect 3642 6560 3962 6561
rect 3642 6496 3650 6560
rect 3714 6496 3730 6560
rect 3794 6496 3810 6560
rect 3874 6496 3890 6560
rect 3954 6496 3962 6560
rect 3642 6495 3962 6496
rect 9040 6560 9360 6561
rect 9040 6496 9048 6560
rect 9112 6496 9128 6560
rect 9192 6496 9208 6560
rect 9272 6496 9288 6560
rect 9352 6496 9360 6560
rect 9040 6495 9360 6496
rect 14437 6560 14757 6561
rect 14437 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14605 6560
rect 14669 6496 14685 6560
rect 14749 6496 14757 6560
rect 14437 6495 14757 6496
rect 0 6218 800 6248
rect 3049 6218 3115 6221
rect 0 6216 3115 6218
rect 0 6160 3054 6216
rect 3110 6160 3115 6216
rect 0 6158 3115 6160
rect 0 6128 800 6158
rect 3049 6155 3115 6158
rect 6341 6016 6661 6017
rect 6341 5952 6349 6016
rect 6413 5952 6429 6016
rect 6493 5952 6509 6016
rect 6573 5952 6589 6016
rect 6653 5952 6661 6016
rect 6341 5951 6661 5952
rect 11738 6016 12058 6017
rect 11738 5952 11746 6016
rect 11810 5952 11826 6016
rect 11890 5952 11906 6016
rect 11970 5952 11986 6016
rect 12050 5952 12058 6016
rect 11738 5951 12058 5952
rect 4613 5810 4679 5813
rect 7649 5810 7715 5813
rect 4613 5808 7715 5810
rect 4613 5752 4618 5808
rect 4674 5752 7654 5808
rect 7710 5752 7715 5808
rect 4613 5750 7715 5752
rect 4613 5747 4679 5750
rect 7649 5747 7715 5750
rect 3642 5472 3962 5473
rect 3642 5408 3650 5472
rect 3714 5408 3730 5472
rect 3794 5408 3810 5472
rect 3874 5408 3890 5472
rect 3954 5408 3962 5472
rect 3642 5407 3962 5408
rect 9040 5472 9360 5473
rect 9040 5408 9048 5472
rect 9112 5408 9128 5472
rect 9192 5408 9208 5472
rect 9272 5408 9288 5472
rect 9352 5408 9360 5472
rect 9040 5407 9360 5408
rect 14437 5472 14757 5473
rect 14437 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14605 5472
rect 14669 5408 14685 5472
rect 14749 5408 14757 5472
rect 14437 5407 14757 5408
rect 6341 4928 6661 4929
rect 6341 4864 6349 4928
rect 6413 4864 6429 4928
rect 6493 4864 6509 4928
rect 6573 4864 6589 4928
rect 6653 4864 6661 4928
rect 6341 4863 6661 4864
rect 11738 4928 12058 4929
rect 11738 4864 11746 4928
rect 11810 4864 11826 4928
rect 11890 4864 11906 4928
rect 11970 4864 11986 4928
rect 12050 4864 12058 4928
rect 11738 4863 12058 4864
rect 15101 4858 15167 4861
rect 17660 4858 18460 4888
rect 15101 4856 18460 4858
rect 15101 4800 15106 4856
rect 15162 4800 18460 4856
rect 15101 4798 18460 4800
rect 15101 4795 15167 4798
rect 17660 4768 18460 4798
rect 3642 4384 3962 4385
rect 3642 4320 3650 4384
rect 3714 4320 3730 4384
rect 3794 4320 3810 4384
rect 3874 4320 3890 4384
rect 3954 4320 3962 4384
rect 3642 4319 3962 4320
rect 9040 4384 9360 4385
rect 9040 4320 9048 4384
rect 9112 4320 9128 4384
rect 9192 4320 9208 4384
rect 9272 4320 9288 4384
rect 9352 4320 9360 4384
rect 9040 4319 9360 4320
rect 14437 4384 14757 4385
rect 14437 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14605 4384
rect 14669 4320 14685 4384
rect 14749 4320 14757 4384
rect 14437 4319 14757 4320
rect 0 4178 800 4208
rect 1393 4178 1459 4181
rect 0 4176 1459 4178
rect 0 4120 1398 4176
rect 1454 4120 1459 4176
rect 0 4118 1459 4120
rect 0 4088 800 4118
rect 1393 4115 1459 4118
rect 6341 3840 6661 3841
rect 6341 3776 6349 3840
rect 6413 3776 6429 3840
rect 6493 3776 6509 3840
rect 6573 3776 6589 3840
rect 6653 3776 6661 3840
rect 6341 3775 6661 3776
rect 11738 3840 12058 3841
rect 11738 3776 11746 3840
rect 11810 3776 11826 3840
rect 11890 3776 11906 3840
rect 11970 3776 11986 3840
rect 12050 3776 12058 3840
rect 11738 3775 12058 3776
rect 6913 3770 6979 3773
rect 8753 3770 8819 3773
rect 6913 3768 8819 3770
rect 6913 3712 6918 3768
rect 6974 3712 8758 3768
rect 8814 3712 8819 3768
rect 6913 3710 8819 3712
rect 6913 3707 6979 3710
rect 8753 3707 8819 3710
rect 3325 3634 3391 3637
rect 8385 3634 8451 3637
rect 3325 3632 8451 3634
rect 3325 3576 3330 3632
rect 3386 3576 8390 3632
rect 8446 3576 8451 3632
rect 3325 3574 8451 3576
rect 3325 3571 3391 3574
rect 8385 3571 8451 3574
rect 5809 3498 5875 3501
rect 6361 3498 6427 3501
rect 5809 3496 6427 3498
rect 5809 3440 5814 3496
rect 5870 3440 6366 3496
rect 6422 3440 6427 3496
rect 5809 3438 6427 3440
rect 5809 3435 5875 3438
rect 6361 3435 6427 3438
rect 3642 3296 3962 3297
rect 3642 3232 3650 3296
rect 3714 3232 3730 3296
rect 3794 3232 3810 3296
rect 3874 3232 3890 3296
rect 3954 3232 3962 3296
rect 3642 3231 3962 3232
rect 9040 3296 9360 3297
rect 9040 3232 9048 3296
rect 9112 3232 9128 3296
rect 9192 3232 9208 3296
rect 9272 3232 9288 3296
rect 9352 3232 9360 3296
rect 9040 3231 9360 3232
rect 14437 3296 14757 3297
rect 14437 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14605 3296
rect 14669 3232 14685 3296
rect 14749 3232 14757 3296
rect 14437 3231 14757 3232
rect 14365 2818 14431 2821
rect 17660 2818 18460 2848
rect 14365 2816 18460 2818
rect 14365 2760 14370 2816
rect 14426 2760 18460 2816
rect 14365 2758 18460 2760
rect 14365 2755 14431 2758
rect 6341 2752 6661 2753
rect 6341 2688 6349 2752
rect 6413 2688 6429 2752
rect 6493 2688 6509 2752
rect 6573 2688 6589 2752
rect 6653 2688 6661 2752
rect 6341 2687 6661 2688
rect 11738 2752 12058 2753
rect 11738 2688 11746 2752
rect 11810 2688 11826 2752
rect 11890 2688 11906 2752
rect 11970 2688 11986 2752
rect 12050 2688 12058 2752
rect 17660 2728 18460 2758
rect 11738 2687 12058 2688
rect 3642 2208 3962 2209
rect 0 2138 800 2168
rect 3642 2144 3650 2208
rect 3714 2144 3730 2208
rect 3794 2144 3810 2208
rect 3874 2144 3890 2208
rect 3954 2144 3962 2208
rect 3642 2143 3962 2144
rect 9040 2208 9360 2209
rect 9040 2144 9048 2208
rect 9112 2144 9128 2208
rect 9192 2144 9208 2208
rect 9272 2144 9288 2208
rect 9352 2144 9360 2208
rect 9040 2143 9360 2144
rect 14437 2208 14757 2209
rect 14437 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14605 2208
rect 14669 2144 14685 2208
rect 14749 2144 14757 2208
rect 14437 2143 14757 2144
rect 2865 2138 2931 2141
rect 0 2136 2931 2138
rect 0 2080 2870 2136
rect 2926 2080 2931 2136
rect 0 2078 2931 2080
rect 0 2048 800 2078
rect 2865 2075 2931 2078
rect 15745 778 15811 781
rect 17660 778 18460 808
rect 15745 776 18460 778
rect 15745 720 15750 776
rect 15806 720 18460 776
rect 15745 718 18460 720
rect 15745 715 15811 718
rect 17660 688 18460 718
<< via3 >>
rect 6349 17980 6413 17984
rect 6349 17924 6353 17980
rect 6353 17924 6409 17980
rect 6409 17924 6413 17980
rect 6349 17920 6413 17924
rect 6429 17980 6493 17984
rect 6429 17924 6433 17980
rect 6433 17924 6489 17980
rect 6489 17924 6493 17980
rect 6429 17920 6493 17924
rect 6509 17980 6573 17984
rect 6509 17924 6513 17980
rect 6513 17924 6569 17980
rect 6569 17924 6573 17980
rect 6509 17920 6573 17924
rect 6589 17980 6653 17984
rect 6589 17924 6593 17980
rect 6593 17924 6649 17980
rect 6649 17924 6653 17980
rect 6589 17920 6653 17924
rect 11746 17980 11810 17984
rect 11746 17924 11750 17980
rect 11750 17924 11806 17980
rect 11806 17924 11810 17980
rect 11746 17920 11810 17924
rect 11826 17980 11890 17984
rect 11826 17924 11830 17980
rect 11830 17924 11886 17980
rect 11886 17924 11890 17980
rect 11826 17920 11890 17924
rect 11906 17980 11970 17984
rect 11906 17924 11910 17980
rect 11910 17924 11966 17980
rect 11966 17924 11970 17980
rect 11906 17920 11970 17924
rect 11986 17980 12050 17984
rect 11986 17924 11990 17980
rect 11990 17924 12046 17980
rect 12046 17924 12050 17980
rect 11986 17920 12050 17924
rect 3650 17436 3714 17440
rect 3650 17380 3654 17436
rect 3654 17380 3710 17436
rect 3710 17380 3714 17436
rect 3650 17376 3714 17380
rect 3730 17436 3794 17440
rect 3730 17380 3734 17436
rect 3734 17380 3790 17436
rect 3790 17380 3794 17436
rect 3730 17376 3794 17380
rect 3810 17436 3874 17440
rect 3810 17380 3814 17436
rect 3814 17380 3870 17436
rect 3870 17380 3874 17436
rect 3810 17376 3874 17380
rect 3890 17436 3954 17440
rect 3890 17380 3894 17436
rect 3894 17380 3950 17436
rect 3950 17380 3954 17436
rect 3890 17376 3954 17380
rect 9048 17436 9112 17440
rect 9048 17380 9052 17436
rect 9052 17380 9108 17436
rect 9108 17380 9112 17436
rect 9048 17376 9112 17380
rect 9128 17436 9192 17440
rect 9128 17380 9132 17436
rect 9132 17380 9188 17436
rect 9188 17380 9192 17436
rect 9128 17376 9192 17380
rect 9208 17436 9272 17440
rect 9208 17380 9212 17436
rect 9212 17380 9268 17436
rect 9268 17380 9272 17436
rect 9208 17376 9272 17380
rect 9288 17436 9352 17440
rect 9288 17380 9292 17436
rect 9292 17380 9348 17436
rect 9348 17380 9352 17436
rect 9288 17376 9352 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 14605 17436 14669 17440
rect 14605 17380 14609 17436
rect 14609 17380 14665 17436
rect 14665 17380 14669 17436
rect 14605 17376 14669 17380
rect 14685 17436 14749 17440
rect 14685 17380 14689 17436
rect 14689 17380 14745 17436
rect 14745 17380 14749 17436
rect 14685 17376 14749 17380
rect 6349 16892 6413 16896
rect 6349 16836 6353 16892
rect 6353 16836 6409 16892
rect 6409 16836 6413 16892
rect 6349 16832 6413 16836
rect 6429 16892 6493 16896
rect 6429 16836 6433 16892
rect 6433 16836 6489 16892
rect 6489 16836 6493 16892
rect 6429 16832 6493 16836
rect 6509 16892 6573 16896
rect 6509 16836 6513 16892
rect 6513 16836 6569 16892
rect 6569 16836 6573 16892
rect 6509 16832 6573 16836
rect 6589 16892 6653 16896
rect 6589 16836 6593 16892
rect 6593 16836 6649 16892
rect 6649 16836 6653 16892
rect 6589 16832 6653 16836
rect 11746 16892 11810 16896
rect 11746 16836 11750 16892
rect 11750 16836 11806 16892
rect 11806 16836 11810 16892
rect 11746 16832 11810 16836
rect 11826 16892 11890 16896
rect 11826 16836 11830 16892
rect 11830 16836 11886 16892
rect 11886 16836 11890 16892
rect 11826 16832 11890 16836
rect 11906 16892 11970 16896
rect 11906 16836 11910 16892
rect 11910 16836 11966 16892
rect 11966 16836 11970 16892
rect 11906 16832 11970 16836
rect 11986 16892 12050 16896
rect 11986 16836 11990 16892
rect 11990 16836 12046 16892
rect 12046 16836 12050 16892
rect 11986 16832 12050 16836
rect 3650 16348 3714 16352
rect 3650 16292 3654 16348
rect 3654 16292 3710 16348
rect 3710 16292 3714 16348
rect 3650 16288 3714 16292
rect 3730 16348 3794 16352
rect 3730 16292 3734 16348
rect 3734 16292 3790 16348
rect 3790 16292 3794 16348
rect 3730 16288 3794 16292
rect 3810 16348 3874 16352
rect 3810 16292 3814 16348
rect 3814 16292 3870 16348
rect 3870 16292 3874 16348
rect 3810 16288 3874 16292
rect 3890 16348 3954 16352
rect 3890 16292 3894 16348
rect 3894 16292 3950 16348
rect 3950 16292 3954 16348
rect 3890 16288 3954 16292
rect 9048 16348 9112 16352
rect 9048 16292 9052 16348
rect 9052 16292 9108 16348
rect 9108 16292 9112 16348
rect 9048 16288 9112 16292
rect 9128 16348 9192 16352
rect 9128 16292 9132 16348
rect 9132 16292 9188 16348
rect 9188 16292 9192 16348
rect 9128 16288 9192 16292
rect 9208 16348 9272 16352
rect 9208 16292 9212 16348
rect 9212 16292 9268 16348
rect 9268 16292 9272 16348
rect 9208 16288 9272 16292
rect 9288 16348 9352 16352
rect 9288 16292 9292 16348
rect 9292 16292 9348 16348
rect 9348 16292 9352 16348
rect 9288 16288 9352 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 14605 16348 14669 16352
rect 14605 16292 14609 16348
rect 14609 16292 14665 16348
rect 14665 16292 14669 16348
rect 14605 16288 14669 16292
rect 14685 16348 14749 16352
rect 14685 16292 14689 16348
rect 14689 16292 14745 16348
rect 14745 16292 14749 16348
rect 14685 16288 14749 16292
rect 6349 15804 6413 15808
rect 6349 15748 6353 15804
rect 6353 15748 6409 15804
rect 6409 15748 6413 15804
rect 6349 15744 6413 15748
rect 6429 15804 6493 15808
rect 6429 15748 6433 15804
rect 6433 15748 6489 15804
rect 6489 15748 6493 15804
rect 6429 15744 6493 15748
rect 6509 15804 6573 15808
rect 6509 15748 6513 15804
rect 6513 15748 6569 15804
rect 6569 15748 6573 15804
rect 6509 15744 6573 15748
rect 6589 15804 6653 15808
rect 6589 15748 6593 15804
rect 6593 15748 6649 15804
rect 6649 15748 6653 15804
rect 6589 15744 6653 15748
rect 11746 15804 11810 15808
rect 11746 15748 11750 15804
rect 11750 15748 11806 15804
rect 11806 15748 11810 15804
rect 11746 15744 11810 15748
rect 11826 15804 11890 15808
rect 11826 15748 11830 15804
rect 11830 15748 11886 15804
rect 11886 15748 11890 15804
rect 11826 15744 11890 15748
rect 11906 15804 11970 15808
rect 11906 15748 11910 15804
rect 11910 15748 11966 15804
rect 11966 15748 11970 15804
rect 11906 15744 11970 15748
rect 11986 15804 12050 15808
rect 11986 15748 11990 15804
rect 11990 15748 12046 15804
rect 12046 15748 12050 15804
rect 11986 15744 12050 15748
rect 3650 15260 3714 15264
rect 3650 15204 3654 15260
rect 3654 15204 3710 15260
rect 3710 15204 3714 15260
rect 3650 15200 3714 15204
rect 3730 15260 3794 15264
rect 3730 15204 3734 15260
rect 3734 15204 3790 15260
rect 3790 15204 3794 15260
rect 3730 15200 3794 15204
rect 3810 15260 3874 15264
rect 3810 15204 3814 15260
rect 3814 15204 3870 15260
rect 3870 15204 3874 15260
rect 3810 15200 3874 15204
rect 3890 15260 3954 15264
rect 3890 15204 3894 15260
rect 3894 15204 3950 15260
rect 3950 15204 3954 15260
rect 3890 15200 3954 15204
rect 9048 15260 9112 15264
rect 9048 15204 9052 15260
rect 9052 15204 9108 15260
rect 9108 15204 9112 15260
rect 9048 15200 9112 15204
rect 9128 15260 9192 15264
rect 9128 15204 9132 15260
rect 9132 15204 9188 15260
rect 9188 15204 9192 15260
rect 9128 15200 9192 15204
rect 9208 15260 9272 15264
rect 9208 15204 9212 15260
rect 9212 15204 9268 15260
rect 9268 15204 9272 15260
rect 9208 15200 9272 15204
rect 9288 15260 9352 15264
rect 9288 15204 9292 15260
rect 9292 15204 9348 15260
rect 9348 15204 9352 15260
rect 9288 15200 9352 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 14605 15260 14669 15264
rect 14605 15204 14609 15260
rect 14609 15204 14665 15260
rect 14665 15204 14669 15260
rect 14605 15200 14669 15204
rect 14685 15260 14749 15264
rect 14685 15204 14689 15260
rect 14689 15204 14745 15260
rect 14745 15204 14749 15260
rect 14685 15200 14749 15204
rect 6349 14716 6413 14720
rect 6349 14660 6353 14716
rect 6353 14660 6409 14716
rect 6409 14660 6413 14716
rect 6349 14656 6413 14660
rect 6429 14716 6493 14720
rect 6429 14660 6433 14716
rect 6433 14660 6489 14716
rect 6489 14660 6493 14716
rect 6429 14656 6493 14660
rect 6509 14716 6573 14720
rect 6509 14660 6513 14716
rect 6513 14660 6569 14716
rect 6569 14660 6573 14716
rect 6509 14656 6573 14660
rect 6589 14716 6653 14720
rect 6589 14660 6593 14716
rect 6593 14660 6649 14716
rect 6649 14660 6653 14716
rect 6589 14656 6653 14660
rect 11746 14716 11810 14720
rect 11746 14660 11750 14716
rect 11750 14660 11806 14716
rect 11806 14660 11810 14716
rect 11746 14656 11810 14660
rect 11826 14716 11890 14720
rect 11826 14660 11830 14716
rect 11830 14660 11886 14716
rect 11886 14660 11890 14716
rect 11826 14656 11890 14660
rect 11906 14716 11970 14720
rect 11906 14660 11910 14716
rect 11910 14660 11966 14716
rect 11966 14660 11970 14716
rect 11906 14656 11970 14660
rect 11986 14716 12050 14720
rect 11986 14660 11990 14716
rect 11990 14660 12046 14716
rect 12046 14660 12050 14716
rect 11986 14656 12050 14660
rect 3650 14172 3714 14176
rect 3650 14116 3654 14172
rect 3654 14116 3710 14172
rect 3710 14116 3714 14172
rect 3650 14112 3714 14116
rect 3730 14172 3794 14176
rect 3730 14116 3734 14172
rect 3734 14116 3790 14172
rect 3790 14116 3794 14172
rect 3730 14112 3794 14116
rect 3810 14172 3874 14176
rect 3810 14116 3814 14172
rect 3814 14116 3870 14172
rect 3870 14116 3874 14172
rect 3810 14112 3874 14116
rect 3890 14172 3954 14176
rect 3890 14116 3894 14172
rect 3894 14116 3950 14172
rect 3950 14116 3954 14172
rect 3890 14112 3954 14116
rect 9048 14172 9112 14176
rect 9048 14116 9052 14172
rect 9052 14116 9108 14172
rect 9108 14116 9112 14172
rect 9048 14112 9112 14116
rect 9128 14172 9192 14176
rect 9128 14116 9132 14172
rect 9132 14116 9188 14172
rect 9188 14116 9192 14172
rect 9128 14112 9192 14116
rect 9208 14172 9272 14176
rect 9208 14116 9212 14172
rect 9212 14116 9268 14172
rect 9268 14116 9272 14172
rect 9208 14112 9272 14116
rect 9288 14172 9352 14176
rect 9288 14116 9292 14172
rect 9292 14116 9348 14172
rect 9348 14116 9352 14172
rect 9288 14112 9352 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 14605 14172 14669 14176
rect 14605 14116 14609 14172
rect 14609 14116 14665 14172
rect 14665 14116 14669 14172
rect 14605 14112 14669 14116
rect 14685 14172 14749 14176
rect 14685 14116 14689 14172
rect 14689 14116 14745 14172
rect 14745 14116 14749 14172
rect 14685 14112 14749 14116
rect 6349 13628 6413 13632
rect 6349 13572 6353 13628
rect 6353 13572 6409 13628
rect 6409 13572 6413 13628
rect 6349 13568 6413 13572
rect 6429 13628 6493 13632
rect 6429 13572 6433 13628
rect 6433 13572 6489 13628
rect 6489 13572 6493 13628
rect 6429 13568 6493 13572
rect 6509 13628 6573 13632
rect 6509 13572 6513 13628
rect 6513 13572 6569 13628
rect 6569 13572 6573 13628
rect 6509 13568 6573 13572
rect 6589 13628 6653 13632
rect 6589 13572 6593 13628
rect 6593 13572 6649 13628
rect 6649 13572 6653 13628
rect 6589 13568 6653 13572
rect 11746 13628 11810 13632
rect 11746 13572 11750 13628
rect 11750 13572 11806 13628
rect 11806 13572 11810 13628
rect 11746 13568 11810 13572
rect 11826 13628 11890 13632
rect 11826 13572 11830 13628
rect 11830 13572 11886 13628
rect 11886 13572 11890 13628
rect 11826 13568 11890 13572
rect 11906 13628 11970 13632
rect 11906 13572 11910 13628
rect 11910 13572 11966 13628
rect 11966 13572 11970 13628
rect 11906 13568 11970 13572
rect 11986 13628 12050 13632
rect 11986 13572 11990 13628
rect 11990 13572 12046 13628
rect 12046 13572 12050 13628
rect 11986 13568 12050 13572
rect 3650 13084 3714 13088
rect 3650 13028 3654 13084
rect 3654 13028 3710 13084
rect 3710 13028 3714 13084
rect 3650 13024 3714 13028
rect 3730 13084 3794 13088
rect 3730 13028 3734 13084
rect 3734 13028 3790 13084
rect 3790 13028 3794 13084
rect 3730 13024 3794 13028
rect 3810 13084 3874 13088
rect 3810 13028 3814 13084
rect 3814 13028 3870 13084
rect 3870 13028 3874 13084
rect 3810 13024 3874 13028
rect 3890 13084 3954 13088
rect 3890 13028 3894 13084
rect 3894 13028 3950 13084
rect 3950 13028 3954 13084
rect 3890 13024 3954 13028
rect 9048 13084 9112 13088
rect 9048 13028 9052 13084
rect 9052 13028 9108 13084
rect 9108 13028 9112 13084
rect 9048 13024 9112 13028
rect 9128 13084 9192 13088
rect 9128 13028 9132 13084
rect 9132 13028 9188 13084
rect 9188 13028 9192 13084
rect 9128 13024 9192 13028
rect 9208 13084 9272 13088
rect 9208 13028 9212 13084
rect 9212 13028 9268 13084
rect 9268 13028 9272 13084
rect 9208 13024 9272 13028
rect 9288 13084 9352 13088
rect 9288 13028 9292 13084
rect 9292 13028 9348 13084
rect 9348 13028 9352 13084
rect 9288 13024 9352 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 14605 13084 14669 13088
rect 14605 13028 14609 13084
rect 14609 13028 14665 13084
rect 14665 13028 14669 13084
rect 14605 13024 14669 13028
rect 14685 13084 14749 13088
rect 14685 13028 14689 13084
rect 14689 13028 14745 13084
rect 14745 13028 14749 13084
rect 14685 13024 14749 13028
rect 6349 12540 6413 12544
rect 6349 12484 6353 12540
rect 6353 12484 6409 12540
rect 6409 12484 6413 12540
rect 6349 12480 6413 12484
rect 6429 12540 6493 12544
rect 6429 12484 6433 12540
rect 6433 12484 6489 12540
rect 6489 12484 6493 12540
rect 6429 12480 6493 12484
rect 6509 12540 6573 12544
rect 6509 12484 6513 12540
rect 6513 12484 6569 12540
rect 6569 12484 6573 12540
rect 6509 12480 6573 12484
rect 6589 12540 6653 12544
rect 6589 12484 6593 12540
rect 6593 12484 6649 12540
rect 6649 12484 6653 12540
rect 6589 12480 6653 12484
rect 11746 12540 11810 12544
rect 11746 12484 11750 12540
rect 11750 12484 11806 12540
rect 11806 12484 11810 12540
rect 11746 12480 11810 12484
rect 11826 12540 11890 12544
rect 11826 12484 11830 12540
rect 11830 12484 11886 12540
rect 11886 12484 11890 12540
rect 11826 12480 11890 12484
rect 11906 12540 11970 12544
rect 11906 12484 11910 12540
rect 11910 12484 11966 12540
rect 11966 12484 11970 12540
rect 11906 12480 11970 12484
rect 11986 12540 12050 12544
rect 11986 12484 11990 12540
rect 11990 12484 12046 12540
rect 12046 12484 12050 12540
rect 11986 12480 12050 12484
rect 3650 11996 3714 12000
rect 3650 11940 3654 11996
rect 3654 11940 3710 11996
rect 3710 11940 3714 11996
rect 3650 11936 3714 11940
rect 3730 11996 3794 12000
rect 3730 11940 3734 11996
rect 3734 11940 3790 11996
rect 3790 11940 3794 11996
rect 3730 11936 3794 11940
rect 3810 11996 3874 12000
rect 3810 11940 3814 11996
rect 3814 11940 3870 11996
rect 3870 11940 3874 11996
rect 3810 11936 3874 11940
rect 3890 11996 3954 12000
rect 3890 11940 3894 11996
rect 3894 11940 3950 11996
rect 3950 11940 3954 11996
rect 3890 11936 3954 11940
rect 9048 11996 9112 12000
rect 9048 11940 9052 11996
rect 9052 11940 9108 11996
rect 9108 11940 9112 11996
rect 9048 11936 9112 11940
rect 9128 11996 9192 12000
rect 9128 11940 9132 11996
rect 9132 11940 9188 11996
rect 9188 11940 9192 11996
rect 9128 11936 9192 11940
rect 9208 11996 9272 12000
rect 9208 11940 9212 11996
rect 9212 11940 9268 11996
rect 9268 11940 9272 11996
rect 9208 11936 9272 11940
rect 9288 11996 9352 12000
rect 9288 11940 9292 11996
rect 9292 11940 9348 11996
rect 9348 11940 9352 11996
rect 9288 11936 9352 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 14605 11996 14669 12000
rect 14605 11940 14609 11996
rect 14609 11940 14665 11996
rect 14665 11940 14669 11996
rect 14605 11936 14669 11940
rect 14685 11996 14749 12000
rect 14685 11940 14689 11996
rect 14689 11940 14745 11996
rect 14745 11940 14749 11996
rect 14685 11936 14749 11940
rect 6349 11452 6413 11456
rect 6349 11396 6353 11452
rect 6353 11396 6409 11452
rect 6409 11396 6413 11452
rect 6349 11392 6413 11396
rect 6429 11452 6493 11456
rect 6429 11396 6433 11452
rect 6433 11396 6489 11452
rect 6489 11396 6493 11452
rect 6429 11392 6493 11396
rect 6509 11452 6573 11456
rect 6509 11396 6513 11452
rect 6513 11396 6569 11452
rect 6569 11396 6573 11452
rect 6509 11392 6573 11396
rect 6589 11452 6653 11456
rect 6589 11396 6593 11452
rect 6593 11396 6649 11452
rect 6649 11396 6653 11452
rect 6589 11392 6653 11396
rect 11746 11452 11810 11456
rect 11746 11396 11750 11452
rect 11750 11396 11806 11452
rect 11806 11396 11810 11452
rect 11746 11392 11810 11396
rect 11826 11452 11890 11456
rect 11826 11396 11830 11452
rect 11830 11396 11886 11452
rect 11886 11396 11890 11452
rect 11826 11392 11890 11396
rect 11906 11452 11970 11456
rect 11906 11396 11910 11452
rect 11910 11396 11966 11452
rect 11966 11396 11970 11452
rect 11906 11392 11970 11396
rect 11986 11452 12050 11456
rect 11986 11396 11990 11452
rect 11990 11396 12046 11452
rect 12046 11396 12050 11452
rect 11986 11392 12050 11396
rect 3650 10908 3714 10912
rect 3650 10852 3654 10908
rect 3654 10852 3710 10908
rect 3710 10852 3714 10908
rect 3650 10848 3714 10852
rect 3730 10908 3794 10912
rect 3730 10852 3734 10908
rect 3734 10852 3790 10908
rect 3790 10852 3794 10908
rect 3730 10848 3794 10852
rect 3810 10908 3874 10912
rect 3810 10852 3814 10908
rect 3814 10852 3870 10908
rect 3870 10852 3874 10908
rect 3810 10848 3874 10852
rect 3890 10908 3954 10912
rect 3890 10852 3894 10908
rect 3894 10852 3950 10908
rect 3950 10852 3954 10908
rect 3890 10848 3954 10852
rect 9048 10908 9112 10912
rect 9048 10852 9052 10908
rect 9052 10852 9108 10908
rect 9108 10852 9112 10908
rect 9048 10848 9112 10852
rect 9128 10908 9192 10912
rect 9128 10852 9132 10908
rect 9132 10852 9188 10908
rect 9188 10852 9192 10908
rect 9128 10848 9192 10852
rect 9208 10908 9272 10912
rect 9208 10852 9212 10908
rect 9212 10852 9268 10908
rect 9268 10852 9272 10908
rect 9208 10848 9272 10852
rect 9288 10908 9352 10912
rect 9288 10852 9292 10908
rect 9292 10852 9348 10908
rect 9348 10852 9352 10908
rect 9288 10848 9352 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 14605 10908 14669 10912
rect 14605 10852 14609 10908
rect 14609 10852 14665 10908
rect 14665 10852 14669 10908
rect 14605 10848 14669 10852
rect 14685 10908 14749 10912
rect 14685 10852 14689 10908
rect 14689 10852 14745 10908
rect 14745 10852 14749 10908
rect 14685 10848 14749 10852
rect 6349 10364 6413 10368
rect 6349 10308 6353 10364
rect 6353 10308 6409 10364
rect 6409 10308 6413 10364
rect 6349 10304 6413 10308
rect 6429 10364 6493 10368
rect 6429 10308 6433 10364
rect 6433 10308 6489 10364
rect 6489 10308 6493 10364
rect 6429 10304 6493 10308
rect 6509 10364 6573 10368
rect 6509 10308 6513 10364
rect 6513 10308 6569 10364
rect 6569 10308 6573 10364
rect 6509 10304 6573 10308
rect 6589 10364 6653 10368
rect 6589 10308 6593 10364
rect 6593 10308 6649 10364
rect 6649 10308 6653 10364
rect 6589 10304 6653 10308
rect 11746 10364 11810 10368
rect 11746 10308 11750 10364
rect 11750 10308 11806 10364
rect 11806 10308 11810 10364
rect 11746 10304 11810 10308
rect 11826 10364 11890 10368
rect 11826 10308 11830 10364
rect 11830 10308 11886 10364
rect 11886 10308 11890 10364
rect 11826 10304 11890 10308
rect 11906 10364 11970 10368
rect 11906 10308 11910 10364
rect 11910 10308 11966 10364
rect 11966 10308 11970 10364
rect 11906 10304 11970 10308
rect 11986 10364 12050 10368
rect 11986 10308 11990 10364
rect 11990 10308 12046 10364
rect 12046 10308 12050 10364
rect 11986 10304 12050 10308
rect 3650 9820 3714 9824
rect 3650 9764 3654 9820
rect 3654 9764 3710 9820
rect 3710 9764 3714 9820
rect 3650 9760 3714 9764
rect 3730 9820 3794 9824
rect 3730 9764 3734 9820
rect 3734 9764 3790 9820
rect 3790 9764 3794 9820
rect 3730 9760 3794 9764
rect 3810 9820 3874 9824
rect 3810 9764 3814 9820
rect 3814 9764 3870 9820
rect 3870 9764 3874 9820
rect 3810 9760 3874 9764
rect 3890 9820 3954 9824
rect 3890 9764 3894 9820
rect 3894 9764 3950 9820
rect 3950 9764 3954 9820
rect 3890 9760 3954 9764
rect 9048 9820 9112 9824
rect 9048 9764 9052 9820
rect 9052 9764 9108 9820
rect 9108 9764 9112 9820
rect 9048 9760 9112 9764
rect 9128 9820 9192 9824
rect 9128 9764 9132 9820
rect 9132 9764 9188 9820
rect 9188 9764 9192 9820
rect 9128 9760 9192 9764
rect 9208 9820 9272 9824
rect 9208 9764 9212 9820
rect 9212 9764 9268 9820
rect 9268 9764 9272 9820
rect 9208 9760 9272 9764
rect 9288 9820 9352 9824
rect 9288 9764 9292 9820
rect 9292 9764 9348 9820
rect 9348 9764 9352 9820
rect 9288 9760 9352 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 14605 9820 14669 9824
rect 14605 9764 14609 9820
rect 14609 9764 14665 9820
rect 14665 9764 14669 9820
rect 14605 9760 14669 9764
rect 14685 9820 14749 9824
rect 14685 9764 14689 9820
rect 14689 9764 14745 9820
rect 14745 9764 14749 9820
rect 14685 9760 14749 9764
rect 6349 9276 6413 9280
rect 6349 9220 6353 9276
rect 6353 9220 6409 9276
rect 6409 9220 6413 9276
rect 6349 9216 6413 9220
rect 6429 9276 6493 9280
rect 6429 9220 6433 9276
rect 6433 9220 6489 9276
rect 6489 9220 6493 9276
rect 6429 9216 6493 9220
rect 6509 9276 6573 9280
rect 6509 9220 6513 9276
rect 6513 9220 6569 9276
rect 6569 9220 6573 9276
rect 6509 9216 6573 9220
rect 6589 9276 6653 9280
rect 6589 9220 6593 9276
rect 6593 9220 6649 9276
rect 6649 9220 6653 9276
rect 6589 9216 6653 9220
rect 11746 9276 11810 9280
rect 11746 9220 11750 9276
rect 11750 9220 11806 9276
rect 11806 9220 11810 9276
rect 11746 9216 11810 9220
rect 11826 9276 11890 9280
rect 11826 9220 11830 9276
rect 11830 9220 11886 9276
rect 11886 9220 11890 9276
rect 11826 9216 11890 9220
rect 11906 9276 11970 9280
rect 11906 9220 11910 9276
rect 11910 9220 11966 9276
rect 11966 9220 11970 9276
rect 11906 9216 11970 9220
rect 11986 9276 12050 9280
rect 11986 9220 11990 9276
rect 11990 9220 12046 9276
rect 12046 9220 12050 9276
rect 11986 9216 12050 9220
rect 3650 8732 3714 8736
rect 3650 8676 3654 8732
rect 3654 8676 3710 8732
rect 3710 8676 3714 8732
rect 3650 8672 3714 8676
rect 3730 8732 3794 8736
rect 3730 8676 3734 8732
rect 3734 8676 3790 8732
rect 3790 8676 3794 8732
rect 3730 8672 3794 8676
rect 3810 8732 3874 8736
rect 3810 8676 3814 8732
rect 3814 8676 3870 8732
rect 3870 8676 3874 8732
rect 3810 8672 3874 8676
rect 3890 8732 3954 8736
rect 3890 8676 3894 8732
rect 3894 8676 3950 8732
rect 3950 8676 3954 8732
rect 3890 8672 3954 8676
rect 9048 8732 9112 8736
rect 9048 8676 9052 8732
rect 9052 8676 9108 8732
rect 9108 8676 9112 8732
rect 9048 8672 9112 8676
rect 9128 8732 9192 8736
rect 9128 8676 9132 8732
rect 9132 8676 9188 8732
rect 9188 8676 9192 8732
rect 9128 8672 9192 8676
rect 9208 8732 9272 8736
rect 9208 8676 9212 8732
rect 9212 8676 9268 8732
rect 9268 8676 9272 8732
rect 9208 8672 9272 8676
rect 9288 8732 9352 8736
rect 9288 8676 9292 8732
rect 9292 8676 9348 8732
rect 9348 8676 9352 8732
rect 9288 8672 9352 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 14605 8732 14669 8736
rect 14605 8676 14609 8732
rect 14609 8676 14665 8732
rect 14665 8676 14669 8732
rect 14605 8672 14669 8676
rect 14685 8732 14749 8736
rect 14685 8676 14689 8732
rect 14689 8676 14745 8732
rect 14745 8676 14749 8732
rect 14685 8672 14749 8676
rect 6349 8188 6413 8192
rect 6349 8132 6353 8188
rect 6353 8132 6409 8188
rect 6409 8132 6413 8188
rect 6349 8128 6413 8132
rect 6429 8188 6493 8192
rect 6429 8132 6433 8188
rect 6433 8132 6489 8188
rect 6489 8132 6493 8188
rect 6429 8128 6493 8132
rect 6509 8188 6573 8192
rect 6509 8132 6513 8188
rect 6513 8132 6569 8188
rect 6569 8132 6573 8188
rect 6509 8128 6573 8132
rect 6589 8188 6653 8192
rect 6589 8132 6593 8188
rect 6593 8132 6649 8188
rect 6649 8132 6653 8188
rect 6589 8128 6653 8132
rect 11746 8188 11810 8192
rect 11746 8132 11750 8188
rect 11750 8132 11806 8188
rect 11806 8132 11810 8188
rect 11746 8128 11810 8132
rect 11826 8188 11890 8192
rect 11826 8132 11830 8188
rect 11830 8132 11886 8188
rect 11886 8132 11890 8188
rect 11826 8128 11890 8132
rect 11906 8188 11970 8192
rect 11906 8132 11910 8188
rect 11910 8132 11966 8188
rect 11966 8132 11970 8188
rect 11906 8128 11970 8132
rect 11986 8188 12050 8192
rect 11986 8132 11990 8188
rect 11990 8132 12046 8188
rect 12046 8132 12050 8188
rect 11986 8128 12050 8132
rect 3650 7644 3714 7648
rect 3650 7588 3654 7644
rect 3654 7588 3710 7644
rect 3710 7588 3714 7644
rect 3650 7584 3714 7588
rect 3730 7644 3794 7648
rect 3730 7588 3734 7644
rect 3734 7588 3790 7644
rect 3790 7588 3794 7644
rect 3730 7584 3794 7588
rect 3810 7644 3874 7648
rect 3810 7588 3814 7644
rect 3814 7588 3870 7644
rect 3870 7588 3874 7644
rect 3810 7584 3874 7588
rect 3890 7644 3954 7648
rect 3890 7588 3894 7644
rect 3894 7588 3950 7644
rect 3950 7588 3954 7644
rect 3890 7584 3954 7588
rect 9048 7644 9112 7648
rect 9048 7588 9052 7644
rect 9052 7588 9108 7644
rect 9108 7588 9112 7644
rect 9048 7584 9112 7588
rect 9128 7644 9192 7648
rect 9128 7588 9132 7644
rect 9132 7588 9188 7644
rect 9188 7588 9192 7644
rect 9128 7584 9192 7588
rect 9208 7644 9272 7648
rect 9208 7588 9212 7644
rect 9212 7588 9268 7644
rect 9268 7588 9272 7644
rect 9208 7584 9272 7588
rect 9288 7644 9352 7648
rect 9288 7588 9292 7644
rect 9292 7588 9348 7644
rect 9348 7588 9352 7644
rect 9288 7584 9352 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 14605 7644 14669 7648
rect 14605 7588 14609 7644
rect 14609 7588 14665 7644
rect 14665 7588 14669 7644
rect 14605 7584 14669 7588
rect 14685 7644 14749 7648
rect 14685 7588 14689 7644
rect 14689 7588 14745 7644
rect 14745 7588 14749 7644
rect 14685 7584 14749 7588
rect 6349 7100 6413 7104
rect 6349 7044 6353 7100
rect 6353 7044 6409 7100
rect 6409 7044 6413 7100
rect 6349 7040 6413 7044
rect 6429 7100 6493 7104
rect 6429 7044 6433 7100
rect 6433 7044 6489 7100
rect 6489 7044 6493 7100
rect 6429 7040 6493 7044
rect 6509 7100 6573 7104
rect 6509 7044 6513 7100
rect 6513 7044 6569 7100
rect 6569 7044 6573 7100
rect 6509 7040 6573 7044
rect 6589 7100 6653 7104
rect 6589 7044 6593 7100
rect 6593 7044 6649 7100
rect 6649 7044 6653 7100
rect 6589 7040 6653 7044
rect 11746 7100 11810 7104
rect 11746 7044 11750 7100
rect 11750 7044 11806 7100
rect 11806 7044 11810 7100
rect 11746 7040 11810 7044
rect 11826 7100 11890 7104
rect 11826 7044 11830 7100
rect 11830 7044 11886 7100
rect 11886 7044 11890 7100
rect 11826 7040 11890 7044
rect 11906 7100 11970 7104
rect 11906 7044 11910 7100
rect 11910 7044 11966 7100
rect 11966 7044 11970 7100
rect 11906 7040 11970 7044
rect 11986 7100 12050 7104
rect 11986 7044 11990 7100
rect 11990 7044 12046 7100
rect 12046 7044 12050 7100
rect 11986 7040 12050 7044
rect 3650 6556 3714 6560
rect 3650 6500 3654 6556
rect 3654 6500 3710 6556
rect 3710 6500 3714 6556
rect 3650 6496 3714 6500
rect 3730 6556 3794 6560
rect 3730 6500 3734 6556
rect 3734 6500 3790 6556
rect 3790 6500 3794 6556
rect 3730 6496 3794 6500
rect 3810 6556 3874 6560
rect 3810 6500 3814 6556
rect 3814 6500 3870 6556
rect 3870 6500 3874 6556
rect 3810 6496 3874 6500
rect 3890 6556 3954 6560
rect 3890 6500 3894 6556
rect 3894 6500 3950 6556
rect 3950 6500 3954 6556
rect 3890 6496 3954 6500
rect 9048 6556 9112 6560
rect 9048 6500 9052 6556
rect 9052 6500 9108 6556
rect 9108 6500 9112 6556
rect 9048 6496 9112 6500
rect 9128 6556 9192 6560
rect 9128 6500 9132 6556
rect 9132 6500 9188 6556
rect 9188 6500 9192 6556
rect 9128 6496 9192 6500
rect 9208 6556 9272 6560
rect 9208 6500 9212 6556
rect 9212 6500 9268 6556
rect 9268 6500 9272 6556
rect 9208 6496 9272 6500
rect 9288 6556 9352 6560
rect 9288 6500 9292 6556
rect 9292 6500 9348 6556
rect 9348 6500 9352 6556
rect 9288 6496 9352 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 14605 6556 14669 6560
rect 14605 6500 14609 6556
rect 14609 6500 14665 6556
rect 14665 6500 14669 6556
rect 14605 6496 14669 6500
rect 14685 6556 14749 6560
rect 14685 6500 14689 6556
rect 14689 6500 14745 6556
rect 14745 6500 14749 6556
rect 14685 6496 14749 6500
rect 6349 6012 6413 6016
rect 6349 5956 6353 6012
rect 6353 5956 6409 6012
rect 6409 5956 6413 6012
rect 6349 5952 6413 5956
rect 6429 6012 6493 6016
rect 6429 5956 6433 6012
rect 6433 5956 6489 6012
rect 6489 5956 6493 6012
rect 6429 5952 6493 5956
rect 6509 6012 6573 6016
rect 6509 5956 6513 6012
rect 6513 5956 6569 6012
rect 6569 5956 6573 6012
rect 6509 5952 6573 5956
rect 6589 6012 6653 6016
rect 6589 5956 6593 6012
rect 6593 5956 6649 6012
rect 6649 5956 6653 6012
rect 6589 5952 6653 5956
rect 11746 6012 11810 6016
rect 11746 5956 11750 6012
rect 11750 5956 11806 6012
rect 11806 5956 11810 6012
rect 11746 5952 11810 5956
rect 11826 6012 11890 6016
rect 11826 5956 11830 6012
rect 11830 5956 11886 6012
rect 11886 5956 11890 6012
rect 11826 5952 11890 5956
rect 11906 6012 11970 6016
rect 11906 5956 11910 6012
rect 11910 5956 11966 6012
rect 11966 5956 11970 6012
rect 11906 5952 11970 5956
rect 11986 6012 12050 6016
rect 11986 5956 11990 6012
rect 11990 5956 12046 6012
rect 12046 5956 12050 6012
rect 11986 5952 12050 5956
rect 3650 5468 3714 5472
rect 3650 5412 3654 5468
rect 3654 5412 3710 5468
rect 3710 5412 3714 5468
rect 3650 5408 3714 5412
rect 3730 5468 3794 5472
rect 3730 5412 3734 5468
rect 3734 5412 3790 5468
rect 3790 5412 3794 5468
rect 3730 5408 3794 5412
rect 3810 5468 3874 5472
rect 3810 5412 3814 5468
rect 3814 5412 3870 5468
rect 3870 5412 3874 5468
rect 3810 5408 3874 5412
rect 3890 5468 3954 5472
rect 3890 5412 3894 5468
rect 3894 5412 3950 5468
rect 3950 5412 3954 5468
rect 3890 5408 3954 5412
rect 9048 5468 9112 5472
rect 9048 5412 9052 5468
rect 9052 5412 9108 5468
rect 9108 5412 9112 5468
rect 9048 5408 9112 5412
rect 9128 5468 9192 5472
rect 9128 5412 9132 5468
rect 9132 5412 9188 5468
rect 9188 5412 9192 5468
rect 9128 5408 9192 5412
rect 9208 5468 9272 5472
rect 9208 5412 9212 5468
rect 9212 5412 9268 5468
rect 9268 5412 9272 5468
rect 9208 5408 9272 5412
rect 9288 5468 9352 5472
rect 9288 5412 9292 5468
rect 9292 5412 9348 5468
rect 9348 5412 9352 5468
rect 9288 5408 9352 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 14605 5468 14669 5472
rect 14605 5412 14609 5468
rect 14609 5412 14665 5468
rect 14665 5412 14669 5468
rect 14605 5408 14669 5412
rect 14685 5468 14749 5472
rect 14685 5412 14689 5468
rect 14689 5412 14745 5468
rect 14745 5412 14749 5468
rect 14685 5408 14749 5412
rect 6349 4924 6413 4928
rect 6349 4868 6353 4924
rect 6353 4868 6409 4924
rect 6409 4868 6413 4924
rect 6349 4864 6413 4868
rect 6429 4924 6493 4928
rect 6429 4868 6433 4924
rect 6433 4868 6489 4924
rect 6489 4868 6493 4924
rect 6429 4864 6493 4868
rect 6509 4924 6573 4928
rect 6509 4868 6513 4924
rect 6513 4868 6569 4924
rect 6569 4868 6573 4924
rect 6509 4864 6573 4868
rect 6589 4924 6653 4928
rect 6589 4868 6593 4924
rect 6593 4868 6649 4924
rect 6649 4868 6653 4924
rect 6589 4864 6653 4868
rect 11746 4924 11810 4928
rect 11746 4868 11750 4924
rect 11750 4868 11806 4924
rect 11806 4868 11810 4924
rect 11746 4864 11810 4868
rect 11826 4924 11890 4928
rect 11826 4868 11830 4924
rect 11830 4868 11886 4924
rect 11886 4868 11890 4924
rect 11826 4864 11890 4868
rect 11906 4924 11970 4928
rect 11906 4868 11910 4924
rect 11910 4868 11966 4924
rect 11966 4868 11970 4924
rect 11906 4864 11970 4868
rect 11986 4924 12050 4928
rect 11986 4868 11990 4924
rect 11990 4868 12046 4924
rect 12046 4868 12050 4924
rect 11986 4864 12050 4868
rect 3650 4380 3714 4384
rect 3650 4324 3654 4380
rect 3654 4324 3710 4380
rect 3710 4324 3714 4380
rect 3650 4320 3714 4324
rect 3730 4380 3794 4384
rect 3730 4324 3734 4380
rect 3734 4324 3790 4380
rect 3790 4324 3794 4380
rect 3730 4320 3794 4324
rect 3810 4380 3874 4384
rect 3810 4324 3814 4380
rect 3814 4324 3870 4380
rect 3870 4324 3874 4380
rect 3810 4320 3874 4324
rect 3890 4380 3954 4384
rect 3890 4324 3894 4380
rect 3894 4324 3950 4380
rect 3950 4324 3954 4380
rect 3890 4320 3954 4324
rect 9048 4380 9112 4384
rect 9048 4324 9052 4380
rect 9052 4324 9108 4380
rect 9108 4324 9112 4380
rect 9048 4320 9112 4324
rect 9128 4380 9192 4384
rect 9128 4324 9132 4380
rect 9132 4324 9188 4380
rect 9188 4324 9192 4380
rect 9128 4320 9192 4324
rect 9208 4380 9272 4384
rect 9208 4324 9212 4380
rect 9212 4324 9268 4380
rect 9268 4324 9272 4380
rect 9208 4320 9272 4324
rect 9288 4380 9352 4384
rect 9288 4324 9292 4380
rect 9292 4324 9348 4380
rect 9348 4324 9352 4380
rect 9288 4320 9352 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 14605 4380 14669 4384
rect 14605 4324 14609 4380
rect 14609 4324 14665 4380
rect 14665 4324 14669 4380
rect 14605 4320 14669 4324
rect 14685 4380 14749 4384
rect 14685 4324 14689 4380
rect 14689 4324 14745 4380
rect 14745 4324 14749 4380
rect 14685 4320 14749 4324
rect 6349 3836 6413 3840
rect 6349 3780 6353 3836
rect 6353 3780 6409 3836
rect 6409 3780 6413 3836
rect 6349 3776 6413 3780
rect 6429 3836 6493 3840
rect 6429 3780 6433 3836
rect 6433 3780 6489 3836
rect 6489 3780 6493 3836
rect 6429 3776 6493 3780
rect 6509 3836 6573 3840
rect 6509 3780 6513 3836
rect 6513 3780 6569 3836
rect 6569 3780 6573 3836
rect 6509 3776 6573 3780
rect 6589 3836 6653 3840
rect 6589 3780 6593 3836
rect 6593 3780 6649 3836
rect 6649 3780 6653 3836
rect 6589 3776 6653 3780
rect 11746 3836 11810 3840
rect 11746 3780 11750 3836
rect 11750 3780 11806 3836
rect 11806 3780 11810 3836
rect 11746 3776 11810 3780
rect 11826 3836 11890 3840
rect 11826 3780 11830 3836
rect 11830 3780 11886 3836
rect 11886 3780 11890 3836
rect 11826 3776 11890 3780
rect 11906 3836 11970 3840
rect 11906 3780 11910 3836
rect 11910 3780 11966 3836
rect 11966 3780 11970 3836
rect 11906 3776 11970 3780
rect 11986 3836 12050 3840
rect 11986 3780 11990 3836
rect 11990 3780 12046 3836
rect 12046 3780 12050 3836
rect 11986 3776 12050 3780
rect 3650 3292 3714 3296
rect 3650 3236 3654 3292
rect 3654 3236 3710 3292
rect 3710 3236 3714 3292
rect 3650 3232 3714 3236
rect 3730 3292 3794 3296
rect 3730 3236 3734 3292
rect 3734 3236 3790 3292
rect 3790 3236 3794 3292
rect 3730 3232 3794 3236
rect 3810 3292 3874 3296
rect 3810 3236 3814 3292
rect 3814 3236 3870 3292
rect 3870 3236 3874 3292
rect 3810 3232 3874 3236
rect 3890 3292 3954 3296
rect 3890 3236 3894 3292
rect 3894 3236 3950 3292
rect 3950 3236 3954 3292
rect 3890 3232 3954 3236
rect 9048 3292 9112 3296
rect 9048 3236 9052 3292
rect 9052 3236 9108 3292
rect 9108 3236 9112 3292
rect 9048 3232 9112 3236
rect 9128 3292 9192 3296
rect 9128 3236 9132 3292
rect 9132 3236 9188 3292
rect 9188 3236 9192 3292
rect 9128 3232 9192 3236
rect 9208 3292 9272 3296
rect 9208 3236 9212 3292
rect 9212 3236 9268 3292
rect 9268 3236 9272 3292
rect 9208 3232 9272 3236
rect 9288 3292 9352 3296
rect 9288 3236 9292 3292
rect 9292 3236 9348 3292
rect 9348 3236 9352 3292
rect 9288 3232 9352 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 14605 3292 14669 3296
rect 14605 3236 14609 3292
rect 14609 3236 14665 3292
rect 14665 3236 14669 3292
rect 14605 3232 14669 3236
rect 14685 3292 14749 3296
rect 14685 3236 14689 3292
rect 14689 3236 14745 3292
rect 14745 3236 14749 3292
rect 14685 3232 14749 3236
rect 6349 2748 6413 2752
rect 6349 2692 6353 2748
rect 6353 2692 6409 2748
rect 6409 2692 6413 2748
rect 6349 2688 6413 2692
rect 6429 2748 6493 2752
rect 6429 2692 6433 2748
rect 6433 2692 6489 2748
rect 6489 2692 6493 2748
rect 6429 2688 6493 2692
rect 6509 2748 6573 2752
rect 6509 2692 6513 2748
rect 6513 2692 6569 2748
rect 6569 2692 6573 2748
rect 6509 2688 6573 2692
rect 6589 2748 6653 2752
rect 6589 2692 6593 2748
rect 6593 2692 6649 2748
rect 6649 2692 6653 2748
rect 6589 2688 6653 2692
rect 11746 2748 11810 2752
rect 11746 2692 11750 2748
rect 11750 2692 11806 2748
rect 11806 2692 11810 2748
rect 11746 2688 11810 2692
rect 11826 2748 11890 2752
rect 11826 2692 11830 2748
rect 11830 2692 11886 2748
rect 11886 2692 11890 2748
rect 11826 2688 11890 2692
rect 11906 2748 11970 2752
rect 11906 2692 11910 2748
rect 11910 2692 11966 2748
rect 11966 2692 11970 2748
rect 11906 2688 11970 2692
rect 11986 2748 12050 2752
rect 11986 2692 11990 2748
rect 11990 2692 12046 2748
rect 12046 2692 12050 2748
rect 11986 2688 12050 2692
rect 3650 2204 3714 2208
rect 3650 2148 3654 2204
rect 3654 2148 3710 2204
rect 3710 2148 3714 2204
rect 3650 2144 3714 2148
rect 3730 2204 3794 2208
rect 3730 2148 3734 2204
rect 3734 2148 3790 2204
rect 3790 2148 3794 2204
rect 3730 2144 3794 2148
rect 3810 2204 3874 2208
rect 3810 2148 3814 2204
rect 3814 2148 3870 2204
rect 3870 2148 3874 2204
rect 3810 2144 3874 2148
rect 3890 2204 3954 2208
rect 3890 2148 3894 2204
rect 3894 2148 3950 2204
rect 3950 2148 3954 2204
rect 3890 2144 3954 2148
rect 9048 2204 9112 2208
rect 9048 2148 9052 2204
rect 9052 2148 9108 2204
rect 9108 2148 9112 2204
rect 9048 2144 9112 2148
rect 9128 2204 9192 2208
rect 9128 2148 9132 2204
rect 9132 2148 9188 2204
rect 9188 2148 9192 2204
rect 9128 2144 9192 2148
rect 9208 2204 9272 2208
rect 9208 2148 9212 2204
rect 9212 2148 9268 2204
rect 9268 2148 9272 2204
rect 9208 2144 9272 2148
rect 9288 2204 9352 2208
rect 9288 2148 9292 2204
rect 9292 2148 9348 2204
rect 9348 2148 9352 2204
rect 9288 2144 9352 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
rect 14605 2204 14669 2208
rect 14605 2148 14609 2204
rect 14609 2148 14665 2204
rect 14665 2148 14669 2204
rect 14605 2144 14669 2148
rect 14685 2204 14749 2208
rect 14685 2148 14689 2204
rect 14689 2148 14745 2204
rect 14745 2148 14749 2204
rect 14685 2144 14749 2148
<< metal4 >>
rect -916 19930 -596 19972
rect -916 19694 -874 19930
rect -638 19694 -596 19930
rect -916 12763 -596 19694
rect -916 12527 -874 12763
rect -638 12527 -596 12763
rect -916 7504 -596 12527
rect -916 7268 -874 7504
rect -638 7268 -596 7504
rect -916 434 -596 7268
rect -256 19270 64 19312
rect -256 19034 -214 19270
rect 22 19034 64 19270
rect -256 15392 64 19034
rect -256 15156 -214 15392
rect 22 15156 64 15392
rect -256 10134 64 15156
rect -256 9898 -214 10134
rect 22 9898 64 10134
rect -256 4875 64 9898
rect -256 4639 -214 4875
rect 22 4639 64 4875
rect -256 1094 64 4639
rect -256 858 -214 1094
rect 22 858 64 1094
rect -256 816 64 858
rect 3642 19270 3963 19972
rect 3642 19034 3684 19270
rect 3920 19034 3963 19270
rect 3642 17440 3963 19034
rect 3642 17376 3650 17440
rect 3714 17376 3730 17440
rect 3794 17376 3810 17440
rect 3874 17376 3890 17440
rect 3954 17376 3963 17440
rect 3642 16352 3963 17376
rect 3642 16288 3650 16352
rect 3714 16288 3730 16352
rect 3794 16288 3810 16352
rect 3874 16288 3890 16352
rect 3954 16288 3963 16352
rect 3642 15392 3963 16288
rect 3642 15264 3684 15392
rect 3920 15264 3963 15392
rect 3642 15200 3650 15264
rect 3954 15200 3963 15264
rect 3642 15156 3684 15200
rect 3920 15156 3963 15200
rect 3642 14176 3963 15156
rect 3642 14112 3650 14176
rect 3714 14112 3730 14176
rect 3794 14112 3810 14176
rect 3874 14112 3890 14176
rect 3954 14112 3963 14176
rect 3642 13088 3963 14112
rect 3642 13024 3650 13088
rect 3714 13024 3730 13088
rect 3794 13024 3810 13088
rect 3874 13024 3890 13088
rect 3954 13024 3963 13088
rect 3642 12000 3963 13024
rect 3642 11936 3650 12000
rect 3714 11936 3730 12000
rect 3794 11936 3810 12000
rect 3874 11936 3890 12000
rect 3954 11936 3963 12000
rect 3642 10912 3963 11936
rect 3642 10848 3650 10912
rect 3714 10848 3730 10912
rect 3794 10848 3810 10912
rect 3874 10848 3890 10912
rect 3954 10848 3963 10912
rect 3642 10134 3963 10848
rect 3642 9898 3684 10134
rect 3920 9898 3963 10134
rect 3642 9824 3963 9898
rect 3642 9760 3650 9824
rect 3714 9760 3730 9824
rect 3794 9760 3810 9824
rect 3874 9760 3890 9824
rect 3954 9760 3963 9824
rect 3642 8736 3963 9760
rect 3642 8672 3650 8736
rect 3714 8672 3730 8736
rect 3794 8672 3810 8736
rect 3874 8672 3890 8736
rect 3954 8672 3963 8736
rect 3642 7648 3963 8672
rect 3642 7584 3650 7648
rect 3714 7584 3730 7648
rect 3794 7584 3810 7648
rect 3874 7584 3890 7648
rect 3954 7584 3963 7648
rect 3642 6560 3963 7584
rect 3642 6496 3650 6560
rect 3714 6496 3730 6560
rect 3794 6496 3810 6560
rect 3874 6496 3890 6560
rect 3954 6496 3963 6560
rect 3642 5472 3963 6496
rect 3642 5408 3650 5472
rect 3714 5408 3730 5472
rect 3794 5408 3810 5472
rect 3874 5408 3890 5472
rect 3954 5408 3963 5472
rect 3642 4875 3963 5408
rect 3642 4639 3684 4875
rect 3920 4639 3963 4875
rect 3642 4384 3963 4639
rect 3642 4320 3650 4384
rect 3714 4320 3730 4384
rect 3794 4320 3810 4384
rect 3874 4320 3890 4384
rect 3954 4320 3963 4384
rect 3642 3296 3963 4320
rect 3642 3232 3650 3296
rect 3714 3232 3730 3296
rect 3794 3232 3810 3296
rect 3874 3232 3890 3296
rect 3954 3232 3963 3296
rect 3642 2208 3963 3232
rect 3642 2144 3650 2208
rect 3714 2144 3730 2208
rect 3794 2144 3810 2208
rect 3874 2144 3890 2208
rect 3954 2144 3963 2208
rect 3642 1094 3963 2144
rect 3642 858 3684 1094
rect 3920 858 3963 1094
rect -916 198 -874 434
rect -638 198 -596 434
rect -916 156 -596 198
rect 3642 156 3963 858
rect 6341 19930 6661 19972
rect 6341 19694 6383 19930
rect 6619 19694 6661 19930
rect 6341 17984 6661 19694
rect 6341 17920 6349 17984
rect 6413 17920 6429 17984
rect 6493 17920 6509 17984
rect 6573 17920 6589 17984
rect 6653 17920 6661 17984
rect 6341 16896 6661 17920
rect 6341 16832 6349 16896
rect 6413 16832 6429 16896
rect 6493 16832 6509 16896
rect 6573 16832 6589 16896
rect 6653 16832 6661 16896
rect 6341 15808 6661 16832
rect 6341 15744 6349 15808
rect 6413 15744 6429 15808
rect 6493 15744 6509 15808
rect 6573 15744 6589 15808
rect 6653 15744 6661 15808
rect 6341 14720 6661 15744
rect 6341 14656 6349 14720
rect 6413 14656 6429 14720
rect 6493 14656 6509 14720
rect 6573 14656 6589 14720
rect 6653 14656 6661 14720
rect 6341 13632 6661 14656
rect 6341 13568 6349 13632
rect 6413 13568 6429 13632
rect 6493 13568 6509 13632
rect 6573 13568 6589 13632
rect 6653 13568 6661 13632
rect 6341 12763 6661 13568
rect 6341 12544 6383 12763
rect 6619 12544 6661 12763
rect 6341 12480 6349 12544
rect 6413 12480 6429 12527
rect 6493 12480 6509 12527
rect 6573 12480 6589 12527
rect 6653 12480 6661 12544
rect 6341 11456 6661 12480
rect 6341 11392 6349 11456
rect 6413 11392 6429 11456
rect 6493 11392 6509 11456
rect 6573 11392 6589 11456
rect 6653 11392 6661 11456
rect 6341 10368 6661 11392
rect 6341 10304 6349 10368
rect 6413 10304 6429 10368
rect 6493 10304 6509 10368
rect 6573 10304 6589 10368
rect 6653 10304 6661 10368
rect 6341 9280 6661 10304
rect 6341 9216 6349 9280
rect 6413 9216 6429 9280
rect 6493 9216 6509 9280
rect 6573 9216 6589 9280
rect 6653 9216 6661 9280
rect 6341 8192 6661 9216
rect 6341 8128 6349 8192
rect 6413 8128 6429 8192
rect 6493 8128 6509 8192
rect 6573 8128 6589 8192
rect 6653 8128 6661 8192
rect 6341 7504 6661 8128
rect 6341 7268 6383 7504
rect 6619 7268 6661 7504
rect 6341 7104 6661 7268
rect 6341 7040 6349 7104
rect 6413 7040 6429 7104
rect 6493 7040 6509 7104
rect 6573 7040 6589 7104
rect 6653 7040 6661 7104
rect 6341 6016 6661 7040
rect 6341 5952 6349 6016
rect 6413 5952 6429 6016
rect 6493 5952 6509 6016
rect 6573 5952 6589 6016
rect 6653 5952 6661 6016
rect 6341 4928 6661 5952
rect 6341 4864 6349 4928
rect 6413 4864 6429 4928
rect 6493 4864 6509 4928
rect 6573 4864 6589 4928
rect 6653 4864 6661 4928
rect 6341 3840 6661 4864
rect 6341 3776 6349 3840
rect 6413 3776 6429 3840
rect 6493 3776 6509 3840
rect 6573 3776 6589 3840
rect 6653 3776 6661 3840
rect 6341 2752 6661 3776
rect 6341 2688 6349 2752
rect 6413 2688 6429 2752
rect 6493 2688 6509 2752
rect 6573 2688 6589 2752
rect 6653 2688 6661 2752
rect 6341 434 6661 2688
rect 6341 198 6383 434
rect 6619 198 6661 434
rect 6341 156 6661 198
rect 9040 19270 9360 19972
rect 9040 19034 9082 19270
rect 9318 19034 9360 19270
rect 9040 17440 9360 19034
rect 9040 17376 9048 17440
rect 9112 17376 9128 17440
rect 9192 17376 9208 17440
rect 9272 17376 9288 17440
rect 9352 17376 9360 17440
rect 9040 16352 9360 17376
rect 9040 16288 9048 16352
rect 9112 16288 9128 16352
rect 9192 16288 9208 16352
rect 9272 16288 9288 16352
rect 9352 16288 9360 16352
rect 9040 15392 9360 16288
rect 9040 15264 9082 15392
rect 9318 15264 9360 15392
rect 9040 15200 9048 15264
rect 9352 15200 9360 15264
rect 9040 15156 9082 15200
rect 9318 15156 9360 15200
rect 9040 14176 9360 15156
rect 9040 14112 9048 14176
rect 9112 14112 9128 14176
rect 9192 14112 9208 14176
rect 9272 14112 9288 14176
rect 9352 14112 9360 14176
rect 9040 13088 9360 14112
rect 9040 13024 9048 13088
rect 9112 13024 9128 13088
rect 9192 13024 9208 13088
rect 9272 13024 9288 13088
rect 9352 13024 9360 13088
rect 9040 12000 9360 13024
rect 9040 11936 9048 12000
rect 9112 11936 9128 12000
rect 9192 11936 9208 12000
rect 9272 11936 9288 12000
rect 9352 11936 9360 12000
rect 9040 10912 9360 11936
rect 9040 10848 9048 10912
rect 9112 10848 9128 10912
rect 9192 10848 9208 10912
rect 9272 10848 9288 10912
rect 9352 10848 9360 10912
rect 9040 10134 9360 10848
rect 9040 9898 9082 10134
rect 9318 9898 9360 10134
rect 9040 9824 9360 9898
rect 9040 9760 9048 9824
rect 9112 9760 9128 9824
rect 9192 9760 9208 9824
rect 9272 9760 9288 9824
rect 9352 9760 9360 9824
rect 9040 8736 9360 9760
rect 9040 8672 9048 8736
rect 9112 8672 9128 8736
rect 9192 8672 9208 8736
rect 9272 8672 9288 8736
rect 9352 8672 9360 8736
rect 9040 7648 9360 8672
rect 9040 7584 9048 7648
rect 9112 7584 9128 7648
rect 9192 7584 9208 7648
rect 9272 7584 9288 7648
rect 9352 7584 9360 7648
rect 9040 6560 9360 7584
rect 9040 6496 9048 6560
rect 9112 6496 9128 6560
rect 9192 6496 9208 6560
rect 9272 6496 9288 6560
rect 9352 6496 9360 6560
rect 9040 5472 9360 6496
rect 9040 5408 9048 5472
rect 9112 5408 9128 5472
rect 9192 5408 9208 5472
rect 9272 5408 9288 5472
rect 9352 5408 9360 5472
rect 9040 4875 9360 5408
rect 9040 4639 9082 4875
rect 9318 4639 9360 4875
rect 9040 4384 9360 4639
rect 9040 4320 9048 4384
rect 9112 4320 9128 4384
rect 9192 4320 9208 4384
rect 9272 4320 9288 4384
rect 9352 4320 9360 4384
rect 9040 3296 9360 4320
rect 9040 3232 9048 3296
rect 9112 3232 9128 3296
rect 9192 3232 9208 3296
rect 9272 3232 9288 3296
rect 9352 3232 9360 3296
rect 9040 2208 9360 3232
rect 9040 2144 9048 2208
rect 9112 2144 9128 2208
rect 9192 2144 9208 2208
rect 9272 2144 9288 2208
rect 9352 2144 9360 2208
rect 9040 1094 9360 2144
rect 9040 858 9082 1094
rect 9318 858 9360 1094
rect 9040 156 9360 858
rect 11738 19930 12059 19972
rect 11738 19694 11780 19930
rect 12016 19694 12059 19930
rect 11738 17984 12059 19694
rect 11738 17920 11746 17984
rect 11810 17920 11826 17984
rect 11890 17920 11906 17984
rect 11970 17920 11986 17984
rect 12050 17920 12059 17984
rect 11738 16896 12059 17920
rect 11738 16832 11746 16896
rect 11810 16832 11826 16896
rect 11890 16832 11906 16896
rect 11970 16832 11986 16896
rect 12050 16832 12059 16896
rect 11738 15808 12059 16832
rect 11738 15744 11746 15808
rect 11810 15744 11826 15808
rect 11890 15744 11906 15808
rect 11970 15744 11986 15808
rect 12050 15744 12059 15808
rect 11738 14720 12059 15744
rect 11738 14656 11746 14720
rect 11810 14656 11826 14720
rect 11890 14656 11906 14720
rect 11970 14656 11986 14720
rect 12050 14656 12059 14720
rect 11738 13632 12059 14656
rect 11738 13568 11746 13632
rect 11810 13568 11826 13632
rect 11890 13568 11906 13632
rect 11970 13568 11986 13632
rect 12050 13568 12059 13632
rect 11738 12763 12059 13568
rect 11738 12544 11780 12763
rect 12016 12544 12059 12763
rect 11738 12480 11746 12544
rect 11810 12480 11826 12527
rect 11890 12480 11906 12527
rect 11970 12480 11986 12527
rect 12050 12480 12059 12544
rect 11738 11456 12059 12480
rect 11738 11392 11746 11456
rect 11810 11392 11826 11456
rect 11890 11392 11906 11456
rect 11970 11392 11986 11456
rect 12050 11392 12059 11456
rect 11738 10368 12059 11392
rect 11738 10304 11746 10368
rect 11810 10304 11826 10368
rect 11890 10304 11906 10368
rect 11970 10304 11986 10368
rect 12050 10304 12059 10368
rect 11738 9280 12059 10304
rect 11738 9216 11746 9280
rect 11810 9216 11826 9280
rect 11890 9216 11906 9280
rect 11970 9216 11986 9280
rect 12050 9216 12059 9280
rect 11738 8192 12059 9216
rect 11738 8128 11746 8192
rect 11810 8128 11826 8192
rect 11890 8128 11906 8192
rect 11970 8128 11986 8192
rect 12050 8128 12059 8192
rect 11738 7504 12059 8128
rect 11738 7268 11780 7504
rect 12016 7268 12059 7504
rect 11738 7104 12059 7268
rect 11738 7040 11746 7104
rect 11810 7040 11826 7104
rect 11890 7040 11906 7104
rect 11970 7040 11986 7104
rect 12050 7040 12059 7104
rect 11738 6016 12059 7040
rect 11738 5952 11746 6016
rect 11810 5952 11826 6016
rect 11890 5952 11906 6016
rect 11970 5952 11986 6016
rect 12050 5952 12059 6016
rect 11738 4928 12059 5952
rect 11738 4864 11746 4928
rect 11810 4864 11826 4928
rect 11890 4864 11906 4928
rect 11970 4864 11986 4928
rect 12050 4864 12059 4928
rect 11738 3840 12059 4864
rect 11738 3776 11746 3840
rect 11810 3776 11826 3840
rect 11890 3776 11906 3840
rect 11970 3776 11986 3840
rect 12050 3776 12059 3840
rect 11738 2752 12059 3776
rect 11738 2688 11746 2752
rect 11810 2688 11826 2752
rect 11890 2688 11906 2752
rect 11970 2688 11986 2752
rect 12050 2688 12059 2752
rect 11738 434 12059 2688
rect 11738 198 11780 434
rect 12016 198 12059 434
rect 11738 156 12059 198
rect 14437 19270 14757 19972
rect 18996 19930 19316 19972
rect 18996 19694 19038 19930
rect 19274 19694 19316 19930
rect 14437 19034 14479 19270
rect 14715 19034 14757 19270
rect 14437 17440 14757 19034
rect 14437 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14605 17440
rect 14669 17376 14685 17440
rect 14749 17376 14757 17440
rect 14437 16352 14757 17376
rect 14437 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14605 16352
rect 14669 16288 14685 16352
rect 14749 16288 14757 16352
rect 14437 15392 14757 16288
rect 14437 15264 14479 15392
rect 14715 15264 14757 15392
rect 14437 15200 14445 15264
rect 14749 15200 14757 15264
rect 14437 15156 14479 15200
rect 14715 15156 14757 15200
rect 14437 14176 14757 15156
rect 14437 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14605 14176
rect 14669 14112 14685 14176
rect 14749 14112 14757 14176
rect 14437 13088 14757 14112
rect 14437 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14605 13088
rect 14669 13024 14685 13088
rect 14749 13024 14757 13088
rect 14437 12000 14757 13024
rect 14437 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14605 12000
rect 14669 11936 14685 12000
rect 14749 11936 14757 12000
rect 14437 10912 14757 11936
rect 14437 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14605 10912
rect 14669 10848 14685 10912
rect 14749 10848 14757 10912
rect 14437 10134 14757 10848
rect 14437 9898 14479 10134
rect 14715 9898 14757 10134
rect 14437 9824 14757 9898
rect 14437 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14605 9824
rect 14669 9760 14685 9824
rect 14749 9760 14757 9824
rect 14437 8736 14757 9760
rect 14437 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14605 8736
rect 14669 8672 14685 8736
rect 14749 8672 14757 8736
rect 14437 7648 14757 8672
rect 14437 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14605 7648
rect 14669 7584 14685 7648
rect 14749 7584 14757 7648
rect 14437 6560 14757 7584
rect 14437 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14605 6560
rect 14669 6496 14685 6560
rect 14749 6496 14757 6560
rect 14437 5472 14757 6496
rect 14437 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14605 5472
rect 14669 5408 14685 5472
rect 14749 5408 14757 5472
rect 14437 4875 14757 5408
rect 14437 4639 14479 4875
rect 14715 4639 14757 4875
rect 14437 4384 14757 4639
rect 14437 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14605 4384
rect 14669 4320 14685 4384
rect 14749 4320 14757 4384
rect 14437 3296 14757 4320
rect 14437 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14605 3296
rect 14669 3232 14685 3296
rect 14749 3232 14757 3296
rect 14437 2208 14757 3232
rect 14437 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14605 2208
rect 14669 2144 14685 2208
rect 14749 2144 14757 2208
rect 14437 1094 14757 2144
rect 14437 858 14479 1094
rect 14715 858 14757 1094
rect 14437 156 14757 858
rect 18336 19270 18656 19312
rect 18336 19034 18378 19270
rect 18614 19034 18656 19270
rect 18336 15392 18656 19034
rect 18336 15156 18378 15392
rect 18614 15156 18656 15392
rect 18336 10134 18656 15156
rect 18336 9898 18378 10134
rect 18614 9898 18656 10134
rect 18336 4875 18656 9898
rect 18336 4639 18378 4875
rect 18614 4639 18656 4875
rect 18336 1094 18656 4639
rect 18336 858 18378 1094
rect 18614 858 18656 1094
rect 18336 816 18656 858
rect 18996 12763 19316 19694
rect 18996 12527 19038 12763
rect 19274 12527 19316 12763
rect 18996 7504 19316 12527
rect 18996 7268 19038 7504
rect 19274 7268 19316 7504
rect 18996 434 19316 7268
rect 18996 198 19038 434
rect 19274 198 19316 434
rect 18996 156 19316 198
<< via4 >>
rect -874 19694 -638 19930
rect -874 12527 -638 12763
rect -874 7268 -638 7504
rect -214 19034 22 19270
rect -214 15156 22 15392
rect -214 9898 22 10134
rect -214 4639 22 4875
rect -214 858 22 1094
rect 3684 19034 3920 19270
rect 3684 15264 3920 15392
rect 3684 15200 3714 15264
rect 3714 15200 3730 15264
rect 3730 15200 3794 15264
rect 3794 15200 3810 15264
rect 3810 15200 3874 15264
rect 3874 15200 3890 15264
rect 3890 15200 3920 15264
rect 3684 15156 3920 15200
rect 3684 9898 3920 10134
rect 3684 4639 3920 4875
rect 3684 858 3920 1094
rect -874 198 -638 434
rect 6383 19694 6619 19930
rect 6383 12544 6619 12763
rect 6383 12527 6413 12544
rect 6413 12527 6429 12544
rect 6429 12527 6493 12544
rect 6493 12527 6509 12544
rect 6509 12527 6573 12544
rect 6573 12527 6589 12544
rect 6589 12527 6619 12544
rect 6383 7268 6619 7504
rect 6383 198 6619 434
rect 9082 19034 9318 19270
rect 9082 15264 9318 15392
rect 9082 15200 9112 15264
rect 9112 15200 9128 15264
rect 9128 15200 9192 15264
rect 9192 15200 9208 15264
rect 9208 15200 9272 15264
rect 9272 15200 9288 15264
rect 9288 15200 9318 15264
rect 9082 15156 9318 15200
rect 9082 9898 9318 10134
rect 9082 4639 9318 4875
rect 9082 858 9318 1094
rect 11780 19694 12016 19930
rect 11780 12544 12016 12763
rect 11780 12527 11810 12544
rect 11810 12527 11826 12544
rect 11826 12527 11890 12544
rect 11890 12527 11906 12544
rect 11906 12527 11970 12544
rect 11970 12527 11986 12544
rect 11986 12527 12016 12544
rect 11780 7268 12016 7504
rect 11780 198 12016 434
rect 19038 19694 19274 19930
rect 14479 19034 14715 19270
rect 14479 15264 14715 15392
rect 14479 15200 14509 15264
rect 14509 15200 14525 15264
rect 14525 15200 14589 15264
rect 14589 15200 14605 15264
rect 14605 15200 14669 15264
rect 14669 15200 14685 15264
rect 14685 15200 14715 15264
rect 14479 15156 14715 15200
rect 14479 9898 14715 10134
rect 14479 4639 14715 4875
rect 14479 858 14715 1094
rect 18378 19034 18614 19270
rect 18378 15156 18614 15392
rect 18378 9898 18614 10134
rect 18378 4639 18614 4875
rect 18378 858 18614 1094
rect 19038 12527 19274 12763
rect 19038 7268 19274 7504
rect 19038 198 19274 434
<< metal5 >>
rect -916 19930 19316 19972
rect -916 19694 -874 19930
rect -638 19694 6383 19930
rect 6619 19694 11780 19930
rect 12016 19694 19038 19930
rect 19274 19694 19316 19930
rect -916 19652 19316 19694
rect -256 19270 18656 19312
rect -256 19034 -214 19270
rect 22 19034 3684 19270
rect 3920 19034 9082 19270
rect 9318 19034 14479 19270
rect 14715 19034 18378 19270
rect 18614 19034 18656 19270
rect -256 18992 18656 19034
rect -916 15392 19316 15435
rect -916 15156 -214 15392
rect 22 15156 3684 15392
rect 3920 15156 9082 15392
rect 9318 15156 14479 15392
rect 14715 15156 18378 15392
rect 18614 15156 19316 15392
rect -916 15114 19316 15156
rect -916 12763 19316 12805
rect -916 12527 -874 12763
rect -638 12527 6383 12763
rect 6619 12527 11780 12763
rect 12016 12527 19038 12763
rect 19274 12527 19316 12763
rect -916 12485 19316 12527
rect -916 10134 19316 10176
rect -916 9898 -214 10134
rect 22 9898 3684 10134
rect 3920 9898 9082 10134
rect 9318 9898 14479 10134
rect 14715 9898 18378 10134
rect 18614 9898 19316 10134
rect -916 9856 19316 9898
rect -916 7504 19316 7547
rect -916 7268 -874 7504
rect -638 7268 6383 7504
rect 6619 7268 11780 7504
rect 12016 7268 19038 7504
rect 19274 7268 19316 7504
rect -916 7226 19316 7268
rect -916 4875 19316 4917
rect -916 4639 -214 4875
rect 22 4639 3684 4875
rect 3920 4639 9082 4875
rect 9318 4639 14479 4875
rect 14715 4639 18378 4875
rect 18614 4639 19316 4875
rect -916 4597 19316 4639
rect -256 1094 18656 1136
rect -256 858 -214 1094
rect 22 858 3684 1094
rect 3920 858 9082 1094
rect 9318 858 14479 1094
rect 14715 858 18378 1094
rect 18614 858 18656 1094
rect -256 816 18656 858
rect -916 434 19316 476
rect -916 198 -874 434
rect -638 198 6383 434
rect 6619 198 11780 434
rect 12016 198 19038 434
rect 19274 198 19316 434
rect -916 156 19316 198
use sky130_fd_sc_hd__decap_6  FILLER_1_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 1932 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1618419204
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1618419204
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ringosc.ibufp11
timestamp 1619507013
transform -1 0 1932 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1619507013
transform -1 0 2392 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 3036 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14
timestamp 1618419204
transform 1 0 2392 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 2760 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfrbp_2  idiv2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 2484 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_4  irb
timestamp 1619507013
transform -1 0 5244 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 5336 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1618419204
transform 1 0 4140 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30
timestamp 1618419204
transform 1 0 3864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36
timestamp 1618419204
transform 1 0 4416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45
timestamp 1618419204
transform 1 0 5244 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_39
timestamp 1618419204
transform 1 0 4692 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1618419204
transform 1 0 5336 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_58
timestamp 1618419204
transform 1 0 6440 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_53
timestamp 1618419204
transform 1 0 5980 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 6532 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1618419204
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1618419204
transform 1 0 6624 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1618419204
transform -1 0 6072 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1618419204
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1618419204
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1618419204
transform -1 0 5980 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_73
timestamp 1618419204
transform 1 0 7820 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1618419204
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[11\].id.delayenb1
timestamp 1619507013
transform -1 0 7912 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_4  ringosc.dstage\[11\].id.delayen0
timestamp 1619507013
transform 1 0 6808 0 1 2720
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74
timestamp 1618419204
transform 1 0 7912 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_82
timestamp 1618419204
transform 1 0 8648 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1618419204
transform 1 0 8280 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _355_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 8372 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_88
timestamp 1618419204
transform 1 0 9200 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1618419204
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86
timestamp 1618419204
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1618419204
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 9568 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp 1618419204
transform 1 0 9568 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1618419204
transform 1 0 10028 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_101
timestamp 1618419204
transform 1 0 10396 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_108
timestamp 1618419204
transform 1 0 11040 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb0
timestamp 1619507013
transform -1 0 11040 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen0
timestamp 1618419204
transform -1 0 11224 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_1_115
timestamp 1618419204
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1618419204
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117
timestamp 1618419204
transform 1 0 11868 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1618419204
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1618419204
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_2  _323_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 12788 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  input1
timestamp 1619507013
transform 1 0 12420 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_127
timestamp 1618419204
transform 1 0 12788 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_136
timestamp 1618419204
transform 1 0 13616 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_132
timestamp 1618419204
transform 1 0 13248 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1618419204
transform 1 0 13156 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_140
timestamp 1618419204
transform 1 0 13984 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1618419204
transform 1 0 14536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1618419204
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1618419204
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1618419204
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfrbp_1  idiv16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 14352 0 1 2720
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_0_150
timestamp 1618419204
transform 1 0 14904 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1618419204
transform 1 0 14996 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_154
timestamp 1618419204
transform 1 0 15272 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1619507013
transform -1 0 15916 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_161
timestamp 1618419204
transform 1 0 15916 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_167
timestamp 1618419204
transform 1 0 16468 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output43
timestamp 1618419204
transform 1 0 16284 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_172
timestamp 1618419204
transform 1 0 16928 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1618419204
transform 1 0 16652 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1618419204
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1618419204
transform -1 0 17296 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1618419204
transform -1 0 17296 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1618419204
transform 1 0 3036 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  ringosc.ibufp10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 2484 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1618419204
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1618419204
transform -1 0 1840 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_8
timestamp 1618419204
transform 1 0 1840 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_15
timestamp 1618419204
transform 1 0 2484 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfrbp_2  idiv4
timestamp 1618419204
transform -1 0 6440 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1618419204
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_25
timestamp 1618419204
transform 1 0 3404 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_30
timestamp 1618419204
transform 1 0 3864 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb0
timestamp 1619507013
transform 1 0 6808 0 -1 3808
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_2_58
timestamp 1618419204
transform 1 0 6440 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1618419204
transform 1 0 7820 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[11\].id.delayen1
timestamp 1618419204
transform 1 0 8188 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb1
timestamp 1619507013
transform 1 0 9476 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1618419204
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_82
timestamp 1618419204
transform 1 0 8648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1618419204
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_98
timestamp 1618419204
transform 1 0 10120 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1618419204
transform 1 0 12420 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1618419204
transform 1 0 10948 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_106
timestamp 1618419204
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_116
timestamp 1618419204
transform 1 0 11776 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_122
timestamp 1618419204
transform 1 0 12328 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1619507013
transform 1 0 13616 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1618419204
transform 1 0 14720 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1618419204
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_132
timestamp 1618419204
transform 1 0 13248 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_139
timestamp 1618419204
transform 1 0 13892 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_144
timestamp 1618419204
transform 1 0 14352 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _325_
timestamp 1618419204
transform 1 0 15916 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1618419204
transform -1 0 17296 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_157
timestamp 1618419204
transform 1 0 15548 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_169
timestamp 1618419204
transform 1 0 16652 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1618419204
transform 1 0 2576 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1618419204
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output41
timestamp 1618419204
transform -1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_7
timestamp 1618419204
transform 1 0 1748 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_15
timestamp 1618419204
transform 1 0 2484 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_19
timestamp 1618419204
transform 1 0 2852 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 3680 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 5704 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_3_27
timestamp 1618419204
transform 1 0 3588 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_41
timestamp 1618419204
transform 1 0 4876 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1618419204
transform -1 0 8188 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.delayen1
timestamp 1618419204
transform 1 0 6808 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1618419204
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50
timestamp 1618419204
transform 1 0 5704 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_56
timestamp 1618419204
transform 1 0 6256 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_58
timestamp 1618419204
transform 1 0 6440 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_67
timestamp 1618419204
transform 1 0 7268 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen0
timestamp 1618419204
transform 1 0 8556 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1618419204
transform 1 0 9384 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1618419204
transform 1 0 10028 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_77
timestamp 1618419204
transform 1 0 8188 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_86
timestamp 1618419204
transform 1 0 9016 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_93
timestamp 1618419204
transform 1 0 9660 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1618419204
transform 1 0 12052 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1618419204
transform 1 0 10856 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1618419204
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_100
timestamp 1618419204
transform 1 0 10304 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_110
timestamp 1618419204
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1618419204
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1619507013
transform -1 0 13800 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfrbp_2  idiv8
timestamp 1618419204
transform 1 0 14260 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_6  FILLER_3_128
timestamp 1618419204
transform 1 0 12880 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_134
timestamp 1618419204
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_138
timestamp 1618419204
transform 1 0 13800 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_142
timestamp 1618419204
transform 1 0 14168 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1618419204
transform -1 0 17296 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1618419204
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_167
timestamp 1618419204
transform 1 0 16468 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_172
timestamp 1618419204
transform 1 0 16928 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen0
timestamp 1618419204
transform -1 0 3220 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb0
timestamp 1619507013
transform 1 0 1748 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1618419204
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1618419204
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_14
timestamp 1618419204
transform 1 0 2392 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_23
timestamp 1618419204
transform 1 0 3220 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb0
timestamp 1619507013
transform -1 0 5612 0 -1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1618419204
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_30
timestamp 1618419204
transform 1 0 3864 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_49
timestamp 1618419204
transform 1 0 5612 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1618419204
transform 1 0 7360 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.delayen0
timestamp 1619507013
transform 1 0 5980 0 -1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_4_64
timestamp 1618419204
transform 1 0 6992 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_71
timestamp 1618419204
transform 1 0 7636 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb0
timestamp 1619507013
transform -1 0 8648 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1618419204
transform -1 0 10304 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1618419204
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1618419204
transform 1 0 9384 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_82
timestamp 1618419204
transform 1 0 8648 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_87
timestamp 1618419204
transform 1 0 9108 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1618419204
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0
timestamp 1618419204
transform 1 0 10948 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen1
timestamp 1618419204
transform 1 0 11684 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_4_100
timestamp 1618419204
transform 1 0 10304 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_106
timestamp 1618419204
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_111
timestamp 1618419204
transform 1 0 11316 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_120
timestamp 1618419204
transform 1 0 12144 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _322_
timestamp 1618419204
transform -1 0 13616 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp 1618419204
transform -1 0 15548 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1618419204
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_136
timestamp 1618419204
transform 1 0 13616 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_142
timestamp 1618419204
transform 1 0 14168 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_144
timestamp 1618419204
transform 1 0 14352 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1618419204
transform 1 0 16192 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1618419204
transform -1 0 17296 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_157
timestamp 1618419204
transform 1 0 15548 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_163
timestamp 1618419204
transform 1 0 16100 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_167
timestamp 1618419204
transform 1 0 16468 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1618419204
transform 1 0 2760 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb1
timestamp 1619507013
transform 1 0 1748 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1618419204
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1618419204
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_14
timestamp 1618419204
transform 1 0 2392 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_21
timestamp 1618419204
transform 1 0 3036 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 4048 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.reseten0
timestamp 1619507013
transform 1 0 4416 0 1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_5_27
timestamp 1618419204
transform 1 0 3588 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_32
timestamp 1618419204
transform 1 0 4048 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1618419204
transform 1 0 5428 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _356_
timestamp 1618419204
transform -1 0 8648 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.iss.delayenb1
timestamp 1619507013
transform 1 0 6808 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1618419204
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_55
timestamp 1618419204
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_58
timestamp 1618419204
transform 1 0 6440 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_69
timestamp 1618419204
transform 1 0 7452 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _377_
timestamp 1618419204
transform -1 0 9844 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb1
timestamp 1619507013
transform -1 0 10856 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_5_82
timestamp 1618419204
transform 1 0 8648 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_95
timestamp 1618419204
transform 1 0 9844 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1618419204
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1618419204
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_106
timestamp 1618419204
transform 1 0 10856 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_115
timestamp 1618419204
transform 1 0 11684 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_122
timestamp 1618419204
transform 1 0 12328 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _324_
timestamp 1618419204
transform -1 0 14904 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb0
timestamp 1619507013
transform -1 0 13340 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_5_133
timestamp 1618419204
transform 1 0 13340 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_141
timestamp 1618419204
transform 1 0 14076 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb1
timestamp 1619507013
transform -1 0 15916 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1618419204
transform -1 0 17296 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1618419204
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_150
timestamp 1618419204
transform 1 0 14904 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_161
timestamp 1618419204
transform 1 0 15916 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1618419204
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_172
timestamp 1618419204
transform 1 0 16928 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1618419204
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1618419204
transform 1 0 1748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1618419204
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1618419204
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1618419204
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen1
timestamp 1618419204
transform 1 0 1840 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _360_
timestamp 1618419204
transform -1 0 2392 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_7_14
timestamp 1618419204
transform 1 0 2392 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_20
timestamp 1618419204
transform 1 0 2944 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_13
timestamp 1618419204
transform 1 0 2300 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1619507013
transform 1 0 2668 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb0
timestamp 1619507013
transform -1 0 3956 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_7_31
timestamp 1618419204
transform 1 0 3956 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_30
timestamp 1618419204
transform 1 0 3864 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_28
timestamp 1618419204
transform 1 0 3680 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1618419204
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_39
timestamp 1618419204
transform 1 0 4692 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_35
timestamp 1618419204
transform 1 0 4324 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1618419204
transform 1 0 4876 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1618419204
transform 1 0 4416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 4876 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_6_48
timestamp 1618419204
transform 1 0 5520 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1
timestamp 1619507013
transform 1 0 5244 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _314_
timestamp 1619507013
transform 1 0 5428 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _321_
timestamp 1619507013
transform 1 0 7268 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1618419204
transform 1 0 5888 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1618419204
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1618419204
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_61
timestamp 1618419204
transform 1 0 6716 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_73
timestamp 1618419204
transform 1 0 7820 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_53
timestamp 1618419204
transform 1 0 5980 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_58
timestamp 1618419204
transform 1 0 6440 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_71
timestamp 1618419204
transform 1 0 7636 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_81
timestamp 1618419204
transform 1 0 8556 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_80
timestamp 1618419204
transform 1 0 8464 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1618419204
transform 1 0 8188 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _306_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 8556 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1618419204
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1618419204
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _312_
timestamp 1619507013
transform -1 0 9476 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_91
timestamp 1618419204
transform 1 0 9476 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_94
timestamp 1618419204
transform 1 0 9752 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1618419204
transform -1 0 9752 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb1
timestamp 1619507013
transform 1 0 9844 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen1
timestamp 1618419204
transform -1 0 10580 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_7_106
timestamp 1618419204
transform 1 0 10856 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_102
timestamp 1618419204
transform 1 0 10488 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_103
timestamp 1618419204
transform 1 0 10580 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1618419204
transform -1 0 11224 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1618419204
transform 1 0 10948 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_115
timestamp 1618419204
transform 1 0 11684 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_110
timestamp 1618419204
transform 1 0 11224 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_110
timestamp 1618419204
transform 1 0 11224 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1618419204
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb1
timestamp 1619507013
transform 1 0 11592 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_7_124
timestamp 1618419204
transform 1 0 12512 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_121
timestamp 1618419204
transform 1 0 12236 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen1
timestamp 1618419204
transform -1 0 12512 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_7_132
timestamp 1618419204
transform 1 0 13248 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_132
timestamp 1618419204
transform 1 0 13248 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 1618419204
transform 1 0 12972 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_137
timestamp 1618419204
transform 1 0 13708 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_139
timestamp 1618419204
transform 1 0 13892 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1618419204
transform 1 0 13616 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1618419204
transform -1 0 13708 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_145
timestamp 1618419204
transform 1 0 14444 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_141
timestamp 1618419204
transform 1 0 14076 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1618419204
transform 1 0 14168 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1618419204
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen0
timestamp 1618419204
transform -1 0 14812 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1618419204
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb0
timestamp 1619507013
transform 1 0 14812 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_7_156
timestamp 1618419204
transform 1 0 15456 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_156
timestamp 1618419204
transform 1 0 15456 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1618419204
transform -1 0 15456 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_165
timestamp 1618419204
transform 1 0 16284 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_165
timestamp 1618419204
transform 1 0 16284 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen1
timestamp 1618419204
transform -1 0 16284 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen0
timestamp 1618419204
transform 1 0 15824 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_7_172
timestamp 1618419204
transform 1 0 16928 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1618419204
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1618419204
transform -1 0 17296 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1618419204
transform -1 0 17296 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1618419204
transform 1 0 1564 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[5\].id.delayen1
timestamp 1618419204
transform 1 0 2944 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1618419204
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1618419204
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_14
timestamp 1618419204
transform 1 0 2392 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 5520 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1619507013
transform -1 0 4876 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1618419204
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_25
timestamp 1618419204
transform 1 0 3404 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_30
timestamp 1618419204
transform 1 0 3864 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_41
timestamp 1618419204
transform 1 0 4876 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_47
timestamp 1618419204
transform 1 0 5428 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _369_
timestamp 1618419204
transform -1 0 8648 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1618419204
transform -1 0 6808 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1619507013
transform -1 0 7452 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_54
timestamp 1618419204
transform 1 0 6072 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_62
timestamp 1618419204
transform 1 0 6808 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_69
timestamp 1618419204
transform 1 0 7452 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1619507013
transform -1 0 10764 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1618419204
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1618419204
transform 1 0 9476 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_82
timestamp 1618419204
transform 1 0 8648 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_87
timestamp 1618419204
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_94
timestamp 1618419204
transform 1 0 9752 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 12512 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[4\].id.delayenb0
timestamp 1619507013
transform -1 0 12144 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_8_105
timestamp 1618419204
transform 1 0 10764 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_120
timestamp 1618419204
transform 1 0 12144 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1618419204
transform 1 0 14720 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen0
timestamp 1618419204
transform 1 0 13432 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1618419204
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_129
timestamp 1618419204
transform 1 0 12972 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_133
timestamp 1618419204
transform 1 0 13340 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_139
timestamp 1618419204
transform 1 0 13892 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_144
timestamp 1618419204
transform 1 0 14352 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1618419204
transform 1 0 16192 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1618419204
transform -1 0 17296 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1618419204
transform 1 0 15456 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_152
timestamp 1618419204
transform 1 0 15088 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_159
timestamp 1618419204
transform 1 0 15732 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_163
timestamp 1618419204
transform 1 0 16100 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_168
timestamp 1618419204
transform 1 0 16560 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_172
timestamp 1618419204
transform 1 0 16928 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1618419204
transform -1 0 2760 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1618419204
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1618419204
transform -1 0 1656 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_6
timestamp 1618419204
transform 1 0 1656 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_18
timestamp 1618419204
transform 1 0 2760 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _372_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 5980 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[5\].id.delayenb1
timestamp 1619507013
transform 1 0 3680 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_9_26
timestamp 1618419204
transform 1 0 3496 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_35
timestamp 1618419204
transform 1 0 4324 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_43
timestamp 1618419204
transform 1 0 5060 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 6808 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1618419204
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_53
timestamp 1618419204
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_58
timestamp 1618419204
transform 1 0 6440 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_69
timestamp 1618419204
transform 1 0 7452 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1619507013
transform 1 0 9016 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _319_
timestamp 1619507013
transform 1 0 8096 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _374_
timestamp 1618419204
transform -1 0 10488 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_75
timestamp 1618419204
transform 1 0 8004 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_82
timestamp 1618419204
transform 1 0 8648 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_89
timestamp 1618419204
transform 1 0 9292 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _368_
timestamp 1618419204
transform 1 0 12052 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1618419204
transform -1 0 11132 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1618419204
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_102
timestamp 1618419204
transform 1 0 10488 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_109
timestamp 1618419204
transform 1 0 11132 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1618419204
transform 1 0 11500 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_115
timestamp 1618419204
transform 1 0 11684 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1618419204
transform 1 0 13248 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_128
timestamp 1618419204
transform 1 0 12880 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_141
timestamp 1618419204
transform 1 0 14076 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_149
timestamp 1618419204
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1618419204
transform -1 0 15364 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1618419204
transform -1 0 17296 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1618419204
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1619507013
transform -1 0 16468 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_155
timestamp 1618419204
transform 1 0 15364 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_163
timestamp 1618419204
transform 1 0 16100 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_167
timestamp 1618419204
transform 1 0 16468 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_172
timestamp 1618419204
transform 1 0 16928 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1618419204
transform 1 0 3128 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb0
timestamp 1619507013
transform 1 0 1380 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1618419204
transform -1 0 2760 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1618419204
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_10
timestamp 1618419204
transform 1 0 2024 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_14
timestamp 1618419204
transform 1 0 2392 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_18
timestamp 1618419204
transform 1 0 2760 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1619507013
transform -1 0 5244 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _354_
timestamp 1618419204
transform -1 0 6440 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1618419204
transform 1 0 4232 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1618419204
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_25
timestamp 1618419204
transform 1 0 3404 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_30
timestamp 1618419204
transform 1 0 3864 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_37
timestamp 1618419204
transform 1 0 4508 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_41
timestamp 1618419204
transform 1 0 4876 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_45
timestamp 1618419204
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _300_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 7176 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _302_
timestamp 1618419204
transform 1 0 7544 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_58
timestamp 1618419204
transform 1 0 6440 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_66
timestamp 1618419204
transform 1 0 7176 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_74
timestamp 1618419204
transform 1 0 7912 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1619507013
transform -1 0 8556 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _315_
timestamp 1619507013
transform -1 0 9936 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1618419204
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_81
timestamp 1618419204
transform 1 0 8556 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1618419204
transform 1 0 8924 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1618419204
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_96
timestamp 1618419204
transform 1 0 9936 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1619507013
transform 1 0 10304 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 11040 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _347_
timestamp 1618419204
transform -1 0 12788 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1618419204
transform 1 0 11868 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_103
timestamp 1618419204
transform 1 0 10580 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_107
timestamp 1618419204
transform 1 0 10948 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_113
timestamp 1618419204
transform 1 0 11500 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_120
timestamp 1618419204
transform 1 0 12144 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb0
timestamp 1619507013
transform 1 0 13156 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1618419204
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1619507013
transform -1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_127
timestamp 1618419204
transform 1 0 12788 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_138
timestamp 1618419204
transform 1 0 13800 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_142
timestamp 1618419204
transform 1 0 14168 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_144
timestamp 1618419204
transform 1 0 14352 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb0
timestamp 1619507013
transform 1 0 15272 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1618419204
transform -1 0 17296 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1618419204
transform 1 0 16376 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_150
timestamp 1618419204
transform 1 0 14904 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_161
timestamp 1618419204
transform 1 0 15916 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_165
timestamp 1618419204
transform 1 0 16284 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_169
timestamp 1618419204
transform 1 0 16652 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb1
timestamp 1619507013
transform -1 0 3220 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1618419204
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output39
timestamp 1618419204
transform -1 0 1748 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_7
timestamp 1618419204
transform 1 0 1748 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp 1618419204
transform 1 0 2484 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_23
timestamp 1618419204
transform 1 0 3220 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _304_
timestamp 1618419204
transform 1 0 5336 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1618419204
transform 1 0 4140 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_31
timestamp 1618419204
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_42
timestamp 1618419204
transform 1 0 4968 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _298_
timestamp 1618419204
transform -1 0 8004 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1618419204
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_53
timestamp 1618419204
transform 1 0 5980 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_58
timestamp 1618419204
transform 1 0 6440 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_66
timestamp 1618419204
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__a31o_1  _308_
timestamp 1618419204
transform 1 0 10028 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__buf_8  repeater46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 8556 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_75
timestamp 1618419204
transform 1 0 8004 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_93
timestamp 1618419204
transform 1 0 9660 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1618419204
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1618419204
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1618419204
transform 1 0 11776 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_104
timestamp 1618419204
transform 1 0 10672 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_112
timestamp 1618419204
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_115
timestamp 1618419204
transform 1 0 11684 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_119
timestamp 1618419204
transform 1 0 12052 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1618419204
transform -1 0 14168 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1618419204
transform 1 0 14628 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_132
timestamp 1618419204
transform 1 0 13248 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_138
timestamp 1618419204
transform 1 0 13800 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_142
timestamp 1618419204
transform 1 0 14168 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_146
timestamp 1618419204
transform 1 0 14536 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen0
timestamp 1618419204
transform 1 0 15272 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1618419204
transform 1 0 16100 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1618419204
transform -1 0 17296 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1618419204
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_150
timestamp 1618419204
transform 1 0 14904 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1618419204
transform 1 0 15732 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_166
timestamp 1618419204
transform 1 0 16376 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_170
timestamp 1618419204
transform 1 0 16744 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_172
timestamp 1618419204
transform 1 0 16928 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen0
timestamp 1618419204
transform 1 0 1840 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen1
timestamp 1618419204
transform -1 0 3220 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1618419204
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1618419204
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1618419204
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_13
timestamp 1618419204
transform 1 0 2300 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_17
timestamp 1618419204
transform 1 0 2668 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_23
timestamp 1618419204
transform 1 0 3220 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _366_
timestamp 1618419204
transform 1 0 4508 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1618419204
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_30
timestamp 1618419204
transform 1 0 3864 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_36
timestamp 1618419204
transform 1 0 4416 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_46
timestamp 1618419204
transform 1 0 5336 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _293_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 6164 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _296_
timestamp 1618419204
transform -1 0 6992 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _301_
timestamp 1618419204
transform 1 0 7360 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_55
timestamp 1618419204
transform 1 0 6164 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_64
timestamp 1618419204
transform 1 0 6992 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_72
timestamp 1618419204
transform 1 0 7728 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 10304 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _317_
timestamp 1619507013
transform -1 0 8648 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1618419204
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_82
timestamp 1618419204
transform 1 0 8648 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1618419204
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _365_
timestamp 1618419204
transform 1 0 10764 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _371_
timestamp 1618419204
transform -1 0 12788 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_100
timestamp 1618419204
transform 1 0 10304 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_104
timestamp 1618419204
transform 1 0 10672 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_114
timestamp 1618419204
transform 1 0 11592 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1618419204
transform 1 0 14720 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb1
timestamp 1619507013
transform 1 0 13248 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1618419204
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_127
timestamp 1618419204
transform 1 0 12788 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_131
timestamp 1618419204
transform 1 0 13156 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_139
timestamp 1618419204
transform 1 0 13892 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_144
timestamp 1618419204
transform 1 0 14352 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb1
timestamp 1619507013
transform 1 0 15456 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1618419204
transform -1 0 17296 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_151
timestamp 1618419204
transform 1 0 14996 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_155
timestamp 1618419204
transform 1 0 15364 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_163
timestamp 1618419204
transform 1 0 16100 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_171
timestamp 1618419204
transform 1 0 16836 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_7
timestamp 1618419204
transform 1 0 1748 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output40
timestamp 1618419204
transform -1 0 1748 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1618419204
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1618419204
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _364_
timestamp 1618419204
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_15
timestamp 1618419204
transform 1 0 2484 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_12
timestamp 1618419204
transform 1 0 2208 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb1
timestamp 1619507013
transform -1 0 3220 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1618419204
transform -1 0 2944 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_23
timestamp 1618419204
transform 1 0 3220 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_20
timestamp 1618419204
transform 1 0 2944 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_36
timestamp 1618419204
transform 1 0 4416 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_30
timestamp 1618419204
transform 1 0 3864 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_30
timestamp 1618419204
transform 1 0 3864 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_26
timestamp 1618419204
transform 1 0 3496 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1618419204
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _294_
timestamp 1618419204
transform 1 0 4508 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1619507013
transform 1 0 3588 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_46
timestamp 1618419204
transform 1 0 5336 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_42
timestamp 1618419204
transform 1 0 4968 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1619507013
transform -1 0 5704 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_8  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 5704 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_14_50
timestamp 1618419204
transform 1 0 5704 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_58
timestamp 1618419204
transform 1 0 6440 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_56
timestamp 1618419204
transform 1 0 6256 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1618419204
transform 1 0 5704 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1618419204
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _305_
timestamp 1618419204
transform 1 0 6072 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_14_65
timestamp 1618419204
transform 1 0 7084 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_61
timestamp 1618419204
transform 1 0 6716 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_67
timestamp 1618419204
transform 1 0 7268 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _310_
timestamp 1619507013
transform -1 0 7636 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _248_
timestamp 1618419204
transform 1 0 6808 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_14_71
timestamp 1618419204
transform 1 0 7636 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_80
timestamp 1618419204
transform 1 0 8464 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_75
timestamp 1618419204
transform 1 0 8004 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _311_
timestamp 1619507013
transform 1 0 8096 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _309_
timestamp 1618419204
transform 1 0 8004 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_14_87
timestamp 1618419204
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_89
timestamp 1618419204
transform 1 0 9292 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_85
timestamp 1618419204
transform 1 0 8924 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1618419204
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__o41a_1  _320_
timestamp 1618419204
transform 1 0 9476 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _254_
timestamp 1618419204
transform 1 0 9384 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_13_97
timestamp 1618419204
transform 1 0 10028 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 1618419204
transform 1 0 11132 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_100
timestamp 1618419204
transform 1 0 10304 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1618419204
transform -1 0 11224 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _290_
timestamp 1618419204
transform 1 0 10672 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_14_116
timestamp 1618419204
transform 1 0 11776 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_115
timestamp 1618419204
transform 1 0 11684 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_110
timestamp 1618419204
transform 1 0 11224 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1619507013
transform -1 0 12236 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1618419204
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 11776 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_120
timestamp 1618419204
transform 1 0 12144 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_121
timestamp 1618419204
transform 1 0 12236 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _292_
timestamp 1618419204
transform 1 0 12236 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_14_133
timestamp 1618419204
transform 1 0 13340 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_126
timestamp 1618419204
transform 1 0 12696 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_134
timestamp 1618419204
transform 1 0 13432 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1618419204
transform 1 0 13064 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1618419204
transform -1 0 13432 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1618419204
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_143
timestamp 1618419204
transform 1 0 14260 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1618419204
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen1
timestamp 1618419204
transform 1 0 13800 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_14_144
timestamp 1618419204
transform 1 0 14352 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_149
timestamp 1618419204
transform 1 0 14812 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1618419204
transform -1 0 14996 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_151
timestamp 1618419204
transform 1 0 14996 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen1
timestamp 1618419204
transform 1 0 15548 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _373_
timestamp 1618419204
transform -1 0 15732 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_162
timestamp 1618419204
transform 1 0 16008 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_167
timestamp 1618419204
transform 1 0 16468 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_163
timestamp 1618419204
transform 1 0 16100 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_159
timestamp 1618419204
transform 1 0 15732 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1618419204
transform 1 0 16192 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1618419204
transform 1 0 16376 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_169
timestamp 1618419204
transform 1 0 16652 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_172
timestamp 1618419204
transform 1 0 16928 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1618419204
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1618419204
transform -1 0 17296 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1618419204
transform -1 0 17296 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1618419204
transform -1 0 2208 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen1
timestamp 1618419204
transform -1 0 3220 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1618419204
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_12
timestamp 1618419204
transform 1 0 2208 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_23
timestamp 1618419204
transform 1 0 3220 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1619507013
transform -1 0 5336 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _273_
timestamp 1618419204
transform 1 0 4232 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1618419204
transform -1 0 3864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_30
timestamp 1618419204
transform 1 0 3864 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_38
timestamp 1618419204
transform 1 0 4600 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_42
timestamp 1618419204
transform 1 0 4968 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_46
timestamp 1618419204
transform 1 0 5336 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1619507013
transform 1 0 7084 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1619507013
transform 1 0 5704 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1618419204
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_53
timestamp 1618419204
transform 1 0 5980 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_58
timestamp 1618419204
transform 1 0 6440 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_64
timestamp 1618419204
transform 1 0 6992 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_68
timestamp 1618419204
transform 1 0 7360 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1619507013
transform 1 0 9936 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1618419204
transform 1 0 8188 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_76
timestamp 1618419204
transform 1 0 8096 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_86
timestamp 1618419204
transform 1 0 9016 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_94
timestamp 1618419204
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_99
timestamp 1618419204
transform 1 0 10212 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _199_
timestamp 1619507013
transform -1 0 11224 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1618419204
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1618419204
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_110
timestamp 1618419204
transform 1 0 11224 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_115
timestamp 1618419204
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_122
timestamp 1618419204
transform 1 0 12328 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _341_
timestamp 1618419204
transform 1 0 12880 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _385_
timestamp 1619507013
transform 1 0 13800 0 1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_6  FILLER_15_131
timestamp 1618419204
transform 1 0 13156 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_137
timestamp 1618419204
transform 1 0 13708 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1618419204
transform -1 0 17296 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1618419204
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_161
timestamp 1618419204
transform 1 0 15916 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1618419204
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_172
timestamp 1618419204
transform 1 0 16928 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen0
timestamp 1618419204
transform -1 0 2944 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb0
timestamp 1619507013
transform 1 0 1472 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1618419204
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1618419204
transform 1 0 1380 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_11
timestamp 1618419204
transform 1 0 2116 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1618419204
transform 1 0 2944 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _392_
timestamp 1619507013
transform 1 0 4232 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1618419204
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_28
timestamp 1618419204
transform 1 0 3680 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_30
timestamp 1618419204
transform 1 0 3864 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _258_
timestamp 1619507013
transform 1 0 6992 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_16_55
timestamp 1618419204
transform 1 0 6164 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_63
timestamp 1618419204
transform 1 0 6900 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_71
timestamp 1618419204
transform 1 0 7636 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _261_
timestamp 1618419204
transform -1 0 8372 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _401_
timestamp 1619507013
transform 1 0 9568 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1618419204
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_79
timestamp 1618419204
transform 1 0 8372 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1618419204
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1618419204
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1618419204
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _386_
timestamp 1619507013
transform 1 0 11776 0 -1 11424
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_16_112
timestamp 1618419204
transform 1 0 11408 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _400_
timestamp 1619507013
transform 1 0 14812 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1618419204
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_139
timestamp 1618419204
transform 1 0 13892 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_144
timestamp 1618419204
transform 1 0 14352 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_148
timestamp 1618419204
transform 1 0 14720 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1618419204
transform -1 0 17296 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_169
timestamp 1618419204
transform 1 0 16652 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1618419204
transform -1 0 2208 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1618419204
transform -1 0 2944 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1618419204
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1618419204
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_12
timestamp 1618419204
transform 1 0 2208 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_20
timestamp 1618419204
transform 1 0 2944 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _246_
timestamp 1619507013
transform 1 0 5336 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1619507013
transform -1 0 3864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 4232 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_26
timestamp 1618419204
transform 1 0 3496 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_30
timestamp 1618419204
transform 1 0 3864 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_42
timestamp 1618419204
transform 1 0 4968 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _260_
timestamp 1618419204
transform 1 0 6808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1618419204
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_53
timestamp 1618419204
transform 1 0 5980 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_58
timestamp 1618419204
transform 1 0 6440 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_70
timestamp 1618419204
transform 1 0 7544 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _395_
timestamp 1619507013
transform 1 0 8464 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_17_78
timestamp 1618419204
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1618419204
transform 1 0 10764 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _343_
timestamp 1618419204
transform -1 0 12328 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1618419204
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_101
timestamp 1618419204
transform 1 0 10396 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_108
timestamp 1618419204
transform 1 0 11040 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_115
timestamp 1618419204
transform 1 0 11684 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_122
timestamp 1618419204
transform 1 0 12328 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1619507013
transform -1 0 14996 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _279_
timestamp 1618419204
transform -1 0 13156 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 14352 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_131
timestamp 1618419204
transform 1 0 13156 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1618419204
transform 1 0 14352 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 15364 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1618419204
transform -1 0 17296 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1618419204
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_151
timestamp 1618419204
transform 1 0 14996 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_163
timestamp 1618419204
transform 1 0 16100 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_172
timestamp 1618419204
transform 1 0 16928 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _267_
timestamp 1618419204
transform 1 0 3128 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1618419204
transform -1 0 2760 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1618419204
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1618419204
transform -1 0 2116 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1618419204
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1618419204
transform 1 0 1748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_11
timestamp 1618419204
transform 1 0 2116 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_18
timestamp 1618419204
transform 1 0 2760 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1619507013
transform -1 0 5244 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _270_
timestamp 1618419204
transform -1 0 4600 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1618419204
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_25
timestamp 1618419204
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_30
timestamp 1618419204
transform 1 0 3864 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_38
timestamp 1618419204
transform 1 0 4600 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_45
timestamp 1618419204
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_49
timestamp 1618419204
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _252_
timestamp 1619507013
transform 1 0 7452 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _256_
timestamp 1619507013
transform 1 0 6348 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1619507013
transform -1 0 5980 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_53
timestamp 1618419204
transform 1 0 5980 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_65
timestamp 1618419204
transform 1 0 7084 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1619507013
transform 1 0 9476 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1618419204
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_76
timestamp 1618419204
transform 1 0 8096 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1618419204
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1618419204
transform 1 0 9108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_94
timestamp 1618419204
transform 1 0 9752 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _223_
timestamp 1619507013
transform 1 0 11776 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 10672 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1618419204
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1618419204
transform 1 0 11408 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_120
timestamp 1618419204
transform 1 0 12144 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_124
timestamp 1618419204
transform 1 0 12512 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1619507013
transform 1 0 13616 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _286_
timestamp 1618419204
transform 1 0 12604 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1618419204
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_132
timestamp 1618419204
transform 1 0 13248 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_139
timestamp 1618419204
transform 1 0 13892 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_144
timestamp 1618419204
transform 1 0 14352 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _200_
timestamp 1619507013
transform -1 0 15732 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1618419204
transform -1 0 17296 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1619507013
transform -1 0 16652 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_159
timestamp 1618419204
transform 1 0 15732 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_165
timestamp 1618419204
transform 1 0 16284 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_169
timestamp 1618419204
transform 1 0 16652 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 2668 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1618419204
transform -1 0 2300 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _391_
timestamp 1619507013
transform 1 0 1380 0 1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1618419204
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1618419204
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1618419204
transform -1 0 1656 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_24
timestamp 1618419204
transform 1 0 3312 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_6
timestamp 1618419204
transform 1 0 1656 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_13
timestamp 1618419204
transform 1 0 2300 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_30
timestamp 1618419204
transform 1 0 3864 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_25
timestamp 1618419204
transform 1 0 3404 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_31
timestamp 1618419204
transform 1 0 3956 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1618419204
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1619507013
transform 1 0 3680 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_39
timestamp 1618419204
transform 1 0 4692 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_35
timestamp 1618419204
transform 1 0 4324 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _269_
timestamp 1618419204
transform -1 0 4692 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _250_
timestamp 1619507013
transform 1 0 4416 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_46
timestamp 1618419204
transform 1 0 5336 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_44
timestamp 1618419204
transform 1 0 5152 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1619507013
transform 1 0 5060 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_58
timestamp 1618419204
transform 1 0 6440 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_50
timestamp 1618419204
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_58
timestamp 1618419204
transform 1 0 6440 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_53
timestamp 1618419204
transform 1 0 5980 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1618419204
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1619507013
transform -1 0 5980 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _251_
timestamp 1619507013
transform -1 0 6440 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_20_67
timestamp 1618419204
transform 1 0 7268 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _265_
timestamp 1618419204
transform 1 0 7176 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _262_
timestamp 1618419204
transform 1 0 6808 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_20_73
timestamp 1618419204
transform 1 0 7820 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_74
timestamp 1618419204
transform 1 0 7912 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _266_
timestamp 1618419204
transform -1 0 8280 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1619507013
transform 1 0 9476 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _394_
timestamp 1619507013
transform 1 0 8280 0 1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1618419204
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_99
timestamp 1618419204
transform 1 0 10212 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_78
timestamp 1618419204
transform 1 0 8280 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_87
timestamp 1618419204
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_94
timestamp 1618419204
transform 1 0 9752 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1618419204
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__o2bb2a_1  _212_
timestamp 1618419204
transform 1 0 10672 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1619507013
transform 1 0 10948 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_112
timestamp 1618419204
transform 1 0 11408 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_115
timestamp 1618419204
transform 1 0 11684 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_110
timestamp 1618419204
transform 1 0 11224 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1618419204
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp 1618419204
transform 1 0 11776 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_119
timestamp 1618419204
transform 1 0 12052 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_122
timestamp 1618419204
transform 1 0 12328 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _207_
timestamp 1619507013
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_132
timestamp 1618419204
transform 1 0 13248 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_130
timestamp 1618419204
transform 1 0 13064 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _285_
timestamp 1618419204
transform -1 0 13064 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 12604 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_20_139
timestamp 1618419204
transform 1 0 13892 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_136
timestamp 1618419204
transform 1 0 13616 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _288_
timestamp 1618419204
transform 1 0 13708 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1619507013
transform 1 0 13616 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_144
timestamp 1618419204
transform 1 0 14352 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_142
timestamp 1618419204
transform 1 0 14168 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1618419204
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1619507013
transform 1 0 14536 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_149
timestamp 1618419204
transform 1 0 14812 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2ai_1  _228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 15364 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_20_155
timestamp 1618419204
transform 1 0 15364 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _210_
timestamp 1619507013
transform -1 0 15824 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_20_164
timestamp 1618419204
transform 1 0 16192 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_160
timestamp 1618419204
transform 1 0 15824 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1618419204
transform 1 0 16192 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _208_
timestamp 1619507013
transform -1 0 16192 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_20_172
timestamp 1618419204
transform 1 0 16928 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_172
timestamp 1618419204
transform 1 0 16928 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_167
timestamp 1618419204
transform 1 0 16468 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1618419204
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1618419204
transform -1 0 17296 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1618419204
transform -1 0 17296 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _244_
timestamp 1619507013
transform 1 0 3312 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _274_
timestamp 1618419204
transform -1 0 2944 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1618419204
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1619507013
transform 1 0 1840 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1618419204
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1618419204
transform 1 0 1748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_11
timestamp 1618419204
transform 1 0 2116 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_20
timestamp 1618419204
transform 1 0 2944 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1619507013
transform 1 0 4324 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _268_
timestamp 1618419204
transform 1 0 5244 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_31
timestamp 1618419204
transform 1 0 3956 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_38
timestamp 1618419204
transform 1 0 4600 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_44
timestamp 1618419204
transform 1 0 5152 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _263_
timestamp 1618419204
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1618419204
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_53
timestamp 1618419204
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_58
timestamp 1618419204
transform 1 0 6440 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_66
timestamp 1618419204
transform 1 0 7176 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_74
timestamp 1618419204
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__o2bb2a_1  _220_
timestamp 1618419204
transform 1 0 9384 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 8832 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_84
timestamp 1618419204
transform 1 0 8832 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_98
timestamp 1618419204
transform 1 0 10120 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _198_
timestamp 1619507013
transform 1 0 10580 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _384_
timestamp 1619507013
transform 1 0 12328 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1618419204
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_102
timestamp 1618419204
transform 1 0 10488 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_110
timestamp 1618419204
transform 1 0 11224 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_115
timestamp 1618419204
transform 1 0 11684 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1618419204
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _399_
timestamp 1619507013
transform 1 0 14628 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_21_142
timestamp 1618419204
transform 1 0 14168 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_146
timestamp 1618419204
transform 1 0 14536 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1618419204
transform -1 0 17296 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1618419204
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_167
timestamp 1618419204
transform 1 0 16468 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_172
timestamp 1618419204
transform 1 0 16928 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _241_
timestamp 1618419204
transform 1 0 2300 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _276_
timestamp 1618419204
transform -1 0 3404 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1618419204
transform -1 0 1932 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1618419204
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1618419204
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_9
timestamp 1618419204
transform 1 0 1932 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_16
timestamp 1618419204
transform 1 0 2576 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _393_
timestamp 1619507013
transform 1 0 4508 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1618419204
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_25
timestamp 1618419204
transform 1 0 3404 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_30
timestamp 1618419204
transform 1 0 3864 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_36
timestamp 1618419204
transform 1 0 4416 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__or3_1  _237_
timestamp 1618419204
transform 1 0 7360 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_22_58
timestamp 1618419204
transform 1 0 6440 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_66
timestamp 1618419204
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_73
timestamp 1618419204
transform 1 0 7820 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _219_
timestamp 1618419204
transform 1 0 9752 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _221_
timestamp 1618419204
transform 1 0 8188 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1618419204
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_82
timestamp 1618419204
transform 1 0 8648 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_87
timestamp 1618419204
transform 1 0 9108 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_93
timestamp 1618419204
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _402_
timestamp 1619507013
transform 1 0 10672 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_22_100
timestamp 1618419204
transform 1 0 10304 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1618419204
transform 1 0 12512 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _289_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 12880 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1618419204
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_136
timestamp 1618419204
transform 1 0 13616 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_142
timestamp 1618419204
transform 1 0 14168 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_144
timestamp 1618419204
transform 1 0 14352 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _201_
timestamp 1619507013
transform -1 0 15548 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _227_
timestamp 1618419204
transform -1 0 16468 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1618419204
transform -1 0 17296 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_157
timestamp 1618419204
transform 1 0 15548 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_167
timestamp 1618419204
transform 1 0 16468 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _390_
timestamp 1619507013
transform 1 0 1380 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1618419204
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_23
timestamp 1618419204
transform 1 0 3220 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _240_
timestamp 1619507013
transform 1 0 3588 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _242_
timestamp 1618419204
transform -1 0 4968 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_34
timestamp 1618419204
transform 1 0 4232 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_42
timestamp 1618419204
transform 1 0 4968 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1619507013
transform 1 0 5704 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 6808 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_4  _238_
timestamp 1619507013
transform 1 0 7912 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1618419204
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_53
timestamp 1618419204
transform 1 0 5980 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_58
timestamp 1618419204
transform 1 0 6440 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_69
timestamp 1618419204
transform 1 0 7452 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_73
timestamp 1618419204
transform 1 0 7820 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _213_
timestamp 1618419204
transform 1 0 10120 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_91
timestamp 1618419204
transform 1 0 9476 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_97
timestamp 1618419204
transform 1 0 10028 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _206_
timestamp 1619507013
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1618419204
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_106
timestamp 1618419204
transform 1 0 10856 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_115
timestamp 1618419204
transform 1 0 11684 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_122
timestamp 1618419204
transform 1 0 12328 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _229_
timestamp 1618419204
transform -1 0 13248 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _231_
timestamp 1618419204
transform -1 0 15364 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 13616 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_128
timestamp 1618419204
transform 1 0 12880 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_132
timestamp 1618419204
transform 1 0 13248 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_142
timestamp 1618419204
transform 1 0 14168 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1619507013
transform 1 0 15732 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1618419204
transform -1 0 17296 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1618419204
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_155
timestamp 1618419204
transform 1 0 15364 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_162
timestamp 1618419204
transform 1 0 16008 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_170
timestamp 1618419204
transform 1 0 16744 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_172
timestamp 1618419204
transform 1 0 16928 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_1  _277_
timestamp 1618419204
transform 1 0 2484 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1618419204
transform -1 0 2116 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1618419204
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1618419204
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1618419204
transform 1 0 1748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_11
timestamp 1618419204
transform 1 0 2116 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_23
timestamp 1618419204
transform 1 0 3220 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1619507013
transform 1 0 4232 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1619507013
transform -1 0 5428 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1618419204
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_30
timestamp 1618419204
transform 1 0 3864 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_37
timestamp 1618419204
transform 1 0 4508 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_43
timestamp 1618419204
transform 1 0 5060 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_47
timestamp 1618419204
transform 1 0 5428 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _202_
timestamp 1619507013
transform -1 0 6440 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 8096 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_58
timestamp 1618419204
transform 1 0 6440 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _214_
timestamp 1618419204
transform 1 0 10028 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1618419204
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_76
timestamp 1618419204
transform 1 0 8096 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1618419204
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_87
timestamp 1618419204
transform 1 0 9108 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_95
timestamp 1618419204
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _236_
timestamp 1618419204
transform -1 0 11224 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _283_
timestamp 1618419204
transform 1 0 11960 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1618419204
transform 1 0 10488 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_110
timestamp 1618419204
transform 1 0 11224 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1619507013
transform -1 0 13892 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _383_
timestamp 1619507013
transform 1 0 14812 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1618419204
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_127
timestamp 1618419204
transform 1 0 12788 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_135
timestamp 1618419204
transform 1 0 13524 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_139
timestamp 1618419204
transform 1 0 13892 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_144
timestamp 1618419204
transform 1 0 14352 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_148
timestamp 1618419204
transform 1 0 14720 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1618419204
transform -1 0 17296 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_169
timestamp 1618419204
transform 1 0 16652 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1619507013
transform -1 0 3036 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1618419204
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1618419204
transform -1 0 2392 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1619507013
transform 1 0 1472 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1618419204
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_7
timestamp 1618419204
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_14
timestamp 1618419204
transform 1 0 2392 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_21
timestamp 1618419204
transform 1 0 3036 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _398_
timestamp 1619507013
transform 1 0 3864 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_25_29
timestamp 1618419204
transform 1 0 3772 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_2  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 6808 0 1 15776
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1618419204
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_50
timestamp 1618419204
transform 1 0 5704 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_56
timestamp 1618419204
transform 1 0 6256 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_58
timestamp 1618419204
transform 1 0 6440 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_72
timestamp 1618419204
transform 1 0 7728 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _216_
timestamp 1618419204
transform 1 0 9752 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_2  _234_
timestamp 1619507013
transform 1 0 8096 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_85
timestamp 1618419204
transform 1 0 8924 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_93
timestamp 1618419204
transform 1 0 9660 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1619507013
transform 1 0 10948 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _387_
timestamp 1619507013
transform 1 0 12420 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1618419204
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1619507013
transform -1 0 12052 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_103
timestamp 1618419204
transform 1 0 10580 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_110
timestamp 1618419204
transform 1 0 11224 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_115
timestamp 1618419204
transform 1 0 11684 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_119
timestamp 1618419204
transform 1 0 12052 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_144
timestamp 1618419204
transform 1 0 14352 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_4  _193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 16468 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1618419204
transform -1 0 17296 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1618419204
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_150
timestamp 1618419204
transform 1 0 14904 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_167
timestamp 1618419204
transform 1 0 16468 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_172
timestamp 1618419204
transform 1 0 16928 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _278_
timestamp 1619507013
transform 1 0 2392 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _338_
timestamp 1618419204
transform -1 0 2024 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _389_
timestamp 1619507013
transform 1 0 1380 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1618419204
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1618419204
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_23
timestamp 1618419204
transform 1 0 3220 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1618419204
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_10
timestamp 1618419204
transform 1 0 2024 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_21
timestamp 1618419204
transform 1 0 3036 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _203_
timestamp 1619507013
transform 1 0 5244 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1619507013
transform 1 0 4600 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 1618419204
transform 1 0 5612 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _396_
timestamp 1619507013
transform 1 0 3404 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1618419204
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_30
timestamp 1618419204
transform 1 0 3864 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_41
timestamp 1618419204
transform 1 0 4876 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_45
timestamp 1618419204
transform 1 0 5244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_58
timestamp 1618419204
transform 1 0 6440 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_56
timestamp 1618419204
transform 1 0 6256 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1618419204
transform 1 0 5888 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_52
timestamp 1618419204
transform 1 0 5888 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1618419204
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_74
timestamp 1618419204
transform 1 0 7912 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_70
timestamp 1618419204
transform 1 0 7544 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_66
timestamp 1618419204
transform 1 0 7176 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1618419204
transform -1 0 7544 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _397_
timestamp 1619507013
transform 1 0 6256 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__a22o_1  _195_
timestamp 1619507013
transform -1 0 10856 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _215_
timestamp 1618419204
transform -1 0 10488 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _403_
timestamp 1619507013
transform -1 0 9844 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1618419204
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_76
timestamp 1618419204
transform 1 0 8096 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_84
timestamp 1618419204
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_87
timestamp 1618419204
transform 1 0 9108 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_93
timestamp 1618419204
transform 1 0 9660 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_95
timestamp 1618419204
transform 1 0 9844 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1619507013
transform 1 0 12052 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _205_
timestamp 1619507013
transform -1 0 11500 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_2  _388_
timestamp 1619507013
transform -1 0 13984 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1618419204
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_102
timestamp 1618419204
transform 1 0 10488 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_113
timestamp 1618419204
transform 1 0 11500 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_122
timestamp 1618419204
transform 1 0 12328 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_106
timestamp 1618419204
transform 1 0 10856 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_115
timestamp 1618419204
transform 1 0 11684 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_136
timestamp 1618419204
transform 1 0 13616 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_129
timestamp 1618419204
transform 1 0 12972 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp 1618419204
transform -1 0 13616 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1618419204
transform -1 0 12972 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_140
timestamp 1618419204
transform 1 0 13984 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_144
timestamp 1618419204
transform 1 0 14352 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_142
timestamp 1618419204
transform 1 0 14168 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1618419204
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _382_
timestamp 1619507013
transform 1 0 14720 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _381_
timestamp 1619507013
transform 1 0 14352 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1618419204
transform -1 0 17296 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1618419204
transform -1 0 17296 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1618419204
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_168
timestamp 1618419204
transform 1 0 16560 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_172
timestamp 1618419204
transform 1 0 16928 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_164
timestamp 1618419204
transform 1 0 16192 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_170
timestamp 1618419204
transform 1 0 16744 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_172
timestamp 1618419204
transform 1 0 16928 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _349_
timestamp 1618419204
transform 1 0 2116 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1618419204
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1619507013
transform 1 0 3128 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output44
timestamp 1618419204
transform -1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_7
timestamp 1618419204
transform 1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_14
timestamp 1618419204
transform 1 0 2392 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _204_
timestamp 1618419204
transform -1 0 5704 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1618419204
transform -1 0 4876 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1618419204
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_25
timestamp 1618419204
transform 1 0 3404 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_30
timestamp 1618419204
transform 1 0 3864 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_41
timestamp 1618419204
transform 1 0 4876 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp 1618419204
transform -1 0 7912 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1618419204
transform 1 0 6440 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1618419204
transform -1 0 7268 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_50
timestamp 1618419204
transform 1 0 5704 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_59
timestamp 1618419204
transform 1 0 6532 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_63
timestamp 1618419204
transform 1 0 6900 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_67
timestamp 1618419204
transform 1 0 7268 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_74
timestamp 1618419204
transform 1 0 7912 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1619507013
transform -1 0 8556 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _218_
timestamp 1618419204
transform -1 0 9844 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1618419204
transform 1 0 9108 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_81
timestamp 1618419204
transform 1 0 8556 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_88
timestamp 1618419204
transform 1 0 9200 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_95
timestamp 1618419204
transform 1 0 9844 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _345_
timestamp 1618419204
transform -1 0 11408 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp 1618419204
transform -1 0 10764 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1618419204
transform 1 0 11776 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1618419204
transform -1 0 12604 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_101
timestamp 1618419204
transform 1 0 10396 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_105
timestamp 1618419204
transform 1 0 10764 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_112
timestamp 1618419204
transform 1 0 11408 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_117
timestamp 1618419204
transform 1 0 11868 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_121
timestamp 1618419204
transform 1 0 12236 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_1  _282_
timestamp 1619507013
transform -1 0 15088 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _339_
timestamp 1618419204
transform -1 0 13248 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp 1618419204
transform -1 0 14076 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1618419204
transform 1 0 14444 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_125
timestamp 1618419204
transform 1 0 12604 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_132
timestamp 1618419204
transform 1 0 13248 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1618419204
transform 1 0 14076 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_146
timestamp 1618419204
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1618419204
transform -1 0 17296 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1618419204
transform -1 0 16652 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output42
timestamp 1618419204
transform 1 0 15548 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1618419204
transform 1 0 15088 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_156
timestamp 1618419204
transform 1 0 15456 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_161
timestamp 1618419204
transform 1 0 15916 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_169
timestamp 1618419204
transform 1 0 16652 0 -1 17952
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 8168 800 8288 6 clockc
port 0 nsew signal tristate
rlabel metal3 s 0 10208 800 10328 6 clockd[0]
port 1 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 clockd[1]
port 2 nsew signal tristate
rlabel metal3 s 17660 17008 18460 17128 6 clockd[2]
port 3 nsew signal tristate
rlabel metal2 s 16578 0 16634 800 6 clockd[3]
port 4 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 clockp[0]
port 5 nsew signal tristate
rlabel metal2 s 1398 0 1454 800 6 clockp[1]
port 6 nsew signal tristate
rlabel metal2 s 12438 0 12494 800 6 dco
port 7 nsew signal input
rlabel metal3 s 17660 12928 18460 13048 6 div[0]
port 8 nsew signal input
rlabel metal2 s 15658 19804 15714 20604 6 div[1]
port 9 nsew signal input
rlabel metal2 s 5998 19804 6054 20604 6 div[2]
port 10 nsew signal input
rlabel metal2 s 478 0 534 800 6 div[3]
port 11 nsew signal input
rlabel metal2 s 11518 19804 11574 20604 6 div[4]
port 12 nsew signal input
rlabel metal2 s 12898 19804 12954 20604 6 ext_trim[0]
port 13 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 ext_trim[10]
port 14 nsew signal input
rlabel metal2 s 1858 19804 1914 20604 6 ext_trim[11]
port 15 nsew signal input
rlabel metal3 s 17660 4768 18460 4888 6 ext_trim[12]
port 16 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 ext_trim[13]
port 17 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 ext_trim[14]
port 18 nsew signal input
rlabel metal3 s 17660 14968 18460 15088 6 ext_trim[15]
port 19 nsew signal input
rlabel metal2 s 3238 19804 3294 20604 6 ext_trim[16]
port 20 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 ext_trim[17]
port 21 nsew signal input
rlabel metal2 s 4618 19804 4674 20604 6 ext_trim[18]
port 22 nsew signal input
rlabel metal3 s 17660 8848 18460 8968 6 ext_trim[19]
port 23 nsew signal input
rlabel metal2 s 10138 19804 10194 20604 6 ext_trim[1]
port 24 nsew signal input
rlabel metal2 s 8758 19804 8814 20604 6 ext_trim[20]
port 25 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 ext_trim[21]
port 26 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 ext_trim[22]
port 27 nsew signal input
rlabel metal3 s 17660 19048 18460 19168 6 ext_trim[23]
port 28 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 ext_trim[24]
port 29 nsew signal input
rlabel metal2 s 7378 19804 7434 20604 6 ext_trim[25]
port 30 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 ext_trim[2]
port 31 nsew signal input
rlabel metal3 s 17660 6808 18460 6928 6 ext_trim[3]
port 32 nsew signal input
rlabel metal3 s 17660 688 18460 808 6 ext_trim[4]
port 33 nsew signal input
rlabel metal3 s 17660 10888 18460 11008 6 ext_trim[5]
port 34 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 ext_trim[6]
port 35 nsew signal input
rlabel metal2 s 478 19804 534 20604 6 ext_trim[7]
port 36 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 ext_trim[8]
port 37 nsew signal input
rlabel metal3 s 17660 2728 18460 2848 6 ext_trim[9]
port 38 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 extclk_sel
port 39 nsew signal input
rlabel metal2 s 14278 19804 14334 20604 6 osc
port 40 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 reset
port 41 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 sel[0]
port 42 nsew signal input
rlabel metal2 s 17038 19804 17094 20604 6 sel[1]
port 43 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 sel[2]
port 44 nsew signal input
rlabel metal4 s 14437 156 14757 19972 6 VPWR
port 45 nsew power bidirectional
rlabel metal4 s 9040 156 9360 19972 6 VPWR
port 46 nsew power bidirectional
rlabel metal4 s 3643 156 3963 19972 6 VPWR
port 47 nsew power bidirectional
rlabel metal4 s 18336 816 18656 19312 6 VPWR
port 48 nsew power bidirectional
rlabel metal4 s -256 816 64 19312 4 VPWR
port 49 nsew power bidirectional
rlabel metal5 s -256 18992 18656 19312 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s -916 15115 19316 15435 6 VPWR
port 51 nsew power bidirectional
rlabel metal5 s -916 9856 19316 10176 6 VPWR
port 52 nsew power bidirectional
rlabel metal5 s -916 4597 19316 4917 6 VPWR
port 53 nsew power bidirectional
rlabel metal5 s -256 816 18656 1136 6 VPWR
port 54 nsew power bidirectional
rlabel metal4 s 18996 156 19316 19972 6 VGND
port 55 nsew ground bidirectional
rlabel metal4 s 11739 156 12059 19972 6 VGND
port 56 nsew ground bidirectional
rlabel metal4 s 6341 156 6661 19972 6 VGND
port 57 nsew ground bidirectional
rlabel metal4 s -916 156 -596 19972 4 VGND
port 58 nsew ground bidirectional
rlabel metal5 s -916 19652 19316 19972 6 VGND
port 59 nsew ground bidirectional
rlabel metal5 s -916 12485 19316 12805 6 VGND
port 60 nsew ground bidirectional
rlabel metal5 s -916 7227 19316 7547 6 VGND
port 61 nsew ground bidirectional
rlabel metal5 s -916 156 19316 476 6 VGND
port 62 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 18460 20604
<< end >>
