VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_pll
  CLASS BLOCK ;
  FOREIGN digital_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 86.230 BY 96.950 ;
  PIN clockp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END clockp[0]
  PIN clockp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 92.950 55.570 96.950 ;
    END
  END clockp[1]
  PIN div[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 92.950 25.670 96.950 ;
    END
  END div[0]
  PIN div[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END div[1]
  PIN div[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 92.950 83.170 96.950 ;
    END
  END div[2]
  PIN div[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END div[3]
  PIN div[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END div[4]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END enable
  PIN osc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 82.230 6.840 86.230 7.440 ;
    END
  END osc
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 82.230 51.040 86.230 51.640 ;
    END
  END resetb
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 67.205 10.640 68.805 84.560 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 42.210 10.640 43.810 84.560 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 17.215 10.640 18.815 84.560 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 71.040 80.500 72.640 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 46.560 80.500 48.160 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 22.080 80.500 23.680 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 54.705 10.640 56.305 84.560 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 29.715 10.640 31.315 84.560 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 58.800 80.500 60.400 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 34.320 80.500 35.920 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 80.500 84.405 ;
      LAYER met1 ;
        RECT 2.370 10.640 83.190 84.560 ;
      LAYER met2 ;
        RECT 2.400 92.670 25.110 92.950 ;
        RECT 25.950 92.670 55.010 92.950 ;
        RECT 55.850 92.670 82.610 92.950 ;
        RECT 2.400 4.280 83.160 92.670 ;
        RECT 2.950 4.000 29.710 4.280 ;
        RECT 30.550 4.000 59.610 4.280 ;
        RECT 60.450 4.000 83.160 4.280 ;
      LAYER met3 ;
        RECT 4.400 88.040 82.230 88.905 ;
        RECT 4.000 52.040 82.230 88.040 ;
        RECT 4.000 50.640 81.830 52.040 ;
        RECT 4.000 45.240 82.230 50.640 ;
        RECT 4.400 43.840 82.230 45.240 ;
        RECT 4.000 7.840 82.230 43.840 ;
        RECT 4.000 6.975 81.830 7.840 ;
      LAYER met4 ;
        RECT 31.715 10.640 41.810 84.560 ;
        RECT 44.210 10.640 54.305 84.560 ;
        RECT 56.705 10.640 66.805 84.560 ;
  END
END digital_pll
END LIBRARY

