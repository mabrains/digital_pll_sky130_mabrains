magic
tech sky130A
magscale 1 2
timestamp 1620212618
<< locali >>
rect 6285 17119 6319 17221
rect 3709 15419 3743 15521
rect 11529 12631 11563 12733
rect 13829 12087 13863 12257
rect 14105 11067 14139 11169
rect 14473 11135 14507 11305
rect 10425 9503 10459 9673
rect 11529 9503 11563 9605
rect 6193 9367 6227 9469
rect 7205 7939 7239 8041
rect 7665 7735 7699 7973
<< viali >>
rect 1501 17833 1535 17867
rect 16865 17765 16899 17799
rect 1593 17697 1627 17731
rect 1869 17697 1903 17731
rect 2329 17697 2363 17731
rect 3249 17697 3283 17731
rect 4253 17697 4287 17731
rect 4813 17697 4847 17731
rect 6009 17697 6043 17731
rect 7573 17697 7607 17731
rect 8769 17697 8803 17731
rect 9413 17697 9447 17731
rect 10149 17697 10183 17731
rect 11713 17697 11747 17731
rect 12357 17697 12391 17731
rect 12909 17697 12943 17731
rect 14381 17697 14415 17731
rect 14749 17629 14783 17663
rect 15025 17629 15059 17663
rect 6193 17561 6227 17595
rect 9229 17561 9263 17595
rect 2053 17493 2087 17527
rect 2145 17493 2179 17527
rect 3433 17493 3467 17527
rect 4445 17493 4479 17527
rect 4629 17493 4663 17527
rect 7389 17493 7423 17527
rect 8953 17493 8987 17527
rect 10333 17493 10367 17527
rect 11529 17493 11563 17527
rect 12541 17493 12575 17527
rect 13093 17493 13127 17527
rect 14197 17493 14231 17527
rect 16497 17493 16531 17527
rect 16773 17493 16807 17527
rect 1593 17289 1627 17323
rect 2881 17289 2915 17323
rect 15393 17289 15427 17323
rect 15945 17289 15979 17323
rect 6285 17221 6319 17255
rect 9965 17221 9999 17255
rect 3709 17153 3743 17187
rect 5273 17153 5307 17187
rect 8309 17153 8343 17187
rect 11713 17153 11747 17187
rect 13921 17153 13955 17187
rect 1777 17085 1811 17119
rect 2605 17085 2639 17119
rect 2743 17085 2777 17119
rect 2973 17085 3007 17119
rect 3249 17085 3283 17119
rect 3433 17085 3467 17119
rect 5641 17085 5675 17119
rect 6285 17085 6319 17119
rect 6653 17085 6687 17119
rect 6837 17085 6871 17119
rect 7021 17085 7055 17119
rect 8033 17085 8067 17119
rect 10149 17085 10183 17119
rect 10333 17085 10367 17119
rect 10517 17085 10551 17119
rect 13645 17085 13679 17119
rect 15669 17085 15703 17119
rect 15761 17085 15795 17119
rect 16221 17085 16255 17119
rect 16589 17085 16623 17119
rect 5457 17017 5491 17051
rect 6745 17017 6779 17051
rect 10241 17017 10275 17051
rect 11989 17017 12023 17051
rect 16773 17017 16807 17051
rect 2421 16949 2455 16983
rect 3065 16949 3099 16983
rect 5181 16949 5215 16983
rect 6469 16949 6503 16983
rect 9781 16949 9815 16983
rect 13461 16949 13495 16983
rect 15485 16949 15519 16983
rect 16037 16949 16071 16983
rect 3341 16745 3375 16779
rect 8125 16745 8159 16779
rect 14565 16745 14599 16779
rect 1685 16677 1719 16711
rect 6561 16677 6595 16711
rect 10241 16677 10275 16711
rect 10333 16677 10367 16711
rect 11161 16677 11195 16711
rect 11621 16677 11655 16711
rect 3433 16609 3467 16643
rect 4629 16609 4663 16643
rect 8309 16609 8343 16643
rect 10057 16609 10091 16643
rect 10425 16609 10459 16643
rect 10701 16609 10735 16643
rect 11069 16609 11103 16643
rect 11437 16609 11471 16643
rect 11713 16609 11747 16643
rect 14381 16609 14415 16643
rect 16037 16609 16071 16643
rect 16221 16609 16255 16643
rect 16681 16609 16715 16643
rect 16773 16609 16807 16643
rect 1409 16541 1443 16575
rect 6285 16541 6319 16575
rect 10793 16541 10827 16575
rect 11437 16473 11471 16507
rect 3157 16405 3191 16439
rect 4813 16405 4847 16439
rect 8033 16405 8067 16439
rect 10609 16405 10643 16439
rect 15761 16405 15795 16439
rect 16773 16201 16807 16235
rect 5733 16133 5767 16167
rect 4169 16065 4203 16099
rect 10241 16065 10275 16099
rect 10609 16065 10643 16099
rect 10885 16065 10919 16099
rect 15025 16065 15059 16099
rect 15301 16065 15335 16099
rect 1409 15997 1443 16031
rect 3893 15997 3927 16031
rect 5917 15997 5951 16031
rect 6009 15997 6043 16031
rect 6285 15997 6319 16031
rect 6561 15997 6595 16031
rect 6653 15997 6687 16031
rect 7021 15997 7055 16031
rect 7205 15997 7239 16031
rect 7297 15997 7331 16031
rect 9505 15997 9539 16031
rect 9689 15997 9723 16031
rect 9965 15997 9999 16031
rect 10149 15997 10183 16031
rect 10333 15997 10367 16031
rect 10517 15997 10551 16031
rect 10793 15997 10827 16031
rect 12449 15997 12483 16031
rect 6101 15929 6135 15963
rect 12725 15929 12759 15963
rect 1593 15861 1627 15895
rect 5641 15861 5675 15895
rect 9505 15861 9539 15895
rect 9781 15861 9815 15895
rect 11253 15861 11287 15895
rect 14197 15861 14231 15895
rect 3893 15657 3927 15691
rect 10057 15657 10091 15691
rect 13553 15657 13587 15691
rect 16129 15657 16163 15691
rect 3065 15589 3099 15623
rect 8217 15589 8251 15623
rect 8861 15589 8895 15623
rect 10241 15589 10275 15623
rect 2145 15521 2179 15555
rect 3249 15521 3283 15555
rect 3341 15521 3375 15555
rect 3617 15521 3651 15555
rect 3709 15521 3743 15555
rect 3893 15521 3927 15555
rect 4077 15521 4111 15555
rect 4813 15521 4847 15555
rect 7205 15521 7239 15555
rect 7573 15521 7607 15555
rect 8401 15521 8435 15555
rect 8493 15521 8527 15555
rect 9321 15521 9355 15555
rect 10425 15521 10459 15555
rect 11989 15521 12023 15555
rect 12173 15521 12207 15555
rect 12265 15521 12299 15555
rect 12541 15521 12575 15555
rect 12817 15521 12851 15555
rect 13001 15521 13035 15555
rect 13369 15521 13403 15555
rect 14565 15521 14599 15555
rect 16313 15521 16347 15555
rect 7297 15453 7331 15487
rect 7757 15453 7791 15487
rect 8033 15453 8067 15487
rect 8677 15453 8711 15487
rect 8769 15453 8803 15487
rect 12357 15453 12391 15487
rect 12909 15453 12943 15487
rect 3709 15385 3743 15419
rect 4905 15385 4939 15419
rect 7941 15385 7975 15419
rect 1961 15317 1995 15351
rect 3525 15317 3559 15351
rect 9229 15317 9263 15351
rect 12725 15317 12759 15351
rect 14473 15317 14507 15351
rect 1409 15113 1443 15147
rect 7481 15113 7515 15147
rect 15485 15113 15519 15147
rect 7849 15045 7883 15079
rect 9689 15045 9723 15079
rect 4077 14977 4111 15011
rect 7297 14977 7331 15011
rect 7573 14977 7607 15011
rect 9505 14977 9539 15011
rect 14013 14977 14047 15011
rect 14565 14977 14599 15011
rect 15025 14977 15059 15011
rect 3157 14909 3191 14943
rect 3433 14909 3467 14943
rect 3735 14909 3769 14943
rect 3893 14909 3927 14943
rect 3985 14909 4019 14943
rect 5457 14909 5491 14943
rect 6837 14909 6871 14943
rect 7389 14909 7423 14943
rect 7481 14909 7515 14943
rect 8493 14909 8527 14943
rect 8677 14909 8711 14943
rect 8861 14909 8895 14943
rect 8953 14909 8987 14943
rect 9321 14909 9355 14943
rect 9781 14909 9815 14943
rect 10609 14909 10643 14943
rect 10885 14909 10919 14943
rect 10977 14909 11011 14943
rect 14197 14909 14231 14943
rect 14473 14909 14507 14943
rect 14766 14909 14800 14943
rect 14933 14909 14967 14943
rect 15117 14909 15151 14943
rect 15301 14909 15335 14943
rect 15393 14909 15427 14943
rect 15577 14909 15611 14943
rect 16773 14909 16807 14943
rect 2881 14841 2915 14875
rect 3249 14841 3283 14875
rect 3525 14841 3559 14875
rect 3617 14841 3651 14875
rect 7021 14841 7055 14875
rect 7941 14841 7975 14875
rect 9505 14841 9539 14875
rect 10793 14841 10827 14875
rect 5641 14773 5675 14807
rect 11161 14773 11195 14807
rect 14381 14773 14415 14807
rect 16589 14773 16623 14807
rect 3341 14569 3375 14603
rect 4077 14569 4111 14603
rect 7757 14569 7791 14603
rect 10425 14569 10459 14603
rect 10701 14569 10735 14603
rect 2973 14501 3007 14535
rect 3157 14501 3191 14535
rect 12173 14501 12207 14535
rect 12909 14501 12943 14535
rect 15117 14501 15151 14535
rect 15209 14501 15243 14535
rect 1409 14433 1443 14467
rect 3709 14433 3743 14467
rect 3985 14433 4019 14467
rect 4537 14433 4571 14467
rect 7849 14433 7883 14467
rect 10484 14433 10518 14467
rect 12449 14433 12483 14467
rect 12725 14433 12759 14467
rect 12817 14433 12851 14467
rect 13093 14433 13127 14467
rect 13185 14433 13219 14467
rect 14933 14433 14967 14467
rect 15301 14433 15335 14467
rect 3433 14365 3467 14399
rect 3617 14365 3651 14399
rect 4813 14365 4847 14399
rect 9965 14365 9999 14399
rect 10609 14297 10643 14331
rect 1593 14229 1627 14263
rect 3525 14229 3559 14263
rect 6285 14229 6319 14263
rect 10057 14229 10091 14263
rect 12541 14229 12575 14263
rect 15485 14229 15519 14263
rect 5273 14025 5307 14059
rect 8125 14025 8159 14059
rect 8861 14025 8895 14059
rect 14105 14025 14139 14059
rect 14473 14025 14507 14059
rect 9413 13957 9447 13991
rect 10701 13957 10735 13991
rect 6101 13889 6135 13923
rect 8309 13889 8343 13923
rect 8769 13889 8803 13923
rect 9965 13889 9999 13923
rect 10149 13889 10183 13923
rect 12357 13889 12391 13923
rect 12633 13889 12667 13923
rect 15025 13889 15059 13923
rect 15301 13889 15335 13923
rect 16773 13889 16807 13923
rect 3985 13821 4019 13855
rect 4077 13821 4111 13855
rect 5457 13821 5491 13855
rect 5917 13821 5951 13855
rect 6009 13821 6043 13855
rect 6193 13821 6227 13855
rect 8401 13821 8435 13855
rect 9229 13821 9263 13855
rect 9594 13821 9628 13855
rect 10057 13821 10091 13855
rect 10333 13821 10367 13855
rect 10609 13821 10643 13855
rect 10701 13821 10735 13855
rect 10885 13821 10919 13855
rect 14657 13821 14691 13855
rect 14933 13821 14967 13855
rect 5549 13753 5583 13787
rect 5641 13753 5675 13787
rect 5779 13753 5813 13787
rect 9045 13753 9079 13787
rect 10517 13753 10551 13787
rect 9597 13685 9631 13719
rect 14841 13685 14875 13719
rect 6377 13481 6411 13515
rect 10701 13481 10735 13515
rect 12909 13481 12943 13515
rect 13461 13481 13495 13515
rect 16313 13481 16347 13515
rect 3525 13413 3559 13447
rect 4721 13413 4755 13447
rect 6469 13413 6503 13447
rect 13001 13413 13035 13447
rect 2237 13345 2271 13379
rect 3709 13345 3743 13379
rect 4077 13345 4111 13379
rect 4169 13345 4203 13379
rect 4445 13345 4479 13379
rect 4905 13345 4939 13379
rect 6009 13345 6043 13379
rect 6193 13345 6227 13379
rect 6745 13345 6779 13379
rect 7389 13345 7423 13379
rect 7665 13345 7699 13379
rect 10977 13345 11011 13379
rect 11253 13345 11287 13379
rect 11621 13345 11655 13379
rect 12817 13345 12851 13379
rect 13277 13345 13311 13379
rect 14933 13345 14967 13379
rect 15117 13345 15151 13379
rect 15485 13345 15519 13379
rect 15577 13345 15611 13379
rect 16497 13345 16531 13379
rect 4353 13277 4387 13311
rect 6469 13277 6503 13311
rect 6653 13277 6687 13311
rect 10885 13277 10919 13311
rect 11345 13277 11379 13311
rect 15301 13277 15335 13311
rect 4537 13209 4571 13243
rect 7757 13209 7791 13243
rect 12633 13209 12667 13243
rect 2053 13141 2087 13175
rect 3341 13141 3375 13175
rect 3893 13141 3927 13175
rect 7481 13141 7515 13175
rect 11529 13141 11563 13175
rect 13185 13141 13219 13175
rect 10701 12937 10735 12971
rect 11253 12937 11287 12971
rect 11713 12937 11747 12971
rect 12909 12937 12943 12971
rect 14473 12937 14507 12971
rect 14933 12937 14967 12971
rect 16589 12937 16623 12971
rect 4813 12869 4847 12903
rect 5089 12869 5123 12903
rect 7849 12869 7883 12903
rect 3249 12801 3283 12835
rect 4721 12801 4755 12835
rect 7941 12801 7975 12835
rect 8125 12801 8159 12835
rect 8309 12801 8343 12835
rect 3525 12733 3559 12767
rect 3617 12733 3651 12767
rect 3985 12733 4019 12767
rect 4077 12733 4111 12767
rect 4445 12733 4479 12767
rect 4629 12733 4663 12767
rect 4905 12733 4939 12767
rect 6653 12733 6687 12767
rect 6837 12733 6871 12767
rect 7021 12733 7055 12767
rect 7205 12733 7239 12767
rect 7353 12733 7387 12767
rect 7573 12733 7607 12767
rect 7670 12733 7704 12767
rect 8217 12733 8251 12767
rect 10882 12733 10916 12767
rect 11345 12733 11379 12767
rect 11529 12733 11563 12767
rect 11989 12733 12023 12767
rect 12081 12733 12115 12767
rect 12265 12733 12299 12767
rect 13001 12733 13035 12767
rect 14381 12733 14415 12767
rect 14749 12733 14783 12767
rect 14933 12733 14967 12767
rect 15209 12733 15243 12767
rect 15301 12733 15335 12767
rect 16773 12733 16807 12767
rect 2973 12665 3007 12699
rect 3341 12665 3375 12699
rect 3709 12665 3743 12699
rect 3847 12665 3881 12699
rect 4169 12665 4203 12699
rect 6745 12665 6779 12699
rect 7481 12665 7515 12699
rect 7941 12665 7975 12699
rect 8585 12665 8619 12699
rect 11713 12665 11747 12699
rect 12173 12665 12207 12699
rect 1501 12597 1535 12631
rect 6469 12597 6503 12631
rect 10057 12597 10091 12631
rect 10885 12597 10919 12631
rect 11529 12597 11563 12631
rect 11897 12597 11931 12631
rect 7297 12393 7331 12427
rect 9505 12393 9539 12427
rect 9689 12393 9723 12427
rect 13001 12393 13035 12427
rect 15761 12393 15795 12427
rect 3893 12325 3927 12359
rect 14013 12325 14047 12359
rect 15393 12325 15427 12359
rect 1409 12257 1443 12291
rect 4169 12257 4203 12291
rect 4261 12257 4295 12291
rect 6377 12257 6411 12291
rect 6653 12257 6687 12291
rect 6837 12257 6871 12291
rect 7481 12257 7515 12291
rect 7573 12257 7607 12291
rect 7849 12257 7883 12291
rect 9413 12257 9447 12291
rect 9873 12257 9907 12291
rect 13185 12257 13219 12291
rect 13369 12257 13403 12291
rect 13737 12257 13771 12291
rect 13829 12257 13863 12291
rect 13921 12257 13955 12291
rect 15209 12257 15243 12291
rect 15485 12257 15519 12291
rect 15577 12257 15611 12291
rect 3893 12189 3927 12223
rect 4077 12189 4111 12223
rect 6561 12189 6595 12223
rect 6745 12189 6779 12223
rect 10333 12189 10367 12223
rect 10609 12189 10643 12223
rect 13461 12189 13495 12223
rect 13645 12189 13679 12223
rect 1593 12053 1627 12087
rect 4353 12053 4387 12087
rect 7021 12053 7055 12087
rect 7757 12053 7791 12087
rect 12081 12053 12115 12087
rect 13369 12053 13403 12087
rect 13553 12053 13587 12087
rect 13829 12053 13863 12087
rect 13369 11849 13403 11883
rect 15393 11849 15427 11883
rect 16589 11781 16623 11815
rect 12817 11713 12851 11747
rect 12909 11713 12943 11747
rect 13829 11713 13863 11747
rect 4399 11645 4433 11679
rect 4629 11645 4663 11679
rect 4757 11645 4791 11679
rect 4905 11645 4939 11679
rect 5181 11645 5215 11679
rect 6745 11645 6779 11679
rect 6838 11645 6872 11679
rect 7021 11645 7055 11679
rect 7210 11645 7244 11679
rect 7481 11645 7515 11679
rect 9505 11645 9539 11679
rect 12725 11645 12759 11679
rect 13001 11645 13035 11679
rect 13277 11645 13311 11679
rect 13553 11645 13587 11679
rect 13737 11645 13771 11679
rect 13921 11645 13955 11679
rect 14105 11645 14139 11679
rect 14565 11645 14599 11679
rect 15574 11645 15608 11679
rect 15945 11645 15979 11679
rect 16037 11645 16071 11679
rect 16773 11645 16807 11679
rect 4537 11577 4571 11611
rect 7113 11577 7147 11611
rect 7573 11577 7607 11611
rect 14289 11577 14323 11611
rect 14381 11577 14415 11611
rect 4261 11509 4295 11543
rect 5089 11509 5123 11543
rect 7389 11509 7423 11543
rect 9689 11509 9723 11543
rect 13185 11509 13219 11543
rect 14749 11509 14783 11543
rect 15577 11509 15611 11543
rect 2513 11305 2547 11339
rect 5181 11305 5215 11339
rect 6837 11305 6871 11339
rect 7021 11305 7055 11339
rect 10885 11305 10919 11339
rect 11069 11305 11103 11339
rect 14473 11305 14507 11339
rect 15117 11305 15151 11339
rect 16957 11305 16991 11339
rect 1961 11237 1995 11271
rect 7757 11237 7791 11271
rect 9413 11237 9447 11271
rect 11345 11237 11379 11271
rect 11437 11237 11471 11271
rect 11989 11237 12023 11271
rect 13737 11237 13771 11271
rect 1501 11169 1535 11203
rect 2053 11169 2087 11203
rect 4261 11169 4295 11203
rect 4353 11169 4387 11203
rect 5365 11169 5399 11203
rect 5457 11169 5491 11203
rect 5733 11169 5767 11203
rect 6929 11169 6963 11203
rect 7205 11169 7239 11203
rect 7297 11169 7331 11203
rect 7573 11169 7607 11203
rect 8033 11169 8067 11203
rect 11253 11169 11287 11203
rect 11621 11169 11655 11203
rect 14105 11169 14139 11203
rect 2145 11101 2179 11135
rect 4537 11101 4571 11135
rect 7757 11101 7791 11135
rect 7941 11101 7975 11135
rect 9137 11101 9171 11135
rect 14013 11101 14047 11135
rect 14841 11237 14875 11271
rect 15485 11237 15519 11271
rect 14565 11169 14599 11203
rect 14749 11169 14783 11203
rect 14933 11169 14967 11203
rect 14473 11101 14507 11135
rect 15209 11101 15243 11135
rect 2513 11033 2547 11067
rect 5641 11033 5675 11067
rect 7481 11033 7515 11067
rect 14105 11033 14139 11067
rect 4445 10965 4479 10999
rect 2145 10761 2179 10795
rect 3065 10761 3099 10795
rect 7021 10761 7055 10795
rect 11437 10761 11471 10795
rect 12909 10761 12943 10795
rect 16405 10761 16439 10795
rect 1593 10625 1627 10659
rect 1685 10625 1719 10659
rect 4169 10625 4203 10659
rect 4445 10625 4479 10659
rect 8677 10625 8711 10659
rect 8861 10625 8895 10659
rect 14105 10625 14139 10659
rect 15853 10625 15887 10659
rect 2697 10557 2731 10591
rect 6929 10557 6963 10591
rect 10241 10557 10275 10591
rect 11253 10557 11287 10591
rect 13093 10557 13127 10591
rect 13829 10557 13863 10591
rect 16221 10557 16255 10591
rect 2881 10489 2915 10523
rect 1777 10421 1811 10455
rect 3157 10421 3191 10455
rect 5917 10421 5951 10455
rect 8217 10421 8251 10455
rect 8585 10421 8619 10455
rect 10333 10421 10367 10455
rect 1501 10217 1535 10251
rect 3617 10217 3651 10251
rect 5273 10217 5307 10251
rect 7205 10217 7239 10251
rect 9137 10217 9171 10251
rect 14933 10217 14967 10251
rect 1593 10081 1627 10115
rect 2605 10081 2639 10115
rect 3157 10081 3191 10115
rect 4077 10081 4111 10115
rect 5089 10081 5123 10115
rect 6377 10081 6411 10115
rect 6469 10081 6503 10115
rect 7113 10081 7147 10115
rect 9413 10081 9447 10115
rect 9873 10081 9907 10115
rect 14749 10081 14783 10115
rect 3249 10013 3283 10047
rect 6285 10013 6319 10047
rect 6561 10013 6595 10047
rect 3617 9945 3651 9979
rect 3893 9945 3927 9979
rect 9597 9945 9631 9979
rect 2605 9877 2639 9911
rect 6101 9877 6135 9911
rect 9505 9877 9539 9911
rect 9689 9877 9723 9911
rect 2789 9673 2823 9707
rect 6101 9673 6135 9707
rect 8033 9673 8067 9707
rect 10425 9673 10459 9707
rect 5733 9605 5767 9639
rect 7021 9605 7055 9639
rect 8401 9605 8435 9639
rect 1869 9537 1903 9571
rect 1961 9537 1995 9571
rect 7205 9537 7239 9571
rect 8125 9537 8159 9571
rect 11529 9605 11563 9639
rect 11713 9605 11747 9639
rect 11069 9537 11103 9571
rect 12265 9537 12299 9571
rect 12817 9537 12851 9571
rect 12909 9537 12943 9571
rect 15025 9537 15059 9571
rect 15209 9537 15243 9571
rect 1777 9469 1811 9503
rect 3985 9469 4019 9503
rect 4445 9469 4479 9503
rect 5273 9469 5307 9503
rect 6009 9469 6043 9503
rect 6101 9469 6135 9503
rect 6193 9469 6227 9503
rect 6837 9469 6871 9503
rect 6929 9469 6963 9503
rect 7297 9469 7331 9503
rect 7573 9469 7607 9503
rect 7757 9469 7791 9503
rect 7849 9469 7883 9503
rect 8033 9469 8067 9503
rect 9137 9469 9171 9503
rect 9229 9469 9263 9503
rect 9413 9469 9447 9503
rect 10425 9469 10459 9503
rect 10517 9469 10551 9503
rect 10701 9469 10735 9503
rect 11253 9469 11287 9503
rect 11529 9469 11563 9503
rect 12081 9469 12115 9503
rect 16773 9469 16807 9503
rect 2697 9401 2731 9435
rect 6469 9401 6503 9435
rect 6653 9401 6687 9435
rect 9597 9401 9631 9435
rect 15301 9401 15335 9435
rect 1409 9333 1443 9367
rect 4077 9333 4111 9367
rect 5365 9333 5399 9367
rect 6193 9333 6227 9367
rect 10609 9333 10643 9367
rect 11437 9333 11471 9367
rect 12173 9333 12207 9367
rect 13001 9333 13035 9367
rect 13369 9333 13403 9367
rect 15669 9333 15703 9367
rect 16589 9333 16623 9367
rect 5089 9129 5123 9163
rect 5733 9129 5767 9163
rect 11621 9129 11655 9163
rect 11989 9129 12023 9163
rect 12633 9129 12667 9163
rect 14749 9129 14783 9163
rect 16497 9129 16531 9163
rect 5365 9061 5399 9095
rect 8861 9061 8895 9095
rect 10977 9061 11011 9095
rect 12265 9061 12299 9095
rect 15945 9061 15979 9095
rect 2973 8993 3007 9027
rect 5549 8993 5583 9027
rect 8125 8993 8159 9027
rect 8401 8993 8435 9027
rect 9137 8993 9171 9027
rect 9413 8993 9447 9027
rect 9597 8993 9631 9027
rect 9965 8993 9999 9027
rect 10149 8993 10183 9027
rect 10517 8993 10551 9027
rect 10609 8993 10643 9027
rect 10793 8993 10827 9027
rect 12449 8993 12483 9027
rect 13369 8993 13403 9027
rect 13921 8993 13955 9027
rect 14381 8993 14415 9027
rect 15025 8993 15059 9027
rect 15485 8993 15519 9027
rect 16037 8993 16071 9027
rect 16773 8993 16807 9027
rect 5089 8925 5123 8959
rect 5181 8925 5215 8959
rect 8217 8925 8251 8959
rect 9505 8925 9539 8959
rect 11345 8925 11379 8959
rect 11529 8925 11563 8959
rect 13829 8925 13863 8959
rect 16129 8925 16163 8959
rect 9873 8857 9907 8891
rect 14749 8857 14783 8891
rect 14841 8857 14875 8891
rect 16497 8857 16531 8891
rect 16589 8857 16623 8891
rect 2881 8789 2915 8823
rect 4629 8789 4663 8823
rect 9321 8789 9355 8823
rect 5365 8585 5399 8619
rect 10885 8585 10919 8619
rect 2237 8517 2271 8551
rect 3617 8517 3651 8551
rect 3709 8517 3743 8551
rect 6101 8517 6135 8551
rect 8125 8517 8159 8551
rect 9229 8517 9263 8551
rect 13277 8517 13311 8551
rect 1869 8449 1903 8483
rect 4629 8449 4663 8483
rect 4721 8449 4755 8483
rect 5549 8449 5583 8483
rect 5641 8449 5675 8483
rect 5825 8449 5859 8483
rect 6285 8449 6319 8483
rect 7021 8449 7055 8483
rect 7481 8449 7515 8483
rect 7757 8449 7791 8483
rect 7941 8449 7975 8483
rect 8309 8449 8343 8483
rect 9597 8449 9631 8483
rect 11253 8449 11287 8483
rect 11437 8449 11471 8483
rect 13093 8449 13127 8483
rect 2605 8381 2639 8415
rect 3157 8381 3191 8415
rect 3249 8381 3283 8415
rect 3893 8381 3927 8415
rect 5733 8381 5767 8415
rect 6009 8381 6043 8415
rect 6469 8381 6503 8415
rect 6929 8381 6963 8415
rect 7573 8381 7607 8415
rect 7665 8381 7699 8415
rect 8033 8381 8067 8415
rect 9413 8381 9447 8415
rect 9505 8381 9539 8415
rect 9682 8381 9716 8415
rect 12817 8381 12851 8415
rect 12909 8381 12943 8415
rect 13461 8381 13495 8415
rect 13921 8381 13955 8415
rect 16129 8381 16163 8415
rect 1409 8313 1443 8347
rect 1593 8313 1627 8347
rect 2697 8313 2731 8347
rect 6285 8313 6319 8347
rect 6653 8313 6687 8347
rect 6837 8313 6871 8347
rect 8309 8313 8343 8347
rect 11345 8313 11379 8347
rect 14105 8313 14139 8347
rect 15945 8313 15979 8347
rect 2237 8245 2271 8279
rect 3617 8245 3651 8279
rect 4169 8245 4203 8279
rect 4537 8245 4571 8279
rect 12449 8245 12483 8279
rect 7205 8041 7239 8075
rect 7573 8041 7607 8075
rect 15945 8041 15979 8075
rect 1869 7973 1903 8007
rect 5825 7973 5859 8007
rect 6009 7973 6043 8007
rect 7665 7973 7699 8007
rect 15117 7973 15151 8007
rect 15761 7973 15795 8007
rect 1409 7905 1443 7939
rect 1961 7905 1995 7939
rect 6653 7905 6687 7939
rect 6929 7905 6963 7939
rect 7205 7905 7239 7939
rect 7297 7905 7331 7939
rect 7389 7905 7423 7939
rect 5733 7837 5767 7871
rect 6745 7837 6779 7871
rect 6837 7837 6871 7871
rect 7573 7837 7607 7871
rect 6285 7769 6319 7803
rect 7941 7905 7975 7939
rect 9965 7905 9999 7939
rect 15301 7905 15335 7939
rect 15853 7905 15887 7939
rect 15945 7905 15979 7939
rect 9321 7837 9355 7871
rect 16313 7837 16347 7871
rect 14933 7769 14967 7803
rect 6469 7701 6503 7735
rect 7665 7701 7699 7735
rect 7849 7701 7883 7735
rect 2513 7497 2547 7531
rect 8217 7497 8251 7531
rect 8953 7497 8987 7531
rect 6561 7429 6595 7463
rect 10333 7429 10367 7463
rect 14197 7429 14231 7463
rect 3893 7361 3927 7395
rect 6929 7361 6963 7395
rect 7941 7361 7975 7395
rect 8125 7361 8159 7395
rect 9873 7361 9907 7395
rect 13829 7361 13863 7395
rect 4261 7293 4295 7327
rect 7113 7293 7147 7327
rect 8033 7293 8067 7327
rect 8401 7293 8435 7327
rect 10885 7293 10919 7327
rect 11437 7293 11471 7327
rect 12449 7293 12483 7327
rect 12633 7293 12667 7327
rect 13185 7293 13219 7327
rect 13737 7293 13771 7327
rect 2605 7225 2639 7259
rect 4353 7225 4387 7259
rect 5181 7225 5215 7259
rect 7021 7225 7055 7259
rect 8769 7225 8803 7259
rect 8974 7225 9008 7259
rect 9781 7225 9815 7259
rect 9873 7225 9907 7259
rect 10977 7225 11011 7259
rect 13645 7225 13679 7259
rect 4261 7157 4295 7191
rect 4445 7157 4479 7191
rect 5089 7157 5123 7191
rect 8585 7157 8619 7191
rect 9137 7157 9171 7191
rect 12817 7157 12851 7191
rect 14197 7157 14231 7191
rect 1961 6953 1995 6987
rect 5457 6953 5491 6987
rect 8309 6953 8343 6987
rect 10885 6953 10919 6987
rect 13645 6953 13679 6987
rect 16405 6953 16439 6987
rect 4445 6885 4479 6919
rect 4997 6885 5031 6919
rect 12541 6885 12575 6919
rect 12725 6885 12759 6919
rect 13737 6885 13771 6919
rect 1869 6817 1903 6851
rect 3893 6817 3927 6851
rect 4537 6817 4571 6851
rect 5089 6817 5123 6851
rect 5365 6817 5399 6851
rect 5641 6817 5675 6851
rect 7481 6817 7515 6851
rect 7665 6817 7699 6851
rect 7757 6817 7791 6851
rect 9229 6817 9263 6851
rect 9413 6817 9447 6851
rect 9873 6817 9907 6851
rect 10333 6817 10367 6851
rect 10425 6817 10459 6851
rect 11161 6817 11195 6851
rect 11345 6817 11379 6851
rect 12081 6817 12115 6851
rect 16313 6817 16347 6851
rect 16957 6817 16991 6851
rect 1685 6749 1719 6783
rect 5917 6749 5951 6783
rect 8033 6749 8067 6783
rect 8217 6749 8251 6783
rect 9137 6749 9171 6783
rect 10517 6749 10551 6783
rect 12817 6749 12851 6783
rect 13829 6749 13863 6783
rect 4353 6681 4387 6715
rect 5181 6681 5215 6715
rect 8677 6681 8711 6715
rect 10885 6681 10919 6715
rect 12265 6681 12299 6715
rect 13277 6681 13311 6715
rect 16773 6681 16807 6715
rect 2329 6613 2363 6647
rect 5825 6613 5859 6647
rect 7297 6613 7331 6647
rect 9597 6613 9631 6647
rect 7941 6409 7975 6443
rect 10885 6409 10919 6443
rect 11069 6409 11103 6443
rect 15393 6409 15427 6443
rect 15853 6409 15887 6443
rect 1685 6273 1719 6307
rect 5549 6273 5583 6307
rect 7389 6273 7423 6307
rect 8033 6273 8067 6307
rect 15485 6273 15519 6307
rect 1961 6205 1995 6239
rect 3157 6205 3191 6239
rect 3893 6205 3927 6239
rect 5733 6205 5767 6239
rect 6009 6205 6043 6239
rect 7205 6205 7239 6239
rect 7941 6205 7975 6239
rect 10701 6205 10735 6239
rect 10977 6205 11011 6239
rect 13553 6205 13587 6239
rect 14841 6205 14875 6239
rect 15393 6205 15427 6239
rect 15853 6205 15887 6239
rect 2973 6137 3007 6171
rect 5917 6137 5951 6171
rect 13369 6137 13403 6171
rect 1869 6069 1903 6103
rect 2329 6069 2363 6103
rect 6837 6069 6871 6103
rect 7297 6069 7331 6103
rect 8309 6069 8343 6103
rect 1593 5865 1627 5899
rect 12081 5865 12115 5899
rect 15853 5865 15887 5899
rect 4261 5797 4295 5831
rect 1409 5729 1443 5763
rect 4629 5729 4663 5763
rect 4813 5729 4847 5763
rect 10241 5729 10275 5763
rect 12449 5729 12483 5763
rect 15761 5729 15795 5763
rect 11713 5661 11747 5695
rect 12081 5593 12115 5627
rect 12265 5593 12299 5627
rect 10149 5525 10183 5559
rect 12541 5321 12575 5355
rect 12725 5321 12759 5355
rect 13737 5321 13771 5355
rect 2789 5253 2823 5287
rect 2881 5253 2915 5287
rect 11069 5253 11103 5287
rect 11161 5253 11195 5287
rect 15853 5253 15887 5287
rect 15945 5253 15979 5287
rect 4445 5185 4479 5219
rect 7113 5185 7147 5219
rect 7941 5185 7975 5219
rect 9137 5185 9171 5219
rect 10241 5185 10275 5219
rect 12081 5185 12115 5219
rect 13369 5185 13403 5219
rect 14749 5185 14783 5219
rect 1777 5117 1811 5151
rect 2329 5117 2363 5151
rect 2421 5117 2455 5151
rect 3065 5117 3099 5151
rect 5365 5117 5399 5151
rect 5457 5117 5491 5151
rect 6837 5117 6871 5151
rect 8217 5117 8251 5151
rect 9413 5117 9447 5151
rect 10057 5117 10091 5151
rect 10609 5117 10643 5151
rect 10701 5117 10735 5151
rect 11345 5117 11379 5151
rect 11713 5117 11747 5151
rect 12265 5117 12299 5151
rect 12725 5117 12759 5151
rect 13277 5117 13311 5151
rect 13737 5117 13771 5151
rect 13921 5117 13955 5151
rect 14565 5117 14599 5151
rect 14841 5117 14875 5151
rect 15393 5117 15427 5151
rect 15485 5117 15519 5151
rect 16129 5117 16163 5151
rect 2237 5049 2271 5083
rect 5089 5049 5123 5083
rect 8125 5049 8159 5083
rect 12449 5049 12483 5083
rect 13829 5049 13863 5083
rect 14933 5049 14967 5083
rect 2789 4981 2823 5015
rect 6469 4981 6503 5015
rect 6929 4981 6963 5015
rect 8585 4981 8619 5015
rect 9321 4981 9355 5015
rect 9781 4981 9815 5015
rect 11069 4981 11103 5015
rect 15853 4981 15887 5015
rect 2789 4777 2823 4811
rect 14933 4777 14967 4811
rect 15301 4777 15335 4811
rect 16773 4777 16807 4811
rect 2237 4709 2271 4743
rect 2881 4709 2915 4743
rect 4629 4709 4663 4743
rect 4813 4709 4847 4743
rect 6653 4709 6687 4743
rect 7757 4709 7791 4743
rect 1777 4641 1811 4675
rect 2329 4641 2363 4675
rect 4353 4641 4387 4675
rect 4905 4641 4939 4675
rect 5641 4641 5675 4675
rect 5825 4641 5859 4675
rect 6009 4641 6043 4675
rect 6929 4641 6963 4675
rect 7021 4641 7055 4675
rect 7573 4641 7607 4675
rect 7665 4641 7699 4675
rect 8217 4641 8251 4675
rect 8769 4641 8803 4675
rect 9505 4641 9539 4675
rect 11069 4641 11103 4675
rect 16957 4641 16991 4675
rect 2421 4573 2455 4607
rect 4445 4573 4479 4607
rect 7389 4573 7423 4607
rect 9137 4573 9171 4607
rect 10885 4573 10919 4607
rect 14657 4573 14691 4607
rect 14841 4573 14875 4607
rect 2789 4505 2823 4539
rect 2973 4505 3007 4539
rect 4169 4437 4203 4471
rect 8769 4437 8803 4471
rect 9505 4437 9539 4471
rect 7021 4233 7055 4267
rect 12081 4165 12115 4199
rect 1409 4097 1443 4131
rect 6653 4097 6687 4131
rect 12725 4097 12759 4131
rect 13277 4097 13311 4131
rect 14289 4097 14323 4131
rect 4169 4029 4203 4063
rect 7021 4029 7055 4063
rect 7297 4029 7331 4063
rect 13461 4029 13495 4063
rect 13737 4029 13771 4063
rect 13829 4029 13863 4063
rect 14197 4029 14231 4063
rect 1593 3961 1627 3995
rect 4721 3961 4755 3995
rect 12541 3961 12575 3995
rect 7113 3893 7147 3927
rect 12449 3893 12483 3927
rect 13185 3893 13219 3927
rect 14381 3893 14415 3927
rect 3433 3689 3467 3723
rect 9781 3689 9815 3723
rect 11069 3689 11103 3723
rect 13737 3689 13771 3723
rect 3341 3621 3375 3655
rect 6837 3621 6871 3655
rect 8585 3621 8619 3655
rect 10517 3621 10551 3655
rect 12909 3621 12943 3655
rect 3985 3553 4019 3587
rect 6101 3553 6135 3587
rect 7021 3553 7055 3587
rect 8401 3553 8435 3587
rect 10149 3553 10183 3587
rect 10425 3553 10459 3587
rect 10977 3553 11011 3587
rect 11437 3553 11471 3587
rect 13277 3553 13311 3587
rect 13553 3553 13587 3587
rect 13645 3553 13679 3587
rect 16773 3553 16807 3587
rect 5733 3485 5767 3519
rect 6009 3485 6043 3519
rect 7389 3485 7423 3519
rect 7757 3485 7791 3519
rect 9413 3485 9447 3519
rect 11069 3485 11103 3519
rect 13093 3485 13127 3519
rect 14749 3485 14783 3519
rect 15025 3485 15059 3519
rect 9781 3417 9815 3451
rect 9965 3417 9999 3451
rect 7389 3349 7423 3383
rect 7481 3145 7515 3179
rect 8125 3145 8159 3179
rect 9965 3145 9999 3179
rect 10609 3145 10643 3179
rect 10793 3145 10827 3179
rect 12449 3145 12483 3179
rect 13277 3145 13311 3179
rect 14197 3145 14231 3179
rect 15393 3145 15427 3179
rect 16589 3145 16623 3179
rect 8401 3077 8435 3111
rect 16313 3077 16347 3111
rect 1777 3009 1811 3043
rect 2513 3009 2547 3043
rect 6469 3009 6503 3043
rect 7205 3009 7239 3043
rect 8953 3009 8987 3043
rect 9321 3009 9355 3043
rect 9505 3009 9539 3043
rect 11437 3009 11471 3043
rect 13093 3009 13127 3043
rect 13829 3009 13863 3043
rect 15117 3009 15151 3043
rect 1409 2941 1443 2975
rect 1869 2941 1903 2975
rect 2283 2941 2317 2975
rect 2386 2941 2420 2975
rect 4537 2941 4571 2975
rect 7297 2941 7331 2975
rect 7481 2941 7515 2975
rect 8033 2941 8067 2975
rect 8309 2941 8343 2975
rect 8769 2941 8803 2975
rect 9597 2941 9631 2975
rect 10057 2941 10091 2975
rect 10609 2941 10643 2975
rect 12909 2941 12943 2975
rect 13737 2941 13771 2975
rect 14289 2941 14323 2975
rect 15025 2941 15059 2975
rect 15577 2941 15611 2975
rect 16497 2941 16531 2975
rect 16773 2941 16807 2975
rect 2789 2873 2823 2907
rect 8861 2873 8895 2907
rect 12817 2873 12851 2907
rect 13645 2873 13679 2907
rect 1593 2805 1627 2839
rect 11161 2805 11195 2839
rect 11253 2805 11287 2839
rect 14565 2805 14599 2839
rect 14933 2805 14967 2839
rect 1869 2601 1903 2635
rect 2237 2601 2271 2635
rect 7113 2601 7147 2635
rect 7389 2601 7423 2635
rect 9689 2601 9723 2635
rect 10609 2601 10643 2635
rect 10701 2601 10735 2635
rect 13645 2601 13679 2635
rect 14933 2601 14967 2635
rect 1593 2533 1627 2567
rect 8585 2533 8619 2567
rect 14657 2533 14691 2567
rect 16681 2533 16715 2567
rect 1777 2465 1811 2499
rect 2053 2465 2087 2499
rect 2789 2465 2823 2499
rect 4169 2465 4203 2499
rect 4905 2465 4939 2499
rect 5733 2465 5767 2499
rect 6929 2465 6963 2499
rect 7297 2465 7331 2499
rect 8401 2465 8435 2499
rect 9873 2465 9907 2499
rect 11253 2465 11287 2499
rect 12541 2465 12575 2499
rect 13461 2465 13495 2499
rect 13645 2465 13679 2499
rect 13829 2465 13863 2499
rect 14197 2465 14231 2499
rect 16957 2465 16991 2499
rect 12817 2397 12851 2431
rect 14013 2397 14047 2431
rect 14841 2397 14875 2431
rect 1409 2329 1443 2363
rect 2973 2329 3007 2363
rect 5089 2329 5123 2363
rect 11069 2329 11103 2363
rect 4353 2261 4387 2295
rect 5549 2261 5583 2295
<< metal1 >>
rect 1104 17978 17296 18000
rect 1104 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 6571 17978
rect 6623 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 11904 17978
rect 11956 17926 11968 17978
rect 12020 17926 17296 17978
rect 1104 17904 17296 17926
rect 1486 17864 1492 17876
rect 1447 17836 1492 17864
rect 1486 17824 1492 17836
rect 1544 17824 1550 17876
rect 474 17756 480 17808
rect 532 17796 538 17808
rect 532 17768 2360 17796
rect 532 17756 538 17768
rect 1578 17728 1584 17740
rect 1539 17700 1584 17728
rect 1578 17688 1584 17700
rect 1636 17688 1642 17740
rect 1854 17728 1860 17740
rect 1815 17700 1860 17728
rect 1854 17688 1860 17700
rect 1912 17688 1918 17740
rect 2332 17737 2360 17768
rect 8772 17768 12388 17796
rect 2317 17731 2375 17737
rect 2317 17697 2329 17731
rect 2363 17697 2375 17731
rect 3234 17728 3240 17740
rect 3195 17700 3240 17728
rect 2317 17691 2375 17697
rect 3234 17688 3240 17700
rect 3292 17688 3298 17740
rect 4246 17737 4252 17740
rect 4241 17728 4252 17737
rect 4207 17700 4252 17728
rect 4241 17691 4252 17700
rect 4246 17688 4252 17691
rect 4304 17688 4310 17740
rect 4614 17688 4620 17740
rect 4672 17728 4678 17740
rect 4801 17731 4859 17737
rect 4801 17728 4813 17731
rect 4672 17700 4813 17728
rect 4672 17688 4678 17700
rect 4801 17697 4813 17700
rect 4847 17697 4859 17731
rect 5994 17728 6000 17740
rect 5955 17700 6000 17728
rect 4801 17691 4859 17697
rect 5994 17688 6000 17700
rect 6052 17688 6058 17740
rect 7374 17688 7380 17740
rect 7432 17728 7438 17740
rect 7561 17731 7619 17737
rect 7561 17728 7573 17731
rect 7432 17700 7573 17728
rect 7432 17688 7438 17700
rect 7561 17697 7573 17700
rect 7607 17697 7619 17731
rect 7561 17691 7619 17697
rect 8294 17688 8300 17740
rect 8352 17728 8358 17740
rect 8772 17737 8800 17768
rect 12360 17740 12388 17768
rect 16022 17756 16028 17808
rect 16080 17756 16086 17808
rect 16853 17799 16911 17805
rect 16853 17765 16865 17799
rect 16899 17796 16911 17799
rect 17034 17796 17040 17808
rect 16899 17768 17040 17796
rect 16899 17765 16911 17768
rect 16853 17759 16911 17765
rect 17034 17756 17040 17768
rect 17092 17756 17098 17808
rect 8757 17731 8815 17737
rect 8757 17728 8769 17731
rect 8352 17700 8769 17728
rect 8352 17688 8358 17700
rect 8757 17697 8769 17700
rect 8803 17697 8815 17731
rect 8757 17691 8815 17697
rect 8846 17688 8852 17740
rect 8904 17728 8910 17740
rect 9401 17731 9459 17737
rect 9401 17728 9413 17731
rect 8904 17700 9413 17728
rect 8904 17688 8910 17700
rect 9401 17697 9413 17700
rect 9447 17697 9459 17731
rect 10134 17728 10140 17740
rect 10095 17700 10140 17728
rect 9401 17691 9459 17697
rect 10134 17688 10140 17700
rect 10192 17688 10198 17740
rect 11514 17688 11520 17740
rect 11572 17728 11578 17740
rect 11701 17731 11759 17737
rect 11701 17728 11713 17731
rect 11572 17700 11713 17728
rect 11572 17688 11578 17700
rect 11701 17697 11713 17700
rect 11747 17697 11759 17731
rect 12342 17728 12348 17740
rect 12255 17700 12348 17728
rect 11701 17691 11759 17697
rect 12342 17688 12348 17700
rect 12400 17688 12406 17740
rect 12894 17728 12900 17740
rect 12855 17700 12900 17728
rect 12894 17688 12900 17700
rect 12952 17688 12958 17740
rect 14274 17688 14280 17740
rect 14332 17728 14338 17740
rect 14369 17731 14427 17737
rect 14369 17728 14381 17731
rect 14332 17700 14381 17728
rect 14332 17688 14338 17700
rect 14369 17697 14381 17700
rect 14415 17697 14427 17731
rect 14369 17691 14427 17697
rect 13446 17620 13452 17672
rect 13504 17660 13510 17672
rect 14737 17663 14795 17669
rect 14737 17660 14749 17663
rect 13504 17632 14749 17660
rect 13504 17620 13510 17632
rect 14737 17629 14749 17632
rect 14783 17629 14795 17663
rect 14737 17623 14795 17629
rect 15013 17663 15071 17669
rect 15013 17629 15025 17663
rect 15059 17660 15071 17663
rect 15378 17660 15384 17672
rect 15059 17632 15384 17660
rect 15059 17629 15071 17632
rect 15013 17623 15071 17629
rect 15378 17620 15384 17632
rect 15436 17620 15442 17672
rect 6181 17595 6239 17601
rect 6181 17561 6193 17595
rect 6227 17592 6239 17595
rect 7558 17592 7564 17604
rect 6227 17564 7564 17592
rect 6227 17561 6239 17564
rect 6181 17555 6239 17561
rect 7558 17552 7564 17564
rect 7616 17552 7622 17604
rect 8570 17552 8576 17604
rect 8628 17592 8634 17604
rect 9217 17595 9275 17601
rect 9217 17592 9229 17595
rect 8628 17564 9229 17592
rect 8628 17552 8634 17564
rect 9217 17561 9229 17564
rect 9263 17561 9275 17595
rect 9217 17555 9275 17561
rect 2038 17524 2044 17536
rect 1999 17496 2044 17524
rect 2038 17484 2044 17496
rect 2096 17484 2102 17536
rect 2133 17527 2191 17533
rect 2133 17493 2145 17527
rect 2179 17524 2191 17527
rect 2222 17524 2228 17536
rect 2179 17496 2228 17524
rect 2179 17493 2191 17496
rect 2133 17487 2191 17493
rect 2222 17484 2228 17496
rect 2280 17484 2286 17536
rect 3234 17484 3240 17536
rect 3292 17524 3298 17536
rect 3421 17527 3479 17533
rect 3421 17524 3433 17527
rect 3292 17496 3433 17524
rect 3292 17484 3298 17496
rect 3421 17493 3433 17496
rect 3467 17493 3479 17527
rect 4430 17524 4436 17536
rect 4391 17496 4436 17524
rect 3421 17487 3479 17493
rect 4430 17484 4436 17496
rect 4488 17484 4494 17536
rect 4522 17484 4528 17536
rect 4580 17524 4586 17536
rect 4617 17527 4675 17533
rect 4617 17524 4629 17527
rect 4580 17496 4629 17524
rect 4580 17484 4586 17496
rect 4617 17493 4629 17496
rect 4663 17493 4675 17527
rect 4617 17487 4675 17493
rect 7098 17484 7104 17536
rect 7156 17524 7162 17536
rect 7377 17527 7435 17533
rect 7377 17524 7389 17527
rect 7156 17496 7389 17524
rect 7156 17484 7162 17496
rect 7377 17493 7389 17496
rect 7423 17493 7435 17527
rect 8938 17524 8944 17536
rect 8899 17496 8944 17524
rect 7377 17487 7435 17493
rect 8938 17484 8944 17496
rect 8996 17484 9002 17536
rect 9858 17484 9864 17536
rect 9916 17524 9922 17536
rect 10321 17527 10379 17533
rect 10321 17524 10333 17527
rect 9916 17496 10333 17524
rect 9916 17484 9922 17496
rect 10321 17493 10333 17496
rect 10367 17493 10379 17527
rect 10321 17487 10379 17493
rect 10410 17484 10416 17536
rect 10468 17524 10474 17536
rect 11517 17527 11575 17533
rect 11517 17524 11529 17527
rect 10468 17496 11529 17524
rect 10468 17484 10474 17496
rect 11517 17493 11529 17496
rect 11563 17493 11575 17527
rect 12526 17524 12532 17536
rect 12487 17496 12532 17524
rect 11517 17487 11575 17493
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 13081 17527 13139 17533
rect 13081 17493 13093 17527
rect 13127 17524 13139 17527
rect 13170 17524 13176 17536
rect 13127 17496 13176 17524
rect 13127 17493 13139 17496
rect 13081 17487 13139 17493
rect 13170 17484 13176 17496
rect 13228 17484 13234 17536
rect 13906 17484 13912 17536
rect 13964 17524 13970 17536
rect 14185 17527 14243 17533
rect 14185 17524 14197 17527
rect 13964 17496 14197 17524
rect 13964 17484 13970 17496
rect 14185 17493 14197 17496
rect 14231 17493 14243 17527
rect 14185 17487 14243 17493
rect 16298 17484 16304 17536
rect 16356 17524 16362 17536
rect 16485 17527 16543 17533
rect 16485 17524 16497 17527
rect 16356 17496 16497 17524
rect 16356 17484 16362 17496
rect 16485 17493 16497 17496
rect 16531 17493 16543 17527
rect 16485 17487 16543 17493
rect 16761 17527 16819 17533
rect 16761 17493 16773 17527
rect 16807 17524 16819 17527
rect 16850 17524 16856 17536
rect 16807 17496 16856 17524
rect 16807 17493 16819 17496
rect 16761 17487 16819 17493
rect 16850 17484 16856 17496
rect 16908 17484 16914 17536
rect 1104 17434 17296 17456
rect 1104 17382 3680 17434
rect 3732 17382 3744 17434
rect 3796 17382 3808 17434
rect 3860 17382 3872 17434
rect 3924 17382 9078 17434
rect 9130 17382 9142 17434
rect 9194 17382 9206 17434
rect 9258 17382 9270 17434
rect 9322 17382 14475 17434
rect 14527 17382 14539 17434
rect 14591 17382 14603 17434
rect 14655 17382 14667 17434
rect 14719 17382 17296 17434
rect 1104 17360 17296 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 2774 17280 2780 17332
rect 2832 17320 2838 17332
rect 2869 17323 2927 17329
rect 2869 17320 2881 17323
rect 2832 17292 2881 17320
rect 2832 17280 2838 17292
rect 2869 17289 2881 17292
rect 2915 17289 2927 17323
rect 4246 17320 4252 17332
rect 2869 17283 2927 17289
rect 3344 17292 4252 17320
rect 2130 17144 2136 17196
rect 2188 17184 2194 17196
rect 3344 17184 3372 17292
rect 4246 17280 4252 17292
rect 4304 17280 4310 17332
rect 15378 17320 15384 17332
rect 15339 17292 15384 17320
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 15933 17323 15991 17329
rect 15933 17289 15945 17323
rect 15979 17320 15991 17323
rect 16022 17320 16028 17332
rect 15979 17292 16028 17320
rect 15979 17289 15991 17292
rect 15933 17283 15991 17289
rect 16022 17280 16028 17292
rect 16080 17280 16086 17332
rect 6273 17255 6331 17261
rect 6273 17221 6285 17255
rect 6319 17252 6331 17255
rect 9953 17255 10011 17261
rect 6319 17224 7052 17252
rect 6319 17221 6331 17224
rect 6273 17215 6331 17221
rect 2188 17156 3372 17184
rect 3697 17187 3755 17193
rect 2188 17144 2194 17156
rect 1762 17116 1768 17128
rect 1723 17088 1768 17116
rect 1762 17076 1768 17088
rect 1820 17076 1826 17128
rect 2590 17116 2596 17128
rect 2551 17088 2596 17116
rect 2590 17076 2596 17088
rect 2648 17076 2654 17128
rect 2731 17119 2789 17125
rect 2731 17085 2743 17119
rect 2777 17116 2789 17119
rect 2866 17116 2872 17128
rect 2777 17088 2872 17116
rect 2777 17085 2789 17088
rect 2731 17079 2789 17085
rect 2866 17076 2872 17088
rect 2924 17076 2930 17128
rect 3252 17125 3280 17156
rect 3697 17153 3709 17187
rect 3743 17184 3755 17187
rect 5261 17187 5319 17193
rect 5261 17184 5273 17187
rect 3743 17156 5273 17184
rect 3743 17153 3755 17156
rect 3697 17147 3755 17153
rect 5261 17153 5273 17156
rect 5307 17153 5319 17187
rect 6730 17184 6736 17196
rect 5261 17147 5319 17153
rect 5460 17156 6736 17184
rect 2961 17119 3019 17125
rect 2961 17085 2973 17119
rect 3007 17085 3019 17119
rect 2961 17079 3019 17085
rect 3237 17119 3295 17125
rect 3237 17085 3249 17119
rect 3283 17085 3295 17119
rect 3418 17116 3424 17128
rect 3379 17088 3424 17116
rect 3237 17079 3295 17085
rect 2976 17048 3004 17079
rect 3418 17076 3424 17088
rect 3476 17076 3482 17128
rect 2976 17020 3464 17048
rect 3436 16992 3464 17020
rect 4430 17008 4436 17060
rect 4488 17008 4494 17060
rect 5460 17057 5488 17156
rect 6730 17144 6736 17156
rect 6788 17184 6794 17196
rect 6788 17156 6868 17184
rect 6788 17144 6794 17156
rect 6840 17125 6868 17156
rect 7024 17128 7052 17224
rect 9953 17221 9965 17255
rect 9999 17221 10011 17255
rect 10962 17252 10968 17264
rect 9953 17215 10011 17221
rect 10244 17224 10968 17252
rect 8297 17187 8355 17193
rect 8297 17153 8309 17187
rect 8343 17184 8355 17187
rect 9968 17184 9996 17215
rect 8343 17156 9996 17184
rect 8343 17153 8355 17156
rect 8297 17147 8355 17153
rect 5629 17119 5687 17125
rect 5629 17085 5641 17119
rect 5675 17116 5687 17119
rect 6273 17119 6331 17125
rect 6273 17116 6285 17119
rect 5675 17088 6285 17116
rect 5675 17085 5687 17088
rect 5629 17079 5687 17085
rect 6273 17085 6285 17088
rect 6319 17085 6331 17119
rect 6273 17079 6331 17085
rect 6641 17119 6699 17125
rect 6641 17085 6653 17119
rect 6687 17085 6699 17119
rect 6641 17079 6699 17085
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17085 6883 17119
rect 7006 17116 7012 17128
rect 6967 17088 7012 17116
rect 6825 17079 6883 17085
rect 5445 17051 5503 17057
rect 5445 17017 5457 17051
rect 5491 17017 5503 17051
rect 5445 17011 5503 17017
rect 1670 16940 1676 16992
rect 1728 16980 1734 16992
rect 2409 16983 2467 16989
rect 2409 16980 2421 16983
rect 1728 16952 2421 16980
rect 1728 16940 1734 16952
rect 2409 16949 2421 16952
rect 2455 16949 2467 16983
rect 3050 16980 3056 16992
rect 3011 16952 3056 16980
rect 2409 16943 2467 16949
rect 3050 16940 3056 16952
rect 3108 16940 3114 16992
rect 3418 16940 3424 16992
rect 3476 16940 3482 16992
rect 5169 16983 5227 16989
rect 5169 16949 5181 16983
rect 5215 16980 5227 16983
rect 5460 16980 5488 17011
rect 5215 16952 5488 16980
rect 5215 16949 5227 16952
rect 5169 16943 5227 16949
rect 6270 16940 6276 16992
rect 6328 16980 6334 16992
rect 6457 16983 6515 16989
rect 6457 16980 6469 16983
rect 6328 16952 6469 16980
rect 6328 16940 6334 16952
rect 6457 16949 6469 16952
rect 6503 16949 6515 16983
rect 6656 16980 6684 17079
rect 7006 17076 7012 17088
rect 7064 17076 7070 17128
rect 8018 17116 8024 17128
rect 7979 17088 8024 17116
rect 8018 17076 8024 17088
rect 8076 17076 8082 17128
rect 10137 17119 10195 17125
rect 10137 17085 10149 17119
rect 10183 17116 10195 17119
rect 10244 17116 10272 17224
rect 10962 17212 10968 17224
rect 11020 17212 11026 17264
rect 15654 17212 15660 17264
rect 15712 17212 15718 17264
rect 11701 17187 11759 17193
rect 11701 17153 11713 17187
rect 11747 17184 11759 17187
rect 13906 17184 13912 17196
rect 11747 17156 13492 17184
rect 13867 17156 13912 17184
rect 11747 17153 11759 17156
rect 11701 17147 11759 17153
rect 13464 17128 13492 17156
rect 13906 17144 13912 17156
rect 13964 17144 13970 17196
rect 15672 17184 15700 17212
rect 15672 17156 16252 17184
rect 10183 17088 10272 17116
rect 10183 17085 10195 17088
rect 10137 17079 10195 17085
rect 10318 17076 10324 17128
rect 10376 17116 10382 17128
rect 10376 17088 10421 17116
rect 10376 17076 10382 17088
rect 10502 17076 10508 17128
rect 10560 17116 10566 17128
rect 11422 17116 11428 17128
rect 10560 17088 11428 17116
rect 10560 17076 10566 17088
rect 11422 17076 11428 17088
rect 11480 17076 11486 17128
rect 13446 17076 13452 17128
rect 13504 17116 13510 17128
rect 13633 17119 13691 17125
rect 13633 17116 13645 17119
rect 13504 17088 13645 17116
rect 13504 17076 13510 17088
rect 13633 17085 13645 17088
rect 13679 17085 13691 17119
rect 13633 17079 13691 17085
rect 15562 17076 15568 17128
rect 15620 17116 15626 17128
rect 15657 17119 15715 17125
rect 15657 17116 15669 17119
rect 15620 17088 15669 17116
rect 15620 17076 15626 17088
rect 15657 17085 15669 17088
rect 15703 17085 15715 17119
rect 15657 17079 15715 17085
rect 15746 17076 15752 17128
rect 15804 17116 15810 17128
rect 16224 17125 16252 17156
rect 16209 17119 16267 17125
rect 15804 17088 15849 17116
rect 15804 17076 15810 17088
rect 16209 17085 16221 17119
rect 16255 17085 16267 17119
rect 16209 17079 16267 17085
rect 16577 17119 16635 17125
rect 16577 17085 16589 17119
rect 16623 17116 16635 17119
rect 17034 17116 17040 17128
rect 16623 17088 17040 17116
rect 16623 17085 16635 17088
rect 16577 17079 16635 17085
rect 17034 17076 17040 17088
rect 17092 17076 17098 17128
rect 6733 17051 6791 17057
rect 6733 17017 6745 17051
rect 6779 17048 6791 17051
rect 7282 17048 7288 17060
rect 6779 17020 7288 17048
rect 6779 17017 6791 17020
rect 6733 17011 6791 17017
rect 7282 17008 7288 17020
rect 7340 17008 7346 17060
rect 8938 17008 8944 17060
rect 8996 17008 9002 17060
rect 10229 17051 10287 17057
rect 10229 17048 10241 17051
rect 9784 17020 10241 17048
rect 6822 16980 6828 16992
rect 6656 16952 6828 16980
rect 6457 16943 6515 16949
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 9784 16989 9812 17020
rect 10229 17017 10241 17020
rect 10275 17017 10287 17051
rect 10229 17011 10287 17017
rect 9769 16983 9827 16989
rect 9769 16949 9781 16983
rect 9815 16949 9827 16983
rect 10244 16980 10272 17011
rect 11514 17008 11520 17060
rect 11572 17048 11578 17060
rect 11977 17051 12035 17057
rect 11977 17048 11989 17051
rect 11572 17020 11989 17048
rect 11572 17008 11578 17020
rect 11977 17017 11989 17020
rect 12023 17017 12035 17051
rect 11977 17011 12035 17017
rect 12526 17008 12532 17060
rect 12584 17008 12590 17060
rect 14550 17008 14556 17060
rect 14608 17008 14614 17060
rect 16758 17048 16764 17060
rect 16719 17020 16764 17048
rect 16758 17008 16764 17020
rect 16816 17008 16822 17060
rect 10594 16980 10600 16992
rect 10244 16952 10600 16980
rect 9769 16943 9827 16949
rect 10594 16940 10600 16952
rect 10652 16940 10658 16992
rect 12618 16940 12624 16992
rect 12676 16980 12682 16992
rect 13449 16983 13507 16989
rect 13449 16980 13461 16983
rect 12676 16952 13461 16980
rect 12676 16940 12682 16952
rect 13449 16949 13461 16952
rect 13495 16949 13507 16983
rect 15470 16980 15476 16992
rect 15431 16952 15476 16980
rect 13449 16943 13507 16949
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 15562 16940 15568 16992
rect 15620 16980 15626 16992
rect 16025 16983 16083 16989
rect 16025 16980 16037 16983
rect 15620 16952 16037 16980
rect 15620 16940 15626 16952
rect 16025 16949 16037 16952
rect 16071 16949 16083 16983
rect 16025 16943 16083 16949
rect 1104 16890 17296 16912
rect 1104 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 6571 16890
rect 6623 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 11904 16890
rect 11956 16838 11968 16890
rect 12020 16838 17296 16890
rect 1104 16816 17296 16838
rect 2590 16736 2596 16788
rect 2648 16776 2654 16788
rect 3329 16779 3387 16785
rect 3329 16776 3341 16779
rect 2648 16748 3341 16776
rect 2648 16736 2654 16748
rect 3329 16745 3341 16748
rect 3375 16745 3387 16779
rect 3329 16739 3387 16745
rect 4246 16736 4252 16788
rect 4304 16776 4310 16788
rect 5442 16776 5448 16788
rect 4304 16748 5448 16776
rect 4304 16736 4310 16748
rect 1670 16708 1676 16720
rect 1631 16680 1676 16708
rect 1670 16668 1676 16680
rect 1728 16668 1734 16720
rect 3050 16708 3056 16720
rect 2898 16680 3056 16708
rect 3050 16668 3056 16680
rect 3108 16668 3114 16720
rect 3418 16640 3424 16652
rect 3379 16612 3424 16640
rect 3418 16600 3424 16612
rect 3476 16600 3482 16652
rect 4632 16649 4660 16748
rect 5442 16736 5448 16748
rect 5500 16776 5506 16788
rect 7834 16776 7840 16788
rect 5500 16748 7840 16776
rect 5500 16736 5506 16748
rect 7834 16736 7840 16748
rect 7892 16736 7898 16788
rect 8113 16779 8171 16785
rect 8113 16745 8125 16779
rect 8159 16745 8171 16779
rect 14550 16776 14556 16788
rect 8113 16739 8171 16745
rect 10244 16748 11192 16776
rect 14511 16748 14556 16776
rect 6270 16668 6276 16720
rect 6328 16708 6334 16720
rect 6549 16711 6607 16717
rect 6549 16708 6561 16711
rect 6328 16680 6561 16708
rect 6328 16668 6334 16680
rect 6549 16677 6561 16680
rect 6595 16677 6607 16711
rect 8128 16708 8156 16739
rect 7774 16680 8156 16708
rect 6549 16671 6607 16677
rect 9950 16668 9956 16720
rect 10008 16708 10014 16720
rect 10244 16717 10272 16748
rect 10229 16711 10287 16717
rect 10229 16708 10241 16711
rect 10008 16680 10241 16708
rect 10008 16668 10014 16680
rect 10229 16677 10241 16680
rect 10275 16677 10287 16711
rect 10229 16671 10287 16677
rect 10318 16668 10324 16720
rect 10376 16708 10382 16720
rect 11164 16717 11192 16748
rect 14550 16736 14556 16748
rect 14608 16736 14614 16788
rect 11149 16711 11207 16717
rect 10376 16680 11100 16708
rect 10376 16668 10382 16680
rect 4617 16643 4675 16649
rect 4617 16609 4629 16643
rect 4663 16609 4675 16643
rect 4617 16603 4675 16609
rect 7834 16600 7840 16652
rect 7892 16640 7898 16652
rect 8294 16640 8300 16652
rect 7892 16612 8300 16640
rect 7892 16600 7898 16612
rect 8294 16600 8300 16612
rect 8352 16600 8358 16652
rect 10045 16643 10103 16649
rect 10045 16609 10057 16643
rect 10091 16609 10103 16643
rect 10045 16603 10103 16609
rect 10413 16643 10471 16649
rect 10413 16609 10425 16643
rect 10459 16640 10471 16643
rect 10594 16640 10600 16652
rect 10459 16612 10600 16640
rect 10459 16609 10471 16612
rect 10413 16603 10471 16609
rect 1397 16575 1455 16581
rect 1397 16541 1409 16575
rect 1443 16572 1455 16575
rect 1762 16572 1768 16584
rect 1443 16544 1768 16572
rect 1443 16541 1455 16544
rect 1397 16535 1455 16541
rect 1762 16532 1768 16544
rect 1820 16572 1826 16584
rect 3510 16572 3516 16584
rect 1820 16544 3516 16572
rect 1820 16532 1826 16544
rect 3510 16532 3516 16544
rect 3568 16532 3574 16584
rect 6273 16575 6331 16581
rect 6273 16541 6285 16575
rect 6319 16572 6331 16575
rect 8018 16572 8024 16584
rect 6319 16544 8024 16572
rect 6319 16541 6331 16544
rect 6273 16535 6331 16541
rect 8018 16532 8024 16544
rect 8076 16532 8082 16584
rect 10060 16572 10088 16603
rect 10594 16600 10600 16612
rect 10652 16640 10658 16652
rect 11072 16649 11100 16680
rect 11149 16677 11161 16711
rect 11195 16708 11207 16711
rect 11609 16711 11667 16717
rect 11609 16708 11621 16711
rect 11195 16680 11621 16708
rect 11195 16677 11207 16680
rect 11149 16671 11207 16677
rect 11609 16677 11621 16680
rect 11655 16677 11667 16711
rect 11609 16671 11667 16677
rect 16224 16680 16804 16708
rect 10689 16643 10747 16649
rect 10689 16640 10701 16643
rect 10652 16612 10701 16640
rect 10652 16600 10658 16612
rect 10689 16609 10701 16612
rect 10735 16609 10747 16643
rect 10689 16603 10747 16609
rect 11057 16643 11115 16649
rect 11057 16609 11069 16643
rect 11103 16609 11115 16643
rect 11422 16640 11428 16652
rect 11383 16612 11428 16640
rect 11057 16603 11115 16609
rect 10134 16572 10140 16584
rect 10047 16544 10140 16572
rect 10134 16532 10140 16544
rect 10192 16572 10198 16584
rect 10781 16575 10839 16581
rect 10781 16572 10793 16575
rect 10192 16544 10793 16572
rect 10192 16532 10198 16544
rect 10781 16541 10793 16544
rect 10827 16541 10839 16575
rect 10781 16535 10839 16541
rect 3145 16439 3203 16445
rect 3145 16405 3157 16439
rect 3191 16436 3203 16439
rect 3418 16436 3424 16448
rect 3191 16408 3424 16436
rect 3191 16405 3203 16408
rect 3145 16399 3203 16405
rect 3418 16396 3424 16408
rect 3476 16396 3482 16448
rect 4798 16436 4804 16448
rect 4759 16408 4804 16436
rect 4798 16396 4804 16408
rect 4856 16396 4862 16448
rect 7282 16396 7288 16448
rect 7340 16436 7346 16448
rect 8021 16439 8079 16445
rect 8021 16436 8033 16439
rect 7340 16408 8033 16436
rect 7340 16396 7346 16408
rect 8021 16405 8033 16408
rect 8067 16405 8079 16439
rect 8021 16399 8079 16405
rect 10597 16439 10655 16445
rect 10597 16405 10609 16439
rect 10643 16436 10655 16439
rect 10686 16436 10692 16448
rect 10643 16408 10692 16436
rect 10643 16405 10655 16408
rect 10597 16399 10655 16405
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 11072 16436 11100 16603
rect 11422 16600 11428 16612
rect 11480 16600 11486 16652
rect 11514 16600 11520 16652
rect 11572 16600 11578 16652
rect 11701 16643 11759 16649
rect 11701 16609 11713 16643
rect 11747 16640 11759 16643
rect 12250 16640 12256 16652
rect 11747 16612 12256 16640
rect 11747 16609 11759 16612
rect 11701 16603 11759 16609
rect 12250 16600 12256 16612
rect 12308 16600 12314 16652
rect 12342 16600 12348 16652
rect 12400 16640 12406 16652
rect 13354 16640 13360 16652
rect 12400 16612 13360 16640
rect 12400 16600 12406 16612
rect 13354 16600 13360 16612
rect 13412 16640 13418 16652
rect 14369 16643 14427 16649
rect 14369 16640 14381 16643
rect 13412 16612 14381 16640
rect 13412 16600 13418 16612
rect 14369 16609 14381 16612
rect 14415 16640 14427 16643
rect 15746 16640 15752 16652
rect 14415 16612 15752 16640
rect 14415 16609 14427 16612
rect 14369 16603 14427 16609
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 16022 16640 16028 16652
rect 15983 16612 16028 16640
rect 16022 16600 16028 16612
rect 16080 16600 16086 16652
rect 16224 16649 16252 16680
rect 16776 16652 16804 16680
rect 16209 16643 16267 16649
rect 16209 16609 16221 16643
rect 16255 16609 16267 16643
rect 16209 16603 16267 16609
rect 16298 16600 16304 16652
rect 16356 16640 16362 16652
rect 16669 16643 16727 16649
rect 16669 16640 16681 16643
rect 16356 16612 16681 16640
rect 16356 16600 16362 16612
rect 16669 16609 16681 16612
rect 16715 16609 16727 16643
rect 16669 16603 16727 16609
rect 16758 16600 16764 16652
rect 16816 16640 16822 16652
rect 16816 16612 16909 16640
rect 16816 16600 16822 16612
rect 11425 16507 11483 16513
rect 11425 16473 11437 16507
rect 11471 16504 11483 16507
rect 11532 16504 11560 16600
rect 11606 16532 11612 16584
rect 11664 16572 11670 16584
rect 12360 16572 12388 16600
rect 11664 16544 12388 16572
rect 11664 16532 11670 16544
rect 11471 16476 11560 16504
rect 11471 16473 11483 16476
rect 11425 16467 11483 16473
rect 12618 16436 12624 16448
rect 11072 16408 12624 16436
rect 12618 16396 12624 16408
rect 12676 16396 12682 16448
rect 15378 16396 15384 16448
rect 15436 16436 15442 16448
rect 15749 16439 15807 16445
rect 15749 16436 15761 16439
rect 15436 16408 15761 16436
rect 15436 16396 15442 16408
rect 15749 16405 15761 16408
rect 15795 16405 15807 16439
rect 15749 16399 15807 16405
rect 1104 16346 17296 16368
rect 1104 16294 3680 16346
rect 3732 16294 3744 16346
rect 3796 16294 3808 16346
rect 3860 16294 3872 16346
rect 3924 16294 9078 16346
rect 9130 16294 9142 16346
rect 9194 16294 9206 16346
rect 9258 16294 9270 16346
rect 9322 16294 14475 16346
rect 14527 16294 14539 16346
rect 14591 16294 14603 16346
rect 14655 16294 14667 16346
rect 14719 16294 17296 16346
rect 1104 16272 17296 16294
rect 7006 16232 7012 16244
rect 5920 16204 7012 16232
rect 5721 16167 5779 16173
rect 5721 16133 5733 16167
rect 5767 16133 5779 16167
rect 5721 16127 5779 16133
rect 4157 16099 4215 16105
rect 4157 16065 4169 16099
rect 4203 16096 4215 16099
rect 5736 16096 5764 16127
rect 4203 16068 5764 16096
rect 4203 16065 4215 16068
rect 4157 16059 4215 16065
rect 1394 16028 1400 16040
rect 1355 16000 1400 16028
rect 1394 15988 1400 16000
rect 1452 15988 1458 16040
rect 3510 15988 3516 16040
rect 3568 16028 3574 16040
rect 5920 16037 5948 16204
rect 7006 16192 7012 16204
rect 7064 16192 7070 16244
rect 16758 16232 16764 16244
rect 16719 16204 16764 16232
rect 16758 16192 16764 16204
rect 16816 16192 16822 16244
rect 7282 16164 7288 16176
rect 6012 16136 7288 16164
rect 6012 16037 6040 16136
rect 7282 16124 7288 16136
rect 7340 16124 7346 16176
rect 10410 16164 10416 16176
rect 9508 16136 10416 16164
rect 6730 16096 6736 16108
rect 6564 16068 6736 16096
rect 3881 16031 3939 16037
rect 3881 16028 3893 16031
rect 3568 16000 3893 16028
rect 3568 15988 3574 16000
rect 3881 15997 3893 16000
rect 3927 15997 3939 16031
rect 3881 15991 3939 15997
rect 5905 16031 5963 16037
rect 5905 15997 5917 16031
rect 5951 15997 5963 16031
rect 5905 15991 5963 15997
rect 5997 16031 6055 16037
rect 5997 15997 6009 16031
rect 6043 15997 6055 16031
rect 5997 15991 6055 15997
rect 6273 16031 6331 16037
rect 6273 15997 6285 16031
rect 6319 16028 6331 16031
rect 6454 16028 6460 16040
rect 6319 16000 6460 16028
rect 6319 15997 6331 16000
rect 6273 15991 6331 15997
rect 3896 15960 3924 15991
rect 6454 15988 6460 16000
rect 6512 15988 6518 16040
rect 6564 16037 6592 16068
rect 6730 16056 6736 16068
rect 6788 16056 6794 16108
rect 6549 16031 6607 16037
rect 6549 15997 6561 16031
rect 6595 15997 6607 16031
rect 6549 15991 6607 15997
rect 6641 16031 6699 16037
rect 6641 15997 6653 16031
rect 6687 15997 6699 16031
rect 7006 16028 7012 16040
rect 6967 16000 7012 16028
rect 6641 15991 6699 15997
rect 4430 15960 4436 15972
rect 3896 15932 4436 15960
rect 4430 15920 4436 15932
rect 4488 15920 4494 15972
rect 4798 15920 4804 15972
rect 4856 15920 4862 15972
rect 6089 15963 6147 15969
rect 6089 15929 6101 15963
rect 6135 15960 6147 15963
rect 6656 15960 6684 15991
rect 7006 15988 7012 16000
rect 7064 15988 7070 16040
rect 7193 16031 7251 16037
rect 7193 15997 7205 16031
rect 7239 15997 7251 16031
rect 7193 15991 7251 15997
rect 6135 15932 6684 15960
rect 7208 15960 7236 15991
rect 7282 15988 7288 16040
rect 7340 16028 7346 16040
rect 9508 16037 9536 16136
rect 10410 16124 10416 16136
rect 10468 16124 10474 16176
rect 10229 16099 10287 16105
rect 10229 16096 10241 16099
rect 9692 16068 10241 16096
rect 9692 16037 9720 16068
rect 10229 16065 10241 16068
rect 10275 16096 10287 16099
rect 10597 16099 10655 16105
rect 10597 16096 10609 16099
rect 10275 16068 10609 16096
rect 10275 16065 10287 16068
rect 10229 16059 10287 16065
rect 10597 16065 10609 16068
rect 10643 16065 10655 16099
rect 10597 16059 10655 16065
rect 10686 16056 10692 16108
rect 10744 16096 10750 16108
rect 10873 16099 10931 16105
rect 10873 16096 10885 16099
rect 10744 16068 10885 16096
rect 10744 16056 10750 16068
rect 10873 16065 10885 16068
rect 10919 16065 10931 16099
rect 13446 16096 13452 16108
rect 10873 16059 10931 16065
rect 12452 16068 13452 16096
rect 12452 16040 12480 16068
rect 13446 16056 13452 16068
rect 13504 16096 13510 16108
rect 15013 16099 15071 16105
rect 15013 16096 15025 16099
rect 13504 16068 15025 16096
rect 13504 16056 13510 16068
rect 15013 16065 15025 16068
rect 15059 16065 15071 16099
rect 15013 16059 15071 16065
rect 15289 16099 15347 16105
rect 15289 16065 15301 16099
rect 15335 16096 15347 16099
rect 16022 16096 16028 16108
rect 15335 16068 16028 16096
rect 15335 16065 15347 16068
rect 15289 16059 15347 16065
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 9493 16031 9551 16037
rect 7340 16000 7385 16028
rect 7340 15988 7346 16000
rect 9493 15997 9505 16031
rect 9539 15997 9551 16031
rect 9493 15991 9551 15997
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 15997 9735 16031
rect 9950 16028 9956 16040
rect 9911 16000 9956 16028
rect 9677 15991 9735 15997
rect 9950 15988 9956 16000
rect 10008 15988 10014 16040
rect 10134 16028 10140 16040
rect 10095 16000 10140 16028
rect 10134 15988 10140 16000
rect 10192 15988 10198 16040
rect 10321 16031 10379 16037
rect 10321 15997 10333 16031
rect 10367 16028 10379 16031
rect 10410 16028 10416 16040
rect 10367 16000 10416 16028
rect 10367 15997 10379 16000
rect 10321 15991 10379 15997
rect 10410 15988 10416 16000
rect 10468 15988 10474 16040
rect 10505 16031 10563 16037
rect 10505 15997 10517 16031
rect 10551 15997 10563 16031
rect 10505 15991 10563 15997
rect 10781 16031 10839 16037
rect 10781 15997 10793 16031
rect 10827 15997 10839 16031
rect 12434 16028 12440 16040
rect 12395 16000 12440 16028
rect 10781 15991 10839 15997
rect 8386 15960 8392 15972
rect 7208 15932 8392 15960
rect 6135 15929 6147 15932
rect 6089 15923 6147 15929
rect 1581 15895 1639 15901
rect 1581 15861 1593 15895
rect 1627 15892 1639 15895
rect 4890 15892 4896 15904
rect 1627 15864 4896 15892
rect 1627 15861 1639 15864
rect 1581 15855 1639 15861
rect 4890 15852 4896 15864
rect 4948 15852 4954 15904
rect 5629 15895 5687 15901
rect 5629 15861 5641 15895
rect 5675 15892 5687 15895
rect 6104 15892 6132 15923
rect 8386 15920 8392 15932
rect 8444 15920 8450 15972
rect 5675 15864 6132 15892
rect 5675 15861 5687 15864
rect 5629 15855 5687 15861
rect 8846 15852 8852 15904
rect 8904 15892 8910 15904
rect 9493 15895 9551 15901
rect 9493 15892 9505 15895
rect 8904 15864 9505 15892
rect 8904 15852 8910 15864
rect 9493 15861 9505 15864
rect 9539 15861 9551 15895
rect 9766 15892 9772 15904
rect 9727 15864 9772 15892
rect 9493 15855 9551 15861
rect 9766 15852 9772 15864
rect 9824 15852 9830 15904
rect 10042 15852 10048 15904
rect 10100 15892 10106 15904
rect 10520 15892 10548 15991
rect 10594 15920 10600 15972
rect 10652 15960 10658 15972
rect 10796 15960 10824 15991
rect 12434 15988 12440 16000
rect 12492 15988 12498 16040
rect 10652 15932 10824 15960
rect 12713 15963 12771 15969
rect 10652 15920 10658 15932
rect 12713 15929 12725 15963
rect 12759 15929 12771 15963
rect 12713 15923 12771 15929
rect 11241 15895 11299 15901
rect 11241 15892 11253 15895
rect 10100 15864 11253 15892
rect 10100 15852 10106 15864
rect 11241 15861 11253 15864
rect 11287 15861 11299 15895
rect 12728 15892 12756 15923
rect 13446 15920 13452 15972
rect 13504 15920 13510 15972
rect 16022 15920 16028 15972
rect 16080 15920 16086 15972
rect 12894 15892 12900 15904
rect 12728 15864 12900 15892
rect 11241 15855 11299 15861
rect 12894 15852 12900 15864
rect 12952 15852 12958 15904
rect 12986 15852 12992 15904
rect 13044 15892 13050 15904
rect 14185 15895 14243 15901
rect 14185 15892 14197 15895
rect 13044 15864 14197 15892
rect 13044 15852 13050 15864
rect 14185 15861 14197 15864
rect 14231 15861 14243 15895
rect 14185 15855 14243 15861
rect 1104 15802 17296 15824
rect 1104 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 6571 15802
rect 6623 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 11904 15802
rect 11956 15750 11968 15802
rect 12020 15750 17296 15802
rect 1104 15728 17296 15750
rect 3510 15648 3516 15700
rect 3568 15688 3574 15700
rect 3881 15691 3939 15697
rect 3881 15688 3893 15691
rect 3568 15660 3893 15688
rect 3568 15648 3574 15660
rect 3881 15657 3893 15660
rect 3927 15657 3939 15691
rect 10042 15688 10048 15700
rect 10003 15660 10048 15688
rect 3881 15651 3939 15657
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 12986 15688 12992 15700
rect 12544 15660 12992 15688
rect 2958 15580 2964 15632
rect 3016 15620 3022 15632
rect 3053 15623 3111 15629
rect 3053 15620 3065 15623
rect 3016 15592 3065 15620
rect 3016 15580 3022 15592
rect 3053 15589 3065 15592
rect 3099 15620 3111 15623
rect 8205 15623 8263 15629
rect 8205 15620 8217 15623
rect 3099 15592 4108 15620
rect 3099 15589 3111 15592
rect 3053 15583 3111 15589
rect 2130 15552 2136 15564
rect 2091 15524 2136 15552
rect 2130 15512 2136 15524
rect 2188 15512 2194 15564
rect 3142 15512 3148 15564
rect 3200 15552 3206 15564
rect 3237 15555 3295 15561
rect 3237 15552 3249 15555
rect 3200 15524 3249 15552
rect 3200 15512 3206 15524
rect 3237 15521 3249 15524
rect 3283 15521 3295 15555
rect 3237 15515 3295 15521
rect 3326 15512 3332 15564
rect 3384 15552 3390 15564
rect 4080 15561 4108 15592
rect 4816 15592 8217 15620
rect 3605 15555 3663 15561
rect 3384 15524 3429 15552
rect 3384 15512 3390 15524
rect 3605 15521 3617 15555
rect 3651 15521 3663 15555
rect 3605 15515 3663 15521
rect 3697 15555 3755 15561
rect 3697 15521 3709 15555
rect 3743 15552 3755 15555
rect 3881 15555 3939 15561
rect 3881 15552 3893 15555
rect 3743 15524 3893 15552
rect 3743 15521 3755 15524
rect 3697 15515 3755 15521
rect 3881 15521 3893 15524
rect 3927 15521 3939 15555
rect 3881 15515 3939 15521
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15521 4123 15555
rect 4065 15515 4123 15521
rect 3620 15484 3648 15515
rect 4706 15512 4712 15564
rect 4764 15552 4770 15564
rect 4816 15561 4844 15592
rect 8205 15589 8217 15592
rect 8251 15589 8263 15623
rect 8846 15620 8852 15632
rect 8807 15592 8852 15620
rect 8205 15583 8263 15589
rect 8846 15580 8852 15592
rect 8904 15580 8910 15632
rect 10229 15623 10287 15629
rect 10229 15589 10241 15623
rect 10275 15620 10287 15623
rect 10686 15620 10692 15632
rect 10275 15592 10692 15620
rect 10275 15589 10287 15592
rect 10229 15583 10287 15589
rect 10686 15580 10692 15592
rect 10744 15580 10750 15632
rect 12268 15592 12434 15620
rect 12268 15564 12296 15592
rect 4801 15555 4859 15561
rect 4801 15552 4813 15555
rect 4764 15524 4813 15552
rect 4764 15512 4770 15524
rect 4801 15521 4813 15524
rect 4847 15521 4859 15555
rect 7190 15552 7196 15564
rect 7151 15524 7196 15552
rect 4801 15515 4859 15521
rect 7190 15512 7196 15524
rect 7248 15512 7254 15564
rect 7558 15552 7564 15564
rect 7519 15524 7564 15552
rect 7558 15512 7564 15524
rect 7616 15512 7622 15564
rect 8386 15552 8392 15564
rect 8347 15524 8392 15552
rect 8386 15512 8392 15524
rect 8444 15512 8450 15564
rect 8481 15555 8539 15561
rect 8481 15521 8493 15555
rect 8527 15552 8539 15555
rect 9309 15555 9367 15561
rect 9309 15552 9321 15555
rect 8527 15524 9321 15552
rect 8527 15521 8539 15524
rect 8481 15515 8539 15521
rect 9309 15521 9321 15524
rect 9355 15552 9367 15555
rect 9766 15552 9772 15564
rect 9355 15524 9772 15552
rect 9355 15521 9367 15524
rect 9309 15515 9367 15521
rect 9766 15512 9772 15524
rect 9824 15512 9830 15564
rect 10413 15555 10471 15561
rect 10413 15521 10425 15555
rect 10459 15552 10471 15555
rect 10594 15552 10600 15564
rect 10459 15524 10600 15552
rect 10459 15521 10471 15524
rect 10413 15515 10471 15521
rect 10594 15512 10600 15524
rect 10652 15512 10658 15564
rect 11974 15552 11980 15564
rect 11935 15524 11980 15552
rect 11974 15512 11980 15524
rect 12032 15512 12038 15564
rect 12161 15555 12219 15561
rect 12161 15521 12173 15555
rect 12207 15521 12219 15555
rect 12161 15515 12219 15521
rect 4338 15484 4344 15496
rect 3620 15456 4344 15484
rect 4338 15444 4344 15456
rect 4396 15444 4402 15496
rect 7282 15484 7288 15496
rect 7243 15456 7288 15484
rect 7282 15444 7288 15456
rect 7340 15444 7346 15496
rect 7745 15487 7803 15493
rect 7745 15453 7757 15487
rect 7791 15484 7803 15487
rect 7834 15484 7840 15496
rect 7791 15456 7840 15484
rect 7791 15453 7803 15456
rect 7745 15447 7803 15453
rect 7834 15444 7840 15456
rect 7892 15444 7898 15496
rect 8021 15487 8079 15493
rect 8021 15453 8033 15487
rect 8067 15484 8079 15487
rect 8110 15484 8116 15496
rect 8067 15456 8116 15484
rect 8067 15453 8079 15456
rect 8021 15447 8079 15453
rect 8110 15444 8116 15456
rect 8168 15444 8174 15496
rect 8665 15487 8723 15493
rect 8665 15453 8677 15487
rect 8711 15453 8723 15487
rect 8665 15447 8723 15453
rect 8757 15487 8815 15493
rect 8757 15453 8769 15487
rect 8803 15484 8815 15487
rect 12066 15484 12072 15496
rect 8803 15456 12072 15484
rect 8803 15453 8815 15456
rect 8757 15447 8815 15453
rect 3418 15376 3424 15428
rect 3476 15416 3482 15428
rect 3697 15419 3755 15425
rect 3697 15416 3709 15419
rect 3476 15388 3709 15416
rect 3476 15376 3482 15388
rect 3697 15385 3709 15388
rect 3743 15385 3755 15419
rect 3697 15379 3755 15385
rect 4062 15376 4068 15428
rect 4120 15416 4126 15428
rect 4893 15419 4951 15425
rect 4893 15416 4905 15419
rect 4120 15388 4905 15416
rect 4120 15376 4126 15388
rect 4893 15385 4905 15388
rect 4939 15385 4951 15419
rect 4893 15379 4951 15385
rect 7929 15419 7987 15425
rect 7929 15385 7941 15419
rect 7975 15416 7987 15419
rect 8680 15416 8708 15447
rect 12066 15444 12072 15456
rect 12124 15444 12130 15496
rect 9490 15416 9496 15428
rect 7975 15388 9496 15416
rect 7975 15385 7987 15388
rect 7929 15379 7987 15385
rect 9490 15376 9496 15388
rect 9548 15376 9554 15428
rect 12176 15416 12204 15515
rect 12250 15512 12256 15564
rect 12308 15552 12314 15564
rect 12406 15552 12434 15592
rect 12544 15561 12572 15660
rect 12986 15648 12992 15660
rect 13044 15648 13050 15700
rect 13446 15648 13452 15700
rect 13504 15688 13510 15700
rect 13541 15691 13599 15697
rect 13541 15688 13553 15691
rect 13504 15660 13553 15688
rect 13504 15648 13510 15660
rect 13541 15657 13553 15660
rect 13587 15657 13599 15691
rect 13541 15651 13599 15657
rect 16022 15648 16028 15700
rect 16080 15688 16086 15700
rect 16117 15691 16175 15697
rect 16117 15688 16129 15691
rect 16080 15660 16129 15688
rect 16080 15648 16086 15660
rect 16117 15657 16129 15660
rect 16163 15657 16175 15691
rect 16117 15651 16175 15657
rect 12529 15555 12587 15561
rect 12308 15524 12353 15552
rect 12406 15524 12480 15552
rect 12308 15512 12314 15524
rect 12342 15484 12348 15496
rect 12303 15456 12348 15484
rect 12342 15444 12348 15456
rect 12400 15444 12406 15496
rect 12452 15484 12480 15524
rect 12529 15521 12541 15555
rect 12575 15521 12587 15555
rect 12529 15515 12587 15521
rect 12802 15512 12808 15564
rect 12860 15552 12866 15564
rect 12986 15552 12992 15564
rect 12860 15524 12905 15552
rect 12947 15524 12992 15552
rect 12860 15512 12866 15524
rect 12986 15512 12992 15524
rect 13044 15512 13050 15564
rect 13354 15552 13360 15564
rect 13315 15524 13360 15552
rect 13354 15512 13360 15524
rect 13412 15512 13418 15564
rect 14553 15555 14611 15561
rect 14553 15521 14565 15555
rect 14599 15552 14611 15555
rect 15286 15552 15292 15564
rect 14599 15524 15292 15552
rect 14599 15521 14611 15524
rect 14553 15515 14611 15521
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 15746 15512 15752 15564
rect 15804 15552 15810 15564
rect 16301 15555 16359 15561
rect 16301 15552 16313 15555
rect 15804 15524 16313 15552
rect 15804 15512 15810 15524
rect 16301 15521 16313 15524
rect 16347 15552 16359 15555
rect 16482 15552 16488 15564
rect 16347 15524 16488 15552
rect 16347 15521 16359 15524
rect 16301 15515 16359 15521
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 12897 15487 12955 15493
rect 12897 15484 12909 15487
rect 12452 15456 12909 15484
rect 12897 15453 12909 15456
rect 12943 15453 12955 15487
rect 12897 15447 12955 15453
rect 12618 15416 12624 15428
rect 12176 15388 12624 15416
rect 12618 15376 12624 15388
rect 12676 15376 12682 15428
rect 1854 15308 1860 15360
rect 1912 15348 1918 15360
rect 1949 15351 2007 15357
rect 1949 15348 1961 15351
rect 1912 15320 1961 15348
rect 1912 15308 1918 15320
rect 1949 15317 1961 15320
rect 1995 15317 2007 15351
rect 1949 15311 2007 15317
rect 3513 15351 3571 15357
rect 3513 15317 3525 15351
rect 3559 15348 3571 15351
rect 4154 15348 4160 15360
rect 3559 15320 4160 15348
rect 3559 15317 3571 15320
rect 3513 15311 3571 15317
rect 4154 15308 4160 15320
rect 4212 15308 4218 15360
rect 8478 15308 8484 15360
rect 8536 15348 8542 15360
rect 9217 15351 9275 15357
rect 9217 15348 9229 15351
rect 8536 15320 9229 15348
rect 8536 15308 8542 15320
rect 9217 15317 9229 15320
rect 9263 15317 9275 15351
rect 9217 15311 9275 15317
rect 12713 15351 12771 15357
rect 12713 15317 12725 15351
rect 12759 15348 12771 15351
rect 12894 15348 12900 15360
rect 12759 15320 12900 15348
rect 12759 15317 12771 15320
rect 12713 15311 12771 15317
rect 12894 15308 12900 15320
rect 12952 15308 12958 15360
rect 13814 15308 13820 15360
rect 13872 15348 13878 15360
rect 14461 15351 14519 15357
rect 14461 15348 14473 15351
rect 13872 15320 14473 15348
rect 13872 15308 13878 15320
rect 14461 15317 14473 15320
rect 14507 15317 14519 15351
rect 14461 15311 14519 15317
rect 1104 15258 17296 15280
rect 1104 15206 3680 15258
rect 3732 15206 3744 15258
rect 3796 15206 3808 15258
rect 3860 15206 3872 15258
rect 3924 15206 9078 15258
rect 9130 15206 9142 15258
rect 9194 15206 9206 15258
rect 9258 15206 9270 15258
rect 9322 15206 14475 15258
rect 14527 15206 14539 15258
rect 14591 15206 14603 15258
rect 14655 15206 14667 15258
rect 14719 15206 17296 15258
rect 1104 15184 17296 15206
rect 1397 15147 1455 15153
rect 1397 15113 1409 15147
rect 1443 15144 1455 15147
rect 3142 15144 3148 15156
rect 1443 15116 3148 15144
rect 1443 15113 1455 15116
rect 1397 15107 1455 15113
rect 3142 15104 3148 15116
rect 3200 15104 3206 15156
rect 4430 15144 4436 15156
rect 3252 15116 4436 15144
rect 3145 14943 3203 14949
rect 3145 14909 3157 14943
rect 3191 14940 3203 14943
rect 3252 14940 3280 15116
rect 4430 15104 4436 15116
rect 4488 15104 4494 15156
rect 7282 15104 7288 15156
rect 7340 15144 7346 15156
rect 7469 15147 7527 15153
rect 7469 15144 7481 15147
rect 7340 15116 7481 15144
rect 7340 15104 7346 15116
rect 7469 15113 7481 15116
rect 7515 15113 7527 15147
rect 10962 15144 10968 15156
rect 7469 15107 7527 15113
rect 7576 15116 10968 15144
rect 3326 15036 3332 15088
rect 3384 15076 3390 15088
rect 4246 15076 4252 15088
rect 3384 15048 4252 15076
rect 3384 15036 3390 15048
rect 4246 15036 4252 15048
rect 4304 15036 4310 15088
rect 6822 15076 6828 15088
rect 6735 15048 6828 15076
rect 6822 15036 6828 15048
rect 6880 15076 6886 15088
rect 7576 15076 7604 15116
rect 10962 15104 10968 15116
rect 11020 15104 11026 15156
rect 12342 15104 12348 15156
rect 12400 15144 12406 15156
rect 12802 15144 12808 15156
rect 12400 15116 12808 15144
rect 12400 15104 12406 15116
rect 12802 15104 12808 15116
rect 12860 15104 12866 15156
rect 14366 15104 14372 15156
rect 14424 15144 14430 15156
rect 15010 15144 15016 15156
rect 14424 15116 15016 15144
rect 14424 15104 14430 15116
rect 15010 15104 15016 15116
rect 15068 15104 15074 15156
rect 15286 15104 15292 15156
rect 15344 15144 15350 15156
rect 15473 15147 15531 15153
rect 15473 15144 15485 15147
rect 15344 15116 15485 15144
rect 15344 15104 15350 15116
rect 15473 15113 15485 15116
rect 15519 15113 15531 15147
rect 15473 15107 15531 15113
rect 6880 15048 7604 15076
rect 7837 15079 7895 15085
rect 6880 15036 6886 15048
rect 7837 15045 7849 15079
rect 7883 15045 7895 15079
rect 7837 15039 7895 15045
rect 9677 15079 9735 15085
rect 9677 15045 9689 15079
rect 9723 15076 9735 15079
rect 9723 15048 14044 15076
rect 9723 15045 9735 15048
rect 9677 15039 9735 15045
rect 4065 15011 4123 15017
rect 3738 14980 4016 15008
rect 3738 14952 3766 14980
rect 3191 14912 3280 14940
rect 3191 14909 3203 14912
rect 3145 14903 3203 14909
rect 3326 14900 3332 14952
rect 3384 14940 3390 14952
rect 3421 14943 3479 14949
rect 3421 14940 3433 14943
rect 3384 14912 3433 14940
rect 3384 14900 3390 14912
rect 3421 14909 3433 14912
rect 3467 14909 3479 14943
rect 3421 14903 3479 14909
rect 3694 14900 3700 14952
rect 3752 14949 3766 14952
rect 3752 14943 3781 14949
rect 3769 14909 3781 14943
rect 3878 14940 3884 14952
rect 3839 14912 3884 14940
rect 3752 14903 3781 14909
rect 3752 14900 3758 14903
rect 3878 14900 3884 14912
rect 3936 14900 3942 14952
rect 3988 14949 4016 14980
rect 4065 14977 4077 15011
rect 4111 15008 4123 15011
rect 4338 15008 4344 15020
rect 4111 14980 4344 15008
rect 4111 14977 4123 14980
rect 4065 14971 4123 14977
rect 3973 14943 4031 14949
rect 3973 14909 3985 14943
rect 4019 14909 4031 14943
rect 3973 14903 4031 14909
rect 1854 14832 1860 14884
rect 1912 14832 1918 14884
rect 2869 14875 2927 14881
rect 2869 14841 2881 14875
rect 2915 14872 2927 14875
rect 3237 14875 3295 14881
rect 3237 14872 3249 14875
rect 2915 14844 3249 14872
rect 2915 14841 2927 14844
rect 2869 14835 2927 14841
rect 3237 14841 3249 14844
rect 3283 14841 3295 14875
rect 3510 14872 3516 14884
rect 3471 14844 3516 14872
rect 3237 14835 3295 14841
rect 3510 14832 3516 14844
rect 3568 14832 3574 14884
rect 3605 14875 3663 14881
rect 3605 14841 3617 14875
rect 3651 14872 3663 14875
rect 4062 14872 4068 14884
rect 3651 14844 4068 14872
rect 3651 14841 3663 14844
rect 3605 14835 3663 14841
rect 2774 14764 2780 14816
rect 2832 14804 2838 14816
rect 3620 14804 3648 14835
rect 4062 14832 4068 14844
rect 4120 14832 4126 14884
rect 2832 14776 3648 14804
rect 2832 14764 2838 14776
rect 3694 14764 3700 14816
rect 3752 14804 3758 14816
rect 4172 14804 4200 14980
rect 4338 14968 4344 14980
rect 4396 14968 4402 15020
rect 5442 14940 5448 14952
rect 5403 14912 5448 14940
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 6840 14949 6868 15036
rect 7190 14968 7196 15020
rect 7248 15008 7254 15020
rect 7285 15011 7343 15017
rect 7285 15008 7297 15011
rect 7248 14980 7297 15008
rect 7248 14968 7254 14980
rect 7285 14977 7297 14980
rect 7331 15008 7343 15011
rect 7561 15011 7619 15017
rect 7561 15008 7573 15011
rect 7331 14980 7573 15008
rect 7331 14977 7343 14980
rect 7285 14971 7343 14977
rect 7561 14977 7573 14980
rect 7607 14977 7619 15011
rect 7852 15008 7880 15039
rect 9490 15008 9496 15020
rect 7852 14980 8984 15008
rect 9451 14980 9496 15008
rect 7561 14971 7619 14977
rect 6825 14943 6883 14949
rect 6825 14909 6837 14943
rect 6871 14909 6883 14943
rect 6825 14903 6883 14909
rect 7377 14943 7435 14949
rect 7377 14909 7389 14943
rect 7423 14909 7435 14943
rect 7377 14903 7435 14909
rect 7469 14943 7527 14949
rect 7469 14909 7481 14943
rect 7515 14940 7527 14943
rect 8110 14940 8116 14952
rect 7515 14912 8116 14940
rect 7515 14909 7527 14912
rect 7469 14903 7527 14909
rect 7006 14872 7012 14884
rect 6967 14844 7012 14872
rect 7006 14832 7012 14844
rect 7064 14832 7070 14884
rect 7392 14872 7420 14903
rect 8110 14900 8116 14912
rect 8168 14900 8174 14952
rect 8478 14940 8484 14952
rect 8439 14912 8484 14940
rect 8478 14900 8484 14912
rect 8536 14900 8542 14952
rect 8662 14940 8668 14952
rect 8623 14912 8668 14940
rect 8662 14900 8668 14912
rect 8720 14900 8726 14952
rect 8846 14940 8852 14952
rect 8807 14912 8852 14940
rect 8846 14900 8852 14912
rect 8904 14900 8910 14952
rect 8956 14949 8984 14980
rect 9490 14968 9496 14980
rect 9548 14968 9554 15020
rect 13814 15008 13820 15020
rect 9784 14980 13820 15008
rect 9784 14949 9812 14980
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 14016 15017 14044 15048
rect 14918 15036 14924 15088
rect 14976 15076 14982 15088
rect 14976 15048 15424 15076
rect 14976 15036 14982 15048
rect 14001 15011 14059 15017
rect 14001 14977 14013 15011
rect 14047 15008 14059 15011
rect 14553 15011 14611 15017
rect 14553 15008 14565 15011
rect 14047 14980 14565 15008
rect 14047 14977 14059 14980
rect 14001 14971 14059 14977
rect 14553 14977 14565 14980
rect 14599 14977 14611 15011
rect 15010 15008 15016 15020
rect 14971 14980 15016 15008
rect 14553 14971 14611 14977
rect 15010 14968 15016 14980
rect 15068 14968 15074 15020
rect 8941 14943 8999 14949
rect 8941 14909 8953 14943
rect 8987 14909 8999 14943
rect 8941 14903 8999 14909
rect 9309 14943 9367 14949
rect 9309 14909 9321 14943
rect 9355 14909 9367 14943
rect 9309 14903 9367 14909
rect 9769 14943 9827 14949
rect 9769 14909 9781 14943
rect 9815 14909 9827 14943
rect 9769 14903 9827 14909
rect 7558 14872 7564 14884
rect 7392 14844 7564 14872
rect 7558 14832 7564 14844
rect 7616 14832 7622 14884
rect 7929 14875 7987 14881
rect 7929 14841 7941 14875
rect 7975 14841 7987 14875
rect 9324 14872 9352 14903
rect 10502 14900 10508 14952
rect 10560 14940 10566 14952
rect 10597 14943 10655 14949
rect 10597 14940 10609 14943
rect 10560 14912 10609 14940
rect 10560 14900 10566 14912
rect 10597 14909 10609 14912
rect 10643 14940 10655 14943
rect 10686 14940 10692 14952
rect 10643 14912 10692 14940
rect 10643 14909 10655 14912
rect 10597 14903 10655 14909
rect 10686 14900 10692 14912
rect 10744 14900 10750 14952
rect 10870 14940 10876 14952
rect 10831 14912 10876 14940
rect 10870 14900 10876 14912
rect 10928 14900 10934 14952
rect 10962 14900 10968 14952
rect 11020 14940 11026 14952
rect 12250 14940 12256 14952
rect 11020 14912 12256 14940
rect 11020 14900 11026 14912
rect 12250 14900 12256 14912
rect 12308 14900 12314 14952
rect 14185 14943 14243 14949
rect 14185 14909 14197 14943
rect 14231 14909 14243 14943
rect 14185 14903 14243 14909
rect 9493 14875 9551 14881
rect 9493 14872 9505 14875
rect 9324 14844 9505 14872
rect 7929 14835 7987 14841
rect 9493 14841 9505 14844
rect 9539 14841 9551 14875
rect 9493 14835 9551 14841
rect 10781 14875 10839 14881
rect 10781 14841 10793 14875
rect 10827 14841 10839 14875
rect 10781 14835 10839 14841
rect 3752 14776 4200 14804
rect 3752 14764 3758 14776
rect 5534 14764 5540 14816
rect 5592 14804 5598 14816
rect 5629 14807 5687 14813
rect 5629 14804 5641 14807
rect 5592 14776 5641 14804
rect 5592 14764 5598 14776
rect 5629 14773 5641 14776
rect 5675 14773 5687 14807
rect 5629 14767 5687 14773
rect 6822 14764 6828 14816
rect 6880 14804 6886 14816
rect 7944 14804 7972 14835
rect 6880 14776 7972 14804
rect 6880 14764 6886 14776
rect 10502 14764 10508 14816
rect 10560 14804 10566 14816
rect 10796 14804 10824 14835
rect 12066 14832 12072 14884
rect 12124 14872 12130 14884
rect 14200 14872 14228 14903
rect 14366 14900 14372 14952
rect 14424 14940 14430 14952
rect 14461 14943 14519 14949
rect 14461 14940 14473 14943
rect 14424 14912 14473 14940
rect 14424 14900 14430 14912
rect 14461 14909 14473 14912
rect 14507 14909 14519 14943
rect 14754 14943 14812 14949
rect 14754 14940 14766 14943
rect 14461 14903 14519 14909
rect 14752 14909 14766 14940
rect 14800 14909 14812 14943
rect 14752 14903 14812 14909
rect 12124 14844 14228 14872
rect 14752 14872 14780 14903
rect 14918 14900 14924 14952
rect 14976 14940 14982 14952
rect 15102 14940 15108 14952
rect 14976 14912 15021 14940
rect 15063 14912 15108 14940
rect 14976 14900 14982 14912
rect 15102 14900 15108 14912
rect 15160 14900 15166 14952
rect 15286 14940 15292 14952
rect 15247 14912 15292 14940
rect 15286 14900 15292 14912
rect 15344 14900 15350 14952
rect 15396 14949 15424 15048
rect 15381 14943 15439 14949
rect 15381 14909 15393 14943
rect 15427 14909 15439 14943
rect 15562 14940 15568 14952
rect 15523 14912 15568 14940
rect 15381 14903 15439 14909
rect 15562 14900 15568 14912
rect 15620 14900 15626 14952
rect 16758 14940 16764 14952
rect 16719 14912 16764 14940
rect 16758 14900 16764 14912
rect 16816 14900 16822 14952
rect 15580 14872 15608 14900
rect 14752 14844 15608 14872
rect 12124 14832 12130 14844
rect 10962 14804 10968 14816
rect 10560 14776 10968 14804
rect 10560 14764 10566 14776
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 11149 14807 11207 14813
rect 11149 14773 11161 14807
rect 11195 14804 11207 14807
rect 12158 14804 12164 14816
rect 11195 14776 12164 14804
rect 11195 14773 11207 14776
rect 11149 14767 11207 14773
rect 12158 14764 12164 14776
rect 12216 14764 12222 14816
rect 14369 14807 14427 14813
rect 14369 14773 14381 14807
rect 14415 14804 14427 14807
rect 15102 14804 15108 14816
rect 14415 14776 15108 14804
rect 14415 14773 14427 14776
rect 14369 14767 14427 14773
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 16577 14807 16635 14813
rect 16577 14773 16589 14807
rect 16623 14804 16635 14807
rect 16666 14804 16672 14816
rect 16623 14776 16672 14804
rect 16623 14773 16635 14776
rect 16577 14767 16635 14773
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 1104 14714 17296 14736
rect 1104 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 6571 14714
rect 6623 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 11904 14714
rect 11956 14662 11968 14714
rect 12020 14662 17296 14714
rect 1104 14640 17296 14662
rect 3326 14600 3332 14612
rect 3287 14572 3332 14600
rect 3326 14560 3332 14572
rect 3384 14560 3390 14612
rect 4065 14603 4123 14609
rect 4065 14569 4077 14603
rect 4111 14600 4123 14603
rect 4246 14600 4252 14612
rect 4111 14572 4252 14600
rect 4111 14569 4123 14572
rect 4065 14563 4123 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 4632 14572 6132 14600
rect 2958 14532 2964 14544
rect 2919 14504 2964 14532
rect 2958 14492 2964 14504
rect 3016 14492 3022 14544
rect 3145 14535 3203 14541
rect 3145 14501 3157 14535
rect 3191 14532 3203 14535
rect 3418 14532 3424 14544
rect 3191 14504 3424 14532
rect 3191 14501 3203 14504
rect 3145 14495 3203 14501
rect 3418 14492 3424 14504
rect 3476 14492 3482 14544
rect 4430 14532 4436 14544
rect 3528 14504 4436 14532
rect 1394 14464 1400 14476
rect 1355 14436 1400 14464
rect 1394 14424 1400 14436
rect 1452 14424 1458 14476
rect 3326 14424 3332 14476
rect 3384 14464 3390 14476
rect 3528 14464 3556 14504
rect 4430 14492 4436 14504
rect 4488 14532 4494 14544
rect 4632 14532 4660 14572
rect 4488 14504 4660 14532
rect 4488 14492 4494 14504
rect 3694 14464 3700 14476
rect 3384 14436 3556 14464
rect 3655 14436 3700 14464
rect 3384 14424 3390 14436
rect 3694 14424 3700 14436
rect 3752 14424 3758 14476
rect 3973 14467 4031 14473
rect 3973 14433 3985 14467
rect 4019 14464 4031 14467
rect 4154 14464 4160 14476
rect 4019 14436 4160 14464
rect 4019 14433 4031 14436
rect 3973 14427 4031 14433
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14396 3479 14399
rect 3510 14396 3516 14408
rect 3467 14368 3516 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 3510 14356 3516 14368
rect 3568 14356 3574 14408
rect 3605 14399 3663 14405
rect 3605 14365 3617 14399
rect 3651 14396 3663 14399
rect 3988 14396 4016 14427
rect 4154 14424 4160 14436
rect 4212 14464 4218 14476
rect 4338 14464 4344 14476
rect 4212 14436 4344 14464
rect 4212 14424 4218 14436
rect 4338 14424 4344 14436
rect 4396 14424 4402 14476
rect 4540 14473 4568 14504
rect 5534 14492 5540 14544
rect 5592 14492 5598 14544
rect 4525 14467 4583 14473
rect 4525 14433 4537 14467
rect 4571 14433 4583 14467
rect 4525 14427 4583 14433
rect 3651 14368 4016 14396
rect 4801 14399 4859 14405
rect 3651 14365 3663 14368
rect 3605 14359 3663 14365
rect 4801 14365 4813 14399
rect 4847 14396 4859 14399
rect 5258 14396 5264 14408
rect 4847 14368 5264 14396
rect 4847 14365 4859 14368
rect 4801 14359 4859 14365
rect 5258 14356 5264 14368
rect 5316 14356 5322 14408
rect 6104 14396 6132 14572
rect 7282 14560 7288 14612
rect 7340 14600 7346 14612
rect 7745 14603 7803 14609
rect 7745 14600 7757 14603
rect 7340 14572 7757 14600
rect 7340 14560 7346 14572
rect 7745 14569 7757 14572
rect 7791 14569 7803 14603
rect 7745 14563 7803 14569
rect 10413 14603 10471 14609
rect 10413 14569 10425 14603
rect 10459 14600 10471 14603
rect 10689 14603 10747 14609
rect 10689 14600 10701 14603
rect 10459 14572 10701 14600
rect 10459 14569 10471 14572
rect 10413 14563 10471 14569
rect 10689 14569 10701 14572
rect 10735 14600 10747 14603
rect 10778 14600 10784 14612
rect 10735 14572 10784 14600
rect 10735 14569 10747 14572
rect 10689 14563 10747 14569
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 12434 14600 12440 14612
rect 10888 14572 12440 14600
rect 7006 14492 7012 14544
rect 7064 14532 7070 14544
rect 10888 14532 10916 14572
rect 12434 14560 12440 14572
rect 12492 14600 12498 14612
rect 12492 14572 13216 14600
rect 12492 14560 12498 14572
rect 7064 14504 10916 14532
rect 7064 14492 7070 14504
rect 7834 14464 7840 14476
rect 7795 14436 7840 14464
rect 7834 14424 7840 14436
rect 7892 14424 7898 14476
rect 10502 14473 10508 14476
rect 10472 14467 10508 14473
rect 10472 14433 10484 14467
rect 10472 14427 10508 14433
rect 10502 14424 10508 14427
rect 10560 14424 10566 14476
rect 9953 14399 10011 14405
rect 6104 14368 8064 14396
rect 8036 14340 8064 14368
rect 9953 14365 9965 14399
rect 9999 14396 10011 14399
rect 10318 14396 10324 14408
rect 9999 14368 10324 14396
rect 9999 14365 10011 14368
rect 9953 14359 10011 14365
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 10686 14356 10692 14408
rect 10744 14396 10750 14408
rect 10888 14396 10916 14504
rect 11606 14492 11612 14544
rect 11664 14492 11670 14544
rect 12158 14532 12164 14544
rect 12119 14504 12164 14532
rect 12158 14492 12164 14504
rect 12216 14492 12222 14544
rect 12897 14535 12955 14541
rect 12897 14501 12909 14535
rect 12943 14532 12955 14535
rect 12986 14532 12992 14544
rect 12943 14504 12992 14532
rect 12943 14501 12955 14504
rect 12897 14495 12955 14501
rect 12986 14492 12992 14504
rect 13044 14492 13050 14544
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 12526 14464 12532 14476
rect 12483 14436 12532 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 12526 14424 12532 14436
rect 12584 14424 12590 14476
rect 12710 14464 12716 14476
rect 12671 14436 12716 14464
rect 12710 14424 12716 14436
rect 12768 14424 12774 14476
rect 12802 14424 12808 14476
rect 12860 14464 12866 14476
rect 13188 14473 13216 14572
rect 14090 14492 14096 14544
rect 14148 14532 14154 14544
rect 15105 14535 15163 14541
rect 15105 14532 15117 14535
rect 14148 14504 15117 14532
rect 14148 14492 14154 14504
rect 15105 14501 15117 14504
rect 15151 14501 15163 14535
rect 15105 14495 15163 14501
rect 15197 14535 15255 14541
rect 15197 14501 15209 14535
rect 15243 14532 15255 14535
rect 15562 14532 15568 14544
rect 15243 14504 15568 14532
rect 15243 14501 15255 14504
rect 15197 14495 15255 14501
rect 15562 14492 15568 14504
rect 15620 14492 15626 14544
rect 13081 14467 13139 14473
rect 12860 14436 12905 14464
rect 12860 14424 12866 14436
rect 13081 14433 13093 14467
rect 13127 14433 13139 14467
rect 13081 14427 13139 14433
rect 13173 14467 13231 14473
rect 13173 14433 13185 14467
rect 13219 14464 13231 14467
rect 14921 14467 14979 14473
rect 14921 14464 14933 14467
rect 13219 14436 14933 14464
rect 13219 14433 13231 14436
rect 13173 14427 13231 14433
rect 14921 14433 14933 14436
rect 14967 14433 14979 14467
rect 14921 14427 14979 14433
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14464 15347 14467
rect 15378 14464 15384 14476
rect 15335 14436 15384 14464
rect 15335 14433 15347 14436
rect 15289 14427 15347 14433
rect 10744 14368 10916 14396
rect 12544 14396 12572 14424
rect 13096 14396 13124 14427
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 14274 14396 14280 14408
rect 12544 14368 13032 14396
rect 13096 14368 14280 14396
rect 10744 14356 10750 14368
rect 8018 14288 8024 14340
rect 8076 14328 8082 14340
rect 9398 14328 9404 14340
rect 8076 14300 9404 14328
rect 8076 14288 8082 14300
rect 9398 14288 9404 14300
rect 9456 14328 9462 14340
rect 10410 14328 10416 14340
rect 9456 14300 10416 14328
rect 9456 14288 9462 14300
rect 10410 14288 10416 14300
rect 10468 14288 10474 14340
rect 10594 14328 10600 14340
rect 10555 14300 10600 14328
rect 10594 14288 10600 14300
rect 10652 14288 10658 14340
rect 13004 14328 13032 14368
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 13354 14328 13360 14340
rect 13004 14300 13360 14328
rect 13354 14288 13360 14300
rect 13412 14288 13418 14340
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14260 1639 14263
rect 1854 14260 1860 14272
rect 1627 14232 1860 14260
rect 1627 14229 1639 14232
rect 1581 14223 1639 14229
rect 1854 14220 1860 14232
rect 1912 14220 1918 14272
rect 3510 14260 3516 14272
rect 3471 14232 3516 14260
rect 3510 14220 3516 14232
rect 3568 14220 3574 14272
rect 5810 14220 5816 14272
rect 5868 14260 5874 14272
rect 6273 14263 6331 14269
rect 6273 14260 6285 14263
rect 5868 14232 6285 14260
rect 5868 14220 5874 14232
rect 6273 14229 6285 14232
rect 6319 14229 6331 14263
rect 10042 14260 10048 14272
rect 10003 14232 10048 14260
rect 6273 14223 6331 14229
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 12529 14263 12587 14269
rect 12529 14229 12541 14263
rect 12575 14260 12587 14263
rect 12618 14260 12624 14272
rect 12575 14232 12624 14260
rect 12575 14229 12587 14232
rect 12529 14223 12587 14229
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 15286 14220 15292 14272
rect 15344 14260 15350 14272
rect 15473 14263 15531 14269
rect 15473 14260 15485 14263
rect 15344 14232 15485 14260
rect 15344 14220 15350 14232
rect 15473 14229 15485 14232
rect 15519 14229 15531 14263
rect 15473 14223 15531 14229
rect 1104 14170 17296 14192
rect 1104 14118 3680 14170
rect 3732 14118 3744 14170
rect 3796 14118 3808 14170
rect 3860 14118 3872 14170
rect 3924 14118 9078 14170
rect 9130 14118 9142 14170
rect 9194 14118 9206 14170
rect 9258 14118 9270 14170
rect 9322 14118 14475 14170
rect 14527 14118 14539 14170
rect 14591 14118 14603 14170
rect 14655 14118 14667 14170
rect 14719 14118 17296 14170
rect 1104 14096 17296 14118
rect 5258 14056 5264 14068
rect 5219 14028 5264 14056
rect 5258 14016 5264 14028
rect 5316 14016 5322 14068
rect 8110 14056 8116 14068
rect 8071 14028 8116 14056
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 8846 14056 8852 14068
rect 8807 14028 8852 14056
rect 8846 14016 8852 14028
rect 8904 14016 8910 14068
rect 10410 14016 10416 14068
rect 10468 14056 10474 14068
rect 13354 14056 13360 14068
rect 10468 14028 13360 14056
rect 10468 14016 10474 14028
rect 2314 13948 2320 14000
rect 2372 13988 2378 14000
rect 2372 13960 6776 13988
rect 2372 13948 2378 13960
rect 6089 13923 6147 13929
rect 6089 13920 6101 13923
rect 5460 13892 6101 13920
rect 3510 13812 3516 13864
rect 3568 13852 3574 13864
rect 3973 13855 4031 13861
rect 3973 13852 3985 13855
rect 3568 13824 3985 13852
rect 3568 13812 3574 13824
rect 3973 13821 3985 13824
rect 4019 13821 4031 13855
rect 3973 13815 4031 13821
rect 4065 13855 4123 13861
rect 4065 13821 4077 13855
rect 4111 13852 4123 13855
rect 4706 13852 4712 13864
rect 4111 13824 4712 13852
rect 4111 13821 4123 13824
rect 4065 13815 4123 13821
rect 4706 13812 4712 13824
rect 4764 13812 4770 13864
rect 5460 13861 5488 13892
rect 6089 13889 6101 13892
rect 6135 13889 6147 13923
rect 6089 13883 6147 13889
rect 5445 13855 5503 13861
rect 5445 13821 5457 13855
rect 5491 13821 5503 13855
rect 5902 13852 5908 13864
rect 5863 13824 5908 13852
rect 5445 13815 5503 13821
rect 5902 13812 5908 13824
rect 5960 13812 5966 13864
rect 5994 13812 6000 13864
rect 6052 13852 6058 13864
rect 6181 13855 6239 13861
rect 6052 13824 6097 13852
rect 6052 13812 6058 13824
rect 6181 13821 6193 13855
rect 6227 13821 6239 13855
rect 6748 13852 6776 13960
rect 8297 13923 8355 13929
rect 8297 13889 8309 13923
rect 8343 13920 8355 13923
rect 8757 13923 8815 13929
rect 8343 13892 8708 13920
rect 8343 13889 8355 13892
rect 8297 13883 8355 13889
rect 8389 13855 8447 13861
rect 8389 13852 8401 13855
rect 6748 13824 8401 13852
rect 6181 13815 6239 13821
rect 8389 13821 8401 13824
rect 8435 13852 8447 13855
rect 8680 13852 8708 13892
rect 8757 13889 8769 13923
rect 8803 13920 8815 13923
rect 8864 13920 8892 14016
rect 9401 13991 9459 13997
rect 9401 13988 9413 13991
rect 8803 13892 8892 13920
rect 9232 13960 9413 13988
rect 8803 13889 8815 13892
rect 8757 13883 8815 13889
rect 9232 13861 9260 13960
rect 9401 13957 9413 13960
rect 9447 13957 9459 13991
rect 9401 13951 9459 13957
rect 10318 13948 10324 14000
rect 10376 13988 10382 14000
rect 10689 13991 10747 13997
rect 10689 13988 10701 13991
rect 10376 13960 10701 13988
rect 10376 13948 10382 13960
rect 10689 13957 10701 13960
rect 10735 13957 10747 13991
rect 10689 13951 10747 13957
rect 9950 13920 9956 13932
rect 9863 13892 9956 13920
rect 9950 13880 9956 13892
rect 10008 13920 10014 13932
rect 10137 13923 10195 13929
rect 10137 13920 10149 13923
rect 10008 13892 10149 13920
rect 10008 13880 10014 13892
rect 10137 13889 10149 13892
rect 10183 13889 10195 13923
rect 10137 13883 10195 13889
rect 12345 13923 12403 13929
rect 12345 13889 12357 13923
rect 12391 13920 12403 13923
rect 12452 13920 12480 14028
rect 13354 14016 13360 14028
rect 13412 14056 13418 14068
rect 14090 14056 14096 14068
rect 13412 14028 13676 14056
rect 14051 14028 14096 14056
rect 13412 14016 13418 14028
rect 12618 13920 12624 13932
rect 12391 13892 12480 13920
rect 12579 13892 12624 13920
rect 12391 13889 12403 13892
rect 12345 13883 12403 13889
rect 12618 13880 12624 13892
rect 12676 13880 12682 13932
rect 13648 13920 13676 14028
rect 14090 14016 14096 14028
rect 14148 14016 14154 14068
rect 14366 14016 14372 14068
rect 14424 14056 14430 14068
rect 14461 14059 14519 14065
rect 14461 14056 14473 14059
rect 14424 14028 14473 14056
rect 14424 14016 14430 14028
rect 14461 14025 14473 14028
rect 14507 14025 14519 14059
rect 14461 14019 14519 14025
rect 14366 13920 14372 13932
rect 13648 13892 14372 13920
rect 14366 13880 14372 13892
rect 14424 13920 14430 13932
rect 15013 13923 15071 13929
rect 15013 13920 15025 13923
rect 14424 13892 15025 13920
rect 14424 13880 14430 13892
rect 15013 13889 15025 13892
rect 15059 13889 15071 13923
rect 15286 13920 15292 13932
rect 15247 13892 15292 13920
rect 15013 13883 15071 13889
rect 15286 13880 15292 13892
rect 15344 13880 15350 13932
rect 15654 13880 15660 13932
rect 15712 13920 15718 13932
rect 16761 13923 16819 13929
rect 16761 13920 16773 13923
rect 15712 13892 16773 13920
rect 15712 13880 15718 13892
rect 16761 13889 16773 13892
rect 16807 13889 16819 13923
rect 16761 13883 16819 13889
rect 9217 13855 9275 13861
rect 9217 13852 9229 13855
rect 8435 13824 8616 13852
rect 8680 13824 9229 13852
rect 8435 13821 8447 13824
rect 8389 13815 8447 13821
rect 5534 13784 5540 13796
rect 5495 13756 5540 13784
rect 5534 13744 5540 13756
rect 5592 13744 5598 13796
rect 5810 13793 5816 13796
rect 5629 13787 5687 13793
rect 5629 13753 5641 13787
rect 5675 13753 5687 13787
rect 5629 13747 5687 13753
rect 5767 13787 5816 13793
rect 5767 13753 5779 13787
rect 5813 13753 5816 13787
rect 5767 13747 5816 13753
rect 3418 13676 3424 13728
rect 3476 13716 3482 13728
rect 4062 13716 4068 13728
rect 3476 13688 4068 13716
rect 3476 13676 3482 13688
rect 4062 13676 4068 13688
rect 4120 13716 4126 13728
rect 4430 13716 4436 13728
rect 4120 13688 4436 13716
rect 4120 13676 4126 13688
rect 4430 13676 4436 13688
rect 4488 13716 4494 13728
rect 5644 13716 5672 13747
rect 5810 13744 5816 13747
rect 5868 13744 5874 13796
rect 6196 13784 6224 13815
rect 6012 13756 6224 13784
rect 8588 13784 8616 13824
rect 9217 13821 9229 13824
rect 9263 13821 9275 13855
rect 9217 13815 9275 13821
rect 9582 13855 9640 13861
rect 9582 13821 9594 13855
rect 9628 13852 9640 13855
rect 10042 13852 10048 13864
rect 9628 13824 10048 13852
rect 9628 13821 9640 13824
rect 9582 13815 9640 13821
rect 10042 13812 10048 13824
rect 10100 13852 10106 13864
rect 10318 13852 10324 13864
rect 10100 13824 10145 13852
rect 10279 13824 10324 13852
rect 10100 13812 10106 13824
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 10597 13855 10655 13861
rect 10597 13821 10609 13855
rect 10643 13852 10655 13855
rect 10689 13855 10747 13861
rect 10689 13852 10701 13855
rect 10643 13824 10701 13852
rect 10643 13821 10655 13824
rect 10597 13815 10655 13821
rect 10689 13821 10701 13824
rect 10735 13852 10747 13855
rect 10778 13852 10784 13864
rect 10735 13824 10784 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 10778 13812 10784 13824
rect 10836 13812 10842 13864
rect 10873 13855 10931 13861
rect 10873 13821 10885 13855
rect 10919 13821 10931 13855
rect 10873 13815 10931 13821
rect 14645 13855 14703 13861
rect 14645 13821 14657 13855
rect 14691 13821 14703 13855
rect 14918 13852 14924 13864
rect 14879 13824 14924 13852
rect 14645 13815 14703 13821
rect 9033 13787 9091 13793
rect 9033 13784 9045 13787
rect 8588 13756 9045 13784
rect 6012 13728 6040 13756
rect 9033 13753 9045 13756
rect 9079 13753 9091 13787
rect 9033 13747 9091 13753
rect 10505 13787 10563 13793
rect 10505 13753 10517 13787
rect 10551 13784 10563 13787
rect 10888 13784 10916 13815
rect 10962 13784 10968 13796
rect 10551 13756 10968 13784
rect 10551 13753 10563 13756
rect 10505 13747 10563 13753
rect 10962 13744 10968 13756
rect 11020 13784 11026 13796
rect 12894 13784 12900 13796
rect 11020 13756 12900 13784
rect 11020 13744 11026 13756
rect 12894 13744 12900 13756
rect 12952 13744 12958 13796
rect 13354 13744 13360 13796
rect 13412 13744 13418 13796
rect 14660 13784 14688 13815
rect 14918 13812 14924 13824
rect 14976 13812 14982 13864
rect 15378 13784 15384 13796
rect 14660 13756 15384 13784
rect 15378 13744 15384 13756
rect 15436 13744 15442 13796
rect 16298 13744 16304 13796
rect 16356 13744 16362 13796
rect 4488 13688 5672 13716
rect 4488 13676 4494 13688
rect 5994 13676 6000 13728
rect 6052 13676 6058 13728
rect 9585 13719 9643 13725
rect 9585 13685 9597 13719
rect 9631 13716 9643 13719
rect 9950 13716 9956 13728
rect 9631 13688 9956 13716
rect 9631 13685 9643 13688
rect 9585 13679 9643 13685
rect 9950 13676 9956 13688
rect 10008 13676 10014 13728
rect 14274 13676 14280 13728
rect 14332 13716 14338 13728
rect 14734 13716 14740 13728
rect 14332 13688 14740 13716
rect 14332 13676 14338 13688
rect 14734 13676 14740 13688
rect 14792 13716 14798 13728
rect 14829 13719 14887 13725
rect 14829 13716 14841 13719
rect 14792 13688 14841 13716
rect 14792 13676 14798 13688
rect 14829 13685 14841 13688
rect 14875 13685 14887 13719
rect 14829 13679 14887 13685
rect 1104 13626 17296 13648
rect 1104 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 6571 13626
rect 6623 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 11904 13626
rect 11956 13574 11968 13626
rect 12020 13574 17296 13626
rect 1104 13552 17296 13574
rect 4246 13472 4252 13524
rect 4304 13512 4310 13524
rect 5442 13512 5448 13524
rect 4304 13484 5448 13512
rect 4304 13472 4310 13484
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 6365 13515 6423 13521
rect 6365 13512 6377 13515
rect 5592 13484 6377 13512
rect 5592 13472 5598 13484
rect 6365 13481 6377 13484
rect 6411 13481 6423 13515
rect 6365 13475 6423 13481
rect 3510 13444 3516 13456
rect 3471 13416 3516 13444
rect 3510 13404 3516 13416
rect 3568 13404 3574 13456
rect 4264 13444 4292 13472
rect 4706 13444 4712 13456
rect 4172 13416 4292 13444
rect 4667 13416 4712 13444
rect 2130 13336 2136 13388
rect 2188 13376 2194 13388
rect 2225 13379 2283 13385
rect 2225 13376 2237 13379
rect 2188 13348 2237 13376
rect 2188 13336 2194 13348
rect 2225 13345 2237 13348
rect 2271 13345 2283 13379
rect 2225 13339 2283 13345
rect 3697 13379 3755 13385
rect 3697 13345 3709 13379
rect 3743 13376 3755 13379
rect 4062 13376 4068 13388
rect 3743 13348 3924 13376
rect 4023 13348 4068 13376
rect 3743 13345 3755 13348
rect 3697 13339 3755 13345
rect 1946 13132 1952 13184
rect 2004 13172 2010 13184
rect 2041 13175 2099 13181
rect 2041 13172 2053 13175
rect 2004 13144 2053 13172
rect 2004 13132 2010 13144
rect 2041 13141 2053 13144
rect 2087 13141 2099 13175
rect 2041 13135 2099 13141
rect 3329 13175 3387 13181
rect 3329 13141 3341 13175
rect 3375 13172 3387 13175
rect 3510 13172 3516 13184
rect 3375 13144 3516 13172
rect 3375 13141 3387 13144
rect 3329 13135 3387 13141
rect 3510 13132 3516 13144
rect 3568 13132 3574 13184
rect 3896 13181 3924 13348
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 4172 13385 4200 13416
rect 4706 13404 4712 13416
rect 4764 13404 4770 13456
rect 4157 13379 4215 13385
rect 4157 13345 4169 13379
rect 4203 13345 4215 13379
rect 4157 13339 4215 13345
rect 4246 13336 4252 13388
rect 4304 13376 4310 13388
rect 4433 13379 4491 13385
rect 4433 13376 4445 13379
rect 4304 13348 4445 13376
rect 4304 13336 4310 13348
rect 4433 13345 4445 13348
rect 4479 13345 4491 13379
rect 4890 13376 4896 13388
rect 4851 13348 4896 13376
rect 4433 13339 4491 13345
rect 4890 13336 4896 13348
rect 4948 13336 4954 13388
rect 5994 13376 6000 13388
rect 5955 13348 6000 13376
rect 5994 13336 6000 13348
rect 6052 13336 6058 13388
rect 6086 13336 6092 13388
rect 6144 13376 6150 13388
rect 6181 13379 6239 13385
rect 6181 13376 6193 13379
rect 6144 13348 6193 13376
rect 6144 13336 6150 13348
rect 6181 13345 6193 13348
rect 6227 13345 6239 13379
rect 6181 13339 6239 13345
rect 4338 13308 4344 13320
rect 4299 13280 4344 13308
rect 4338 13268 4344 13280
rect 4396 13268 4402 13320
rect 3970 13200 3976 13252
rect 4028 13240 4034 13252
rect 4525 13243 4583 13249
rect 4525 13240 4537 13243
rect 4028 13212 4537 13240
rect 4028 13200 4034 13212
rect 4525 13209 4537 13212
rect 4571 13209 4583 13243
rect 6196 13240 6224 13339
rect 6380 13308 6408 13475
rect 7834 13472 7840 13524
rect 7892 13512 7898 13524
rect 10689 13515 10747 13521
rect 10689 13512 10701 13515
rect 7892 13484 10701 13512
rect 7892 13472 7898 13484
rect 10689 13481 10701 13484
rect 10735 13481 10747 13515
rect 10689 13475 10747 13481
rect 12710 13472 12716 13524
rect 12768 13512 12774 13524
rect 12897 13515 12955 13521
rect 12897 13512 12909 13515
rect 12768 13484 12909 13512
rect 12768 13472 12774 13484
rect 12897 13481 12909 13484
rect 12943 13481 12955 13515
rect 12897 13475 12955 13481
rect 13354 13472 13360 13524
rect 13412 13512 13418 13524
rect 13449 13515 13507 13521
rect 13449 13512 13461 13515
rect 13412 13484 13461 13512
rect 13412 13472 13418 13484
rect 13449 13481 13461 13484
rect 13495 13481 13507 13515
rect 16298 13512 16304 13524
rect 16259 13484 16304 13512
rect 13449 13475 13507 13481
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 6457 13447 6515 13453
rect 6457 13413 6469 13447
rect 6503 13444 6515 13447
rect 6503 13416 7696 13444
rect 6503 13413 6515 13416
rect 6457 13407 6515 13413
rect 7668 13388 7696 13416
rect 12250 13404 12256 13456
rect 12308 13444 12314 13456
rect 12989 13447 13047 13453
rect 12989 13444 13001 13447
rect 12308 13416 13001 13444
rect 12308 13404 12314 13416
rect 12989 13413 13001 13416
rect 13035 13444 13047 13447
rect 13538 13444 13544 13456
rect 13035 13416 13544 13444
rect 13035 13413 13047 13416
rect 12989 13407 13047 13413
rect 13538 13404 13544 13416
rect 13596 13444 13602 13456
rect 15194 13444 15200 13456
rect 13596 13416 15200 13444
rect 13596 13404 13602 13416
rect 15194 13404 15200 13416
rect 15252 13404 15258 13456
rect 6730 13376 6736 13388
rect 6691 13348 6736 13376
rect 6730 13336 6736 13348
rect 6788 13336 6794 13388
rect 7377 13379 7435 13385
rect 7377 13345 7389 13379
rect 7423 13376 7435 13379
rect 7466 13376 7472 13388
rect 7423 13348 7472 13376
rect 7423 13345 7435 13348
rect 7377 13339 7435 13345
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 7650 13336 7656 13388
rect 7708 13376 7714 13388
rect 10965 13379 11023 13385
rect 7708 13348 7801 13376
rect 7708 13336 7714 13348
rect 10965 13345 10977 13379
rect 11011 13376 11023 13379
rect 11241 13379 11299 13385
rect 11241 13376 11253 13379
rect 11011 13348 11253 13376
rect 11011 13345 11023 13348
rect 10965 13339 11023 13345
rect 11241 13345 11253 13348
rect 11287 13376 11299 13379
rect 11422 13376 11428 13388
rect 11287 13348 11428 13376
rect 11287 13345 11299 13348
rect 11241 13339 11299 13345
rect 11422 13336 11428 13348
rect 11480 13336 11486 13388
rect 11609 13379 11667 13385
rect 11609 13345 11621 13379
rect 11655 13345 11667 13379
rect 11609 13339 11667 13345
rect 12805 13379 12863 13385
rect 12805 13345 12817 13379
rect 12851 13376 12863 13379
rect 12894 13376 12900 13388
rect 12851 13348 12900 13376
rect 12851 13345 12863 13348
rect 12805 13339 12863 13345
rect 6457 13311 6515 13317
rect 6457 13308 6469 13311
rect 6380 13280 6469 13308
rect 6457 13277 6469 13280
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 6641 13311 6699 13317
rect 6641 13277 6653 13311
rect 6687 13308 6699 13311
rect 6822 13308 6828 13320
rect 6687 13280 6828 13308
rect 6687 13277 6699 13280
rect 6641 13271 6699 13277
rect 6546 13240 6552 13252
rect 6196 13212 6552 13240
rect 4525 13203 4583 13209
rect 6546 13200 6552 13212
rect 6604 13200 6610 13252
rect 3881 13175 3939 13181
rect 3881 13141 3893 13175
rect 3927 13172 3939 13175
rect 4062 13172 4068 13184
rect 3927 13144 4068 13172
rect 3927 13141 3939 13144
rect 3881 13135 3939 13141
rect 4062 13132 4068 13144
rect 4120 13132 4126 13184
rect 4246 13132 4252 13184
rect 4304 13172 4310 13184
rect 4614 13172 4620 13184
rect 4304 13144 4620 13172
rect 4304 13132 4310 13144
rect 4614 13132 4620 13144
rect 4672 13172 4678 13184
rect 4982 13172 4988 13184
rect 4672 13144 4988 13172
rect 4672 13132 4678 13144
rect 4982 13132 4988 13144
rect 5040 13172 5046 13184
rect 5902 13172 5908 13184
rect 5040 13144 5908 13172
rect 5040 13132 5046 13144
rect 5902 13132 5908 13144
rect 5960 13132 5966 13184
rect 6178 13132 6184 13184
rect 6236 13172 6242 13184
rect 6656 13172 6684 13271
rect 6822 13268 6828 13280
rect 6880 13268 6886 13320
rect 10873 13311 10931 13317
rect 10873 13277 10885 13311
rect 10919 13308 10931 13311
rect 11333 13311 11391 13317
rect 11333 13308 11345 13311
rect 10919 13280 11345 13308
rect 10919 13277 10931 13280
rect 10873 13271 10931 13277
rect 11333 13277 11345 13280
rect 11379 13308 11391 13311
rect 11624 13308 11652 13339
rect 12894 13336 12900 13348
rect 12952 13336 12958 13388
rect 13262 13376 13268 13388
rect 13223 13348 13268 13376
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 14734 13336 14740 13388
rect 14792 13376 14798 13388
rect 14921 13379 14979 13385
rect 14921 13376 14933 13379
rect 14792 13348 14933 13376
rect 14792 13336 14798 13348
rect 14921 13345 14933 13348
rect 14967 13345 14979 13379
rect 14921 13339 14979 13345
rect 15010 13336 15016 13388
rect 15068 13376 15074 13388
rect 15105 13379 15163 13385
rect 15105 13376 15117 13379
rect 15068 13348 15117 13376
rect 15068 13336 15074 13348
rect 15105 13345 15117 13348
rect 15151 13376 15163 13379
rect 15473 13379 15531 13385
rect 15473 13376 15485 13379
rect 15151 13348 15485 13376
rect 15151 13345 15163 13348
rect 15105 13339 15163 13345
rect 15473 13345 15485 13348
rect 15519 13345 15531 13379
rect 15473 13339 15531 13345
rect 15562 13336 15568 13388
rect 15620 13376 15626 13388
rect 15620 13348 15665 13376
rect 15620 13336 15626 13348
rect 16206 13336 16212 13388
rect 16264 13376 16270 13388
rect 16482 13376 16488 13388
rect 16264 13348 16488 13376
rect 16264 13336 16270 13348
rect 16482 13336 16488 13348
rect 16540 13336 16546 13388
rect 13630 13308 13636 13320
rect 11379 13280 13636 13308
rect 11379 13277 11391 13280
rect 11333 13271 11391 13277
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 15289 13311 15347 13317
rect 15289 13277 15301 13311
rect 15335 13308 15347 13311
rect 15378 13308 15384 13320
rect 15335 13280 15384 13308
rect 15335 13277 15347 13280
rect 15289 13271 15347 13277
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 7374 13200 7380 13252
rect 7432 13240 7438 13252
rect 7745 13243 7803 13249
rect 7745 13240 7757 13243
rect 7432 13212 7757 13240
rect 7432 13200 7438 13212
rect 7745 13209 7757 13212
rect 7791 13209 7803 13243
rect 7745 13203 7803 13209
rect 12621 13243 12679 13249
rect 12621 13209 12633 13243
rect 12667 13240 12679 13243
rect 12986 13240 12992 13252
rect 12667 13212 12992 13240
rect 12667 13209 12679 13212
rect 12621 13203 12679 13209
rect 12986 13200 12992 13212
rect 13044 13200 13050 13252
rect 6236 13144 6684 13172
rect 7469 13175 7527 13181
rect 6236 13132 6242 13144
rect 7469 13141 7481 13175
rect 7515 13172 7527 13175
rect 7558 13172 7564 13184
rect 7515 13144 7564 13172
rect 7515 13141 7527 13144
rect 7469 13135 7527 13141
rect 7558 13132 7564 13144
rect 7616 13132 7622 13184
rect 11238 13132 11244 13184
rect 11296 13172 11302 13184
rect 11517 13175 11575 13181
rect 11517 13172 11529 13175
rect 11296 13144 11529 13172
rect 11296 13132 11302 13144
rect 11517 13141 11529 13144
rect 11563 13141 11575 13175
rect 11517 13135 11575 13141
rect 12710 13132 12716 13184
rect 12768 13172 12774 13184
rect 13173 13175 13231 13181
rect 13173 13172 13185 13175
rect 12768 13144 13185 13172
rect 12768 13132 12774 13144
rect 13173 13141 13185 13144
rect 13219 13141 13231 13175
rect 13173 13135 13231 13141
rect 1104 13082 17296 13104
rect 1104 13030 3680 13082
rect 3732 13030 3744 13082
rect 3796 13030 3808 13082
rect 3860 13030 3872 13082
rect 3924 13030 9078 13082
rect 9130 13030 9142 13082
rect 9194 13030 9206 13082
rect 9258 13030 9270 13082
rect 9322 13030 14475 13082
rect 14527 13030 14539 13082
rect 14591 13030 14603 13082
rect 14655 13030 14667 13082
rect 14719 13030 17296 13082
rect 1104 13008 17296 13030
rect 7006 12968 7012 12980
rect 4540 12940 7012 12968
rect 3970 12900 3976 12912
rect 3712 12872 3976 12900
rect 3237 12835 3295 12841
rect 3237 12801 3249 12835
rect 3283 12832 3295 12835
rect 3326 12832 3332 12844
rect 3283 12804 3332 12832
rect 3283 12801 3295 12804
rect 3237 12795 3295 12801
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 3510 12764 3516 12776
rect 3471 12736 3516 12764
rect 3510 12724 3516 12736
rect 3568 12724 3574 12776
rect 3605 12767 3663 12773
rect 3605 12733 3617 12767
rect 3651 12764 3663 12767
rect 3712 12764 3740 12872
rect 3970 12860 3976 12872
rect 4028 12860 4034 12912
rect 4246 12832 4252 12844
rect 3988 12804 4252 12832
rect 3988 12773 4016 12804
rect 4246 12792 4252 12804
rect 4304 12792 4310 12844
rect 3651 12736 3740 12764
rect 3973 12767 4031 12773
rect 3651 12733 3663 12736
rect 3605 12727 3663 12733
rect 3973 12733 3985 12767
rect 4019 12733 4031 12767
rect 3973 12727 4031 12733
rect 4062 12724 4068 12776
rect 4120 12764 4126 12776
rect 4120 12736 4165 12764
rect 4120 12724 4126 12736
rect 4338 12724 4344 12776
rect 4396 12764 4402 12776
rect 4433 12767 4491 12773
rect 4433 12764 4445 12767
rect 4396 12736 4445 12764
rect 4396 12724 4402 12736
rect 4433 12733 4445 12736
rect 4479 12733 4491 12767
rect 4540 12764 4568 12940
rect 7006 12928 7012 12940
rect 7064 12928 7070 12980
rect 10042 12928 10048 12980
rect 10100 12968 10106 12980
rect 10689 12971 10747 12977
rect 10689 12968 10701 12971
rect 10100 12940 10701 12968
rect 10100 12928 10106 12940
rect 10689 12937 10701 12940
rect 10735 12937 10747 12971
rect 11238 12968 11244 12980
rect 11199 12940 11244 12968
rect 10689 12931 10747 12937
rect 11238 12928 11244 12940
rect 11296 12928 11302 12980
rect 11422 12928 11428 12980
rect 11480 12968 11486 12980
rect 11701 12971 11759 12977
rect 11701 12968 11713 12971
rect 11480 12940 11713 12968
rect 11480 12928 11486 12940
rect 11701 12937 11713 12940
rect 11747 12937 11759 12971
rect 12894 12968 12900 12980
rect 12855 12940 12900 12968
rect 11701 12931 11759 12937
rect 12894 12928 12900 12940
rect 12952 12928 12958 12980
rect 14274 12928 14280 12980
rect 14332 12968 14338 12980
rect 14461 12971 14519 12977
rect 14461 12968 14473 12971
rect 14332 12940 14473 12968
rect 14332 12928 14338 12940
rect 14461 12937 14473 12940
rect 14507 12937 14519 12971
rect 14461 12931 14519 12937
rect 14826 12928 14832 12980
rect 14884 12968 14890 12980
rect 14921 12971 14979 12977
rect 14921 12968 14933 12971
rect 14884 12940 14933 12968
rect 14884 12928 14890 12940
rect 14921 12937 14933 12940
rect 14967 12937 14979 12971
rect 14921 12931 14979 12937
rect 15102 12928 15108 12980
rect 15160 12968 15166 12980
rect 16577 12971 16635 12977
rect 16577 12968 16589 12971
rect 15160 12940 16589 12968
rect 15160 12928 15166 12940
rect 16577 12937 16589 12940
rect 16623 12937 16635 12971
rect 16577 12931 16635 12937
rect 4614 12860 4620 12912
rect 4672 12900 4678 12912
rect 4801 12903 4859 12909
rect 4801 12900 4813 12903
rect 4672 12872 4813 12900
rect 4672 12860 4678 12872
rect 4801 12869 4813 12872
rect 4847 12869 4859 12903
rect 4801 12863 4859 12869
rect 5077 12903 5135 12909
rect 5077 12869 5089 12903
rect 5123 12900 5135 12903
rect 6546 12900 6552 12912
rect 5123 12872 6552 12900
rect 5123 12869 5135 12872
rect 5077 12863 5135 12869
rect 6546 12860 6552 12872
rect 6604 12860 6610 12912
rect 6822 12860 6828 12912
rect 6880 12900 6886 12912
rect 7837 12903 7895 12909
rect 6880 12872 6960 12900
rect 6880 12860 6886 12872
rect 4706 12832 4712 12844
rect 4667 12804 4712 12832
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 6270 12792 6276 12844
rect 6328 12832 6334 12844
rect 6730 12832 6736 12844
rect 6328 12804 6736 12832
rect 6328 12792 6334 12804
rect 6730 12792 6736 12804
rect 6788 12832 6794 12844
rect 6788 12804 6868 12832
rect 6788 12792 6794 12804
rect 4617 12767 4675 12773
rect 4617 12764 4629 12767
rect 4540 12736 4629 12764
rect 4433 12727 4491 12733
rect 4617 12733 4629 12736
rect 4663 12733 4675 12767
rect 4890 12764 4896 12776
rect 4803 12736 4896 12764
rect 4617 12727 4675 12733
rect 4890 12724 4896 12736
rect 4948 12724 4954 12776
rect 5442 12724 5448 12776
rect 5500 12764 5506 12776
rect 6840 12773 6868 12804
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 5500 12736 6653 12764
rect 5500 12724 5506 12736
rect 6641 12733 6653 12736
rect 6687 12733 6699 12767
rect 6641 12727 6699 12733
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12733 6883 12767
rect 6932 12764 6960 12872
rect 7837 12869 7849 12903
rect 7883 12869 7895 12903
rect 7837 12863 7895 12869
rect 7852 12832 7880 12863
rect 11514 12860 11520 12912
rect 11572 12860 11578 12912
rect 7929 12835 7987 12841
rect 7929 12832 7941 12835
rect 7852 12804 7941 12832
rect 7929 12801 7941 12804
rect 7975 12801 7987 12835
rect 8110 12832 8116 12844
rect 8071 12804 8116 12832
rect 7929 12795 7987 12801
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 8297 12835 8355 12841
rect 8297 12801 8309 12835
rect 8343 12832 8355 12835
rect 9306 12832 9312 12844
rect 8343 12804 9312 12832
rect 8343 12801 8355 12804
rect 8297 12795 8355 12801
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 11532 12832 11560 12860
rect 11256 12804 12296 12832
rect 7009 12767 7067 12773
rect 7009 12764 7021 12767
rect 6932 12736 7021 12764
rect 6825 12727 6883 12733
rect 7009 12733 7021 12736
rect 7055 12733 7067 12767
rect 7190 12764 7196 12776
rect 7151 12736 7196 12764
rect 7009 12727 7067 12733
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 7374 12773 7380 12776
rect 7341 12767 7380 12773
rect 7341 12733 7353 12767
rect 7341 12727 7380 12733
rect 7374 12724 7380 12727
rect 7432 12724 7438 12776
rect 7558 12764 7564 12776
rect 7519 12736 7564 12764
rect 7558 12724 7564 12736
rect 7616 12724 7622 12776
rect 7650 12724 7656 12776
rect 7708 12773 7714 12776
rect 7708 12764 7716 12773
rect 8202 12764 8208 12776
rect 7708 12736 7753 12764
rect 8163 12736 8208 12764
rect 7708 12727 7716 12736
rect 7708 12724 7714 12727
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 9674 12724 9680 12776
rect 9732 12724 9738 12776
rect 10870 12767 10928 12773
rect 10870 12733 10882 12767
rect 10916 12764 10928 12767
rect 11256 12764 11284 12804
rect 10916 12736 11284 12764
rect 11333 12767 11391 12773
rect 10916 12733 10928 12736
rect 10870 12727 10928 12733
rect 11333 12733 11345 12767
rect 11379 12733 11391 12767
rect 11333 12727 11391 12733
rect 11517 12767 11575 12773
rect 11517 12733 11529 12767
rect 11563 12764 11575 12767
rect 11977 12767 12035 12773
rect 11977 12764 11989 12767
rect 11563 12736 11989 12764
rect 11563 12733 11575 12736
rect 11517 12727 11575 12733
rect 11977 12733 11989 12736
rect 12023 12764 12035 12767
rect 12066 12764 12072 12776
rect 12023 12736 12072 12764
rect 12023 12733 12035 12736
rect 11977 12727 12035 12733
rect 1946 12656 1952 12708
rect 2004 12656 2010 12708
rect 2961 12699 3019 12705
rect 2961 12665 2973 12699
rect 3007 12696 3019 12699
rect 3329 12699 3387 12705
rect 3329 12696 3341 12699
rect 3007 12668 3341 12696
rect 3007 12665 3019 12668
rect 2961 12659 3019 12665
rect 3329 12665 3341 12668
rect 3375 12665 3387 12699
rect 3329 12659 3387 12665
rect 3418 12656 3424 12708
rect 3476 12696 3482 12708
rect 3878 12705 3884 12708
rect 3697 12699 3755 12705
rect 3697 12696 3709 12699
rect 3476 12668 3709 12696
rect 3476 12656 3482 12668
rect 3697 12665 3709 12668
rect 3743 12665 3755 12699
rect 3697 12659 3755 12665
rect 3835 12699 3884 12705
rect 3835 12665 3847 12699
rect 3881 12665 3884 12699
rect 3835 12659 3884 12665
rect 3850 12656 3884 12659
rect 3936 12656 3942 12708
rect 4157 12699 4215 12705
rect 4157 12665 4169 12699
rect 4203 12696 4215 12699
rect 4908 12696 4936 12724
rect 4203 12668 4936 12696
rect 4203 12665 4215 12668
rect 4157 12659 4215 12665
rect 5810 12656 5816 12708
rect 5868 12696 5874 12708
rect 6733 12699 6791 12705
rect 6733 12696 6745 12699
rect 5868 12668 6745 12696
rect 5868 12656 5874 12668
rect 6733 12665 6745 12668
rect 6779 12665 6791 12699
rect 7466 12696 7472 12708
rect 7427 12668 7472 12696
rect 6733 12659 6791 12665
rect 7466 12656 7472 12668
rect 7524 12656 7530 12708
rect 7929 12699 7987 12705
rect 7929 12665 7941 12699
rect 7975 12696 7987 12699
rect 8573 12699 8631 12705
rect 8573 12696 8585 12699
rect 7975 12668 8585 12696
rect 7975 12665 7987 12668
rect 7929 12659 7987 12665
rect 8573 12665 8585 12668
rect 8619 12665 8631 12699
rect 11348 12696 11376 12727
rect 12066 12724 12072 12736
rect 12124 12724 12130 12776
rect 12268 12773 12296 12804
rect 12253 12767 12311 12773
rect 12253 12733 12265 12767
rect 12299 12733 12311 12767
rect 12986 12764 12992 12776
rect 12947 12736 12992 12764
rect 12253 12727 12311 12733
rect 11701 12699 11759 12705
rect 11701 12696 11713 12699
rect 11348 12668 11713 12696
rect 8573 12659 8631 12665
rect 11701 12665 11713 12668
rect 11747 12696 11759 12699
rect 12161 12699 12219 12705
rect 12161 12696 12173 12699
rect 11747 12668 12173 12696
rect 11747 12665 11759 12668
rect 11701 12659 11759 12665
rect 12161 12665 12173 12668
rect 12207 12665 12219 12699
rect 12161 12659 12219 12665
rect 1489 12631 1547 12637
rect 1489 12597 1501 12631
rect 1535 12628 1547 12631
rect 3850 12628 3878 12656
rect 1535 12600 3878 12628
rect 1535 12597 1547 12600
rect 1489 12591 1547 12597
rect 5994 12588 6000 12640
rect 6052 12628 6058 12640
rect 6457 12631 6515 12637
rect 6457 12628 6469 12631
rect 6052 12600 6469 12628
rect 6052 12588 6058 12600
rect 6457 12597 6469 12600
rect 6503 12628 6515 12631
rect 6822 12628 6828 12640
rect 6503 12600 6828 12628
rect 6503 12597 6515 12600
rect 6457 12591 6515 12597
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 9398 12588 9404 12640
rect 9456 12628 9462 12640
rect 10045 12631 10103 12637
rect 10045 12628 10057 12631
rect 9456 12600 10057 12628
rect 9456 12588 9462 12600
rect 10045 12597 10057 12600
rect 10091 12597 10103 12631
rect 10045 12591 10103 12597
rect 10873 12631 10931 12637
rect 10873 12597 10885 12631
rect 10919 12628 10931 12631
rect 11517 12631 11575 12637
rect 11517 12628 11529 12631
rect 10919 12600 11529 12628
rect 10919 12597 10931 12600
rect 10873 12591 10931 12597
rect 11517 12597 11529 12600
rect 11563 12597 11575 12631
rect 11517 12591 11575 12597
rect 11885 12631 11943 12637
rect 11885 12597 11897 12631
rect 11931 12628 11943 12631
rect 12268 12628 12296 12727
rect 12986 12724 12992 12736
rect 13044 12724 13050 12776
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 14369 12767 14427 12773
rect 14369 12764 14381 12767
rect 14148 12736 14381 12764
rect 14148 12724 14154 12736
rect 14369 12733 14381 12736
rect 14415 12733 14427 12767
rect 14369 12727 14427 12733
rect 14737 12767 14795 12773
rect 14737 12733 14749 12767
rect 14783 12733 14795 12767
rect 14737 12727 14795 12733
rect 14921 12767 14979 12773
rect 14921 12733 14933 12767
rect 14967 12764 14979 12767
rect 15194 12764 15200 12776
rect 14967 12736 15200 12764
rect 14967 12733 14979 12736
rect 14921 12727 14979 12733
rect 14752 12696 14780 12727
rect 15194 12724 15200 12736
rect 15252 12724 15258 12776
rect 15289 12767 15347 12773
rect 15289 12733 15301 12767
rect 15335 12764 15347 12767
rect 15378 12764 15384 12776
rect 15335 12736 15384 12764
rect 15335 12733 15347 12736
rect 15289 12727 15347 12733
rect 15304 12696 15332 12727
rect 15378 12724 15384 12736
rect 15436 12724 15442 12776
rect 16758 12764 16764 12776
rect 16719 12736 16764 12764
rect 16758 12724 16764 12736
rect 16816 12724 16822 12776
rect 14752 12668 15332 12696
rect 11931 12600 12296 12628
rect 11931 12597 11943 12600
rect 11885 12591 11943 12597
rect 1104 12538 17296 12560
rect 1104 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 6571 12538
rect 6623 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 11904 12538
rect 11956 12486 11968 12538
rect 12020 12486 17296 12538
rect 1104 12464 17296 12486
rect 6380 12396 7236 12424
rect 3881 12359 3939 12365
rect 3881 12325 3893 12359
rect 3927 12356 3939 12359
rect 3927 12328 4292 12356
rect 3927 12325 3939 12328
rect 3881 12319 3939 12325
rect 4264 12300 4292 12328
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 4154 12288 4160 12300
rect 4115 12260 4160 12288
rect 4154 12248 4160 12260
rect 4212 12248 4218 12300
rect 4246 12248 4252 12300
rect 4304 12288 4310 12300
rect 6380 12297 6408 12396
rect 6730 12356 6736 12368
rect 6656 12328 6736 12356
rect 6656 12297 6684 12328
rect 6730 12316 6736 12328
rect 6788 12316 6794 12368
rect 7208 12356 7236 12396
rect 7282 12384 7288 12436
rect 7340 12424 7346 12436
rect 7466 12424 7472 12436
rect 7340 12396 7472 12424
rect 7340 12384 7346 12396
rect 7466 12384 7472 12396
rect 7524 12384 7530 12436
rect 8202 12384 8208 12436
rect 8260 12424 8266 12436
rect 9493 12427 9551 12433
rect 9493 12424 9505 12427
rect 8260 12396 9505 12424
rect 8260 12384 8266 12396
rect 9493 12393 9505 12396
rect 9539 12393 9551 12427
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 9493 12387 9551 12393
rect 9508 12356 9536 12387
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 12986 12424 12992 12436
rect 12947 12396 12992 12424
rect 12986 12384 12992 12396
rect 13044 12384 13050 12436
rect 13630 12384 13636 12436
rect 13688 12424 13694 12436
rect 15749 12427 15807 12433
rect 15749 12424 15761 12427
rect 13688 12396 15761 12424
rect 13688 12384 13694 12396
rect 15749 12393 15761 12396
rect 15795 12393 15807 12427
rect 15749 12387 15807 12393
rect 9582 12356 9588 12368
rect 7208 12328 7604 12356
rect 9508 12328 9588 12356
rect 6365 12291 6423 12297
rect 6365 12288 6377 12291
rect 4304 12260 4397 12288
rect 6196 12260 6377 12288
rect 4304 12248 4310 12260
rect 6196 12232 6224 12260
rect 6365 12257 6377 12260
rect 6411 12257 6423 12291
rect 6365 12251 6423 12257
rect 6641 12291 6699 12297
rect 6641 12257 6653 12291
rect 6687 12257 6699 12291
rect 6822 12288 6828 12300
rect 6783 12260 6828 12288
rect 6641 12251 6699 12257
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 7282 12248 7288 12300
rect 7340 12248 7346 12300
rect 7576 12297 7604 12328
rect 9582 12316 9588 12328
rect 9640 12316 9646 12368
rect 11238 12316 11244 12368
rect 11296 12316 11302 12368
rect 14001 12359 14059 12365
rect 14001 12356 14013 12359
rect 13188 12328 14013 12356
rect 7469 12291 7527 12297
rect 7469 12257 7481 12291
rect 7515 12257 7527 12291
rect 7469 12251 7527 12257
rect 7561 12291 7619 12297
rect 7561 12257 7573 12291
rect 7607 12257 7619 12291
rect 7561 12251 7619 12257
rect 7837 12291 7895 12297
rect 7837 12257 7849 12291
rect 7883 12288 7895 12291
rect 8202 12288 8208 12300
rect 7883 12260 8208 12288
rect 7883 12257 7895 12260
rect 7837 12251 7895 12257
rect 3881 12223 3939 12229
rect 3881 12189 3893 12223
rect 3927 12220 3939 12223
rect 3970 12220 3976 12232
rect 3927 12192 3976 12220
rect 3927 12189 3939 12192
rect 3881 12183 3939 12189
rect 3970 12180 3976 12192
rect 4028 12180 4034 12232
rect 4065 12223 4123 12229
rect 4065 12189 4077 12223
rect 4111 12220 4123 12223
rect 4338 12220 4344 12232
rect 4111 12192 4344 12220
rect 4111 12189 4123 12192
rect 4065 12183 4123 12189
rect 4338 12180 4344 12192
rect 4396 12220 4402 12232
rect 5534 12220 5540 12232
rect 4396 12192 5540 12220
rect 4396 12180 4402 12192
rect 5534 12180 5540 12192
rect 5592 12220 5598 12232
rect 6178 12220 6184 12232
rect 5592 12192 6184 12220
rect 5592 12180 5598 12192
rect 6178 12180 6184 12192
rect 6236 12180 6242 12232
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12220 6791 12223
rect 7300 12220 7328 12248
rect 6779 12192 7328 12220
rect 6779 12189 6791 12192
rect 6733 12183 6791 12189
rect 6564 12152 6592 12183
rect 7374 12180 7380 12232
rect 7432 12220 7438 12232
rect 7484 12220 7512 12251
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 9398 12288 9404 12300
rect 9359 12260 9404 12288
rect 9398 12248 9404 12260
rect 9456 12248 9462 12300
rect 9490 12248 9496 12300
rect 9548 12288 9554 12300
rect 13188 12297 13216 12328
rect 9861 12291 9919 12297
rect 9861 12288 9873 12291
rect 9548 12260 9873 12288
rect 9548 12248 9554 12260
rect 9861 12257 9873 12260
rect 9907 12257 9919 12291
rect 9861 12251 9919 12257
rect 13173 12291 13231 12297
rect 13173 12257 13185 12291
rect 13219 12257 13231 12291
rect 13354 12288 13360 12300
rect 13315 12260 13360 12288
rect 13173 12251 13231 12257
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 13740 12297 13768 12328
rect 14001 12325 14013 12328
rect 14047 12356 14059 12359
rect 14090 12356 14096 12368
rect 14047 12328 14096 12356
rect 14047 12325 14059 12328
rect 14001 12319 14059 12325
rect 14090 12316 14096 12328
rect 14148 12316 14154 12368
rect 15378 12356 15384 12368
rect 15339 12328 15384 12356
rect 15378 12316 15384 12328
rect 15436 12316 15442 12368
rect 13725 12291 13783 12297
rect 13725 12257 13737 12291
rect 13771 12257 13783 12291
rect 13725 12251 13783 12257
rect 13817 12291 13875 12297
rect 13817 12257 13829 12291
rect 13863 12288 13875 12291
rect 13909 12291 13967 12297
rect 13909 12288 13921 12291
rect 13863 12260 13921 12288
rect 13863 12257 13875 12260
rect 13817 12251 13875 12257
rect 13909 12257 13921 12260
rect 13955 12288 13967 12291
rect 15194 12288 15200 12300
rect 13955 12260 15056 12288
rect 15155 12260 15200 12288
rect 13955 12257 13967 12260
rect 13909 12251 13967 12257
rect 9416 12220 9444 12248
rect 10321 12223 10379 12229
rect 10321 12220 10333 12223
rect 7432 12192 9444 12220
rect 9646 12192 10333 12220
rect 7432 12180 7438 12192
rect 7282 12152 7288 12164
rect 6564 12124 7288 12152
rect 7282 12112 7288 12124
rect 7340 12112 7346 12164
rect 9398 12112 9404 12164
rect 9456 12152 9462 12164
rect 9646 12152 9674 12192
rect 10321 12189 10333 12192
rect 10367 12189 10379 12223
rect 10321 12183 10379 12189
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12220 10655 12223
rect 11054 12220 11060 12232
rect 10643 12192 11060 12220
rect 10643 12189 10655 12192
rect 10597 12183 10655 12189
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 13372 12220 13400 12248
rect 13449 12223 13507 12229
rect 13449 12220 13461 12223
rect 13372 12192 13461 12220
rect 13449 12189 13461 12192
rect 13495 12189 13507 12223
rect 13449 12183 13507 12189
rect 13633 12223 13691 12229
rect 13633 12189 13645 12223
rect 13679 12220 13691 12223
rect 14274 12220 14280 12232
rect 13679 12192 14280 12220
rect 13679 12189 13691 12192
rect 13633 12183 13691 12189
rect 13648 12152 13676 12183
rect 13924 12164 13952 12192
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 15028 12220 15056 12260
rect 15194 12248 15200 12260
rect 15252 12248 15258 12300
rect 15470 12288 15476 12300
rect 15431 12260 15476 12288
rect 15470 12248 15476 12260
rect 15528 12248 15534 12300
rect 15565 12291 15623 12297
rect 15565 12257 15577 12291
rect 15611 12288 15623 12291
rect 15654 12288 15660 12300
rect 15611 12260 15660 12288
rect 15611 12257 15623 12260
rect 15565 12251 15623 12257
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 15488 12220 15516 12248
rect 15028 12192 15516 12220
rect 9456 12124 9674 12152
rect 13372 12124 13676 12152
rect 9456 12112 9462 12124
rect 1578 12084 1584 12096
rect 1539 12056 1584 12084
rect 1578 12044 1584 12056
rect 1636 12044 1642 12096
rect 4341 12087 4399 12093
rect 4341 12053 4353 12087
rect 4387 12084 4399 12087
rect 4706 12084 4712 12096
rect 4387 12056 4712 12084
rect 4387 12053 4399 12056
rect 4341 12047 4399 12053
rect 4706 12044 4712 12056
rect 4764 12044 4770 12096
rect 7006 12084 7012 12096
rect 6967 12056 7012 12084
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 7466 12044 7472 12096
rect 7524 12084 7530 12096
rect 7745 12087 7803 12093
rect 7745 12084 7757 12087
rect 7524 12056 7757 12084
rect 7524 12044 7530 12056
rect 7745 12053 7757 12056
rect 7791 12053 7803 12087
rect 7745 12047 7803 12053
rect 11330 12044 11336 12096
rect 11388 12084 11394 12096
rect 12066 12084 12072 12096
rect 11388 12056 12072 12084
rect 11388 12044 11394 12056
rect 12066 12044 12072 12056
rect 12124 12044 12130 12096
rect 13372 12093 13400 12124
rect 13906 12112 13912 12164
rect 13964 12112 13970 12164
rect 13357 12087 13415 12093
rect 13357 12053 13369 12087
rect 13403 12053 13415 12087
rect 13357 12047 13415 12053
rect 13446 12044 13452 12096
rect 13504 12084 13510 12096
rect 13541 12087 13599 12093
rect 13541 12084 13553 12087
rect 13504 12056 13553 12084
rect 13504 12044 13510 12056
rect 13541 12053 13553 12056
rect 13587 12053 13599 12087
rect 13541 12047 13599 12053
rect 13722 12044 13728 12096
rect 13780 12084 13786 12096
rect 13817 12087 13875 12093
rect 13817 12084 13829 12087
rect 13780 12056 13829 12084
rect 13780 12044 13786 12056
rect 13817 12053 13829 12056
rect 13863 12053 13875 12087
rect 13817 12047 13875 12053
rect 1104 11994 17296 12016
rect 1104 11942 3680 11994
rect 3732 11942 3744 11994
rect 3796 11942 3808 11994
rect 3860 11942 3872 11994
rect 3924 11942 9078 11994
rect 9130 11942 9142 11994
rect 9194 11942 9206 11994
rect 9258 11942 9270 11994
rect 9322 11942 14475 11994
rect 14527 11942 14539 11994
rect 14591 11942 14603 11994
rect 14655 11942 14667 11994
rect 14719 11942 17296 11994
rect 1104 11920 17296 11942
rect 4430 11840 4436 11892
rect 4488 11880 4494 11892
rect 8110 11880 8116 11892
rect 4488 11852 8116 11880
rect 4488 11840 4494 11852
rect 8110 11840 8116 11852
rect 8168 11840 8174 11892
rect 13354 11880 13360 11892
rect 12406 11852 13216 11880
rect 13315 11852 13360 11880
rect 5074 11772 5080 11824
rect 5132 11812 5138 11824
rect 12406 11812 12434 11852
rect 5132 11784 12434 11812
rect 5132 11772 5138 11784
rect 12986 11772 12992 11824
rect 13044 11772 13050 11824
rect 13188 11812 13216 11852
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 15381 11883 15439 11889
rect 15381 11880 15393 11883
rect 15252 11852 15393 11880
rect 15252 11840 15258 11852
rect 15381 11849 15393 11852
rect 15427 11849 15439 11883
rect 15381 11843 15439 11849
rect 16577 11815 16635 11821
rect 16577 11812 16589 11815
rect 13188 11784 16589 11812
rect 16577 11781 16589 11784
rect 16623 11781 16635 11815
rect 16577 11775 16635 11781
rect 5000 11716 6776 11744
rect 5000 11688 5028 11716
rect 4246 11636 4252 11688
rect 4304 11676 4310 11688
rect 4387 11679 4445 11685
rect 4387 11676 4399 11679
rect 4304 11648 4399 11676
rect 4304 11636 4310 11648
rect 4387 11645 4399 11648
rect 4433 11645 4445 11679
rect 4614 11676 4620 11688
rect 4575 11648 4620 11676
rect 4387 11639 4445 11645
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 4706 11636 4712 11688
rect 4764 11685 4770 11688
rect 4764 11679 4803 11685
rect 4791 11645 4803 11679
rect 4764 11639 4803 11645
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11676 4951 11679
rect 4982 11676 4988 11688
rect 4939 11648 4988 11676
rect 4939 11645 4951 11648
rect 4893 11639 4951 11645
rect 4764 11636 4770 11639
rect 4982 11636 4988 11648
rect 5040 11636 5046 11688
rect 5166 11676 5172 11688
rect 5079 11648 5172 11676
rect 4525 11611 4583 11617
rect 4525 11577 4537 11611
rect 4571 11577 4583 11611
rect 4632 11608 4660 11636
rect 5092 11608 5120 11648
rect 5166 11636 5172 11648
rect 5224 11636 5230 11688
rect 6748 11685 6776 11716
rect 7024 11716 7512 11744
rect 7024 11688 7052 11716
rect 6733 11679 6791 11685
rect 6733 11645 6745 11679
rect 6779 11645 6791 11679
rect 6733 11639 6791 11645
rect 6822 11636 6828 11688
rect 6880 11676 6886 11688
rect 7006 11676 7012 11688
rect 6880 11648 6925 11676
rect 6967 11648 7012 11676
rect 6880 11636 6886 11648
rect 7006 11636 7012 11648
rect 7064 11636 7070 11688
rect 7190 11676 7196 11688
rect 7248 11685 7254 11688
rect 7484 11685 7512 11716
rect 12250 11704 12256 11756
rect 12308 11744 12314 11756
rect 12805 11747 12863 11753
rect 12805 11744 12817 11747
rect 12308 11716 12817 11744
rect 12308 11704 12314 11716
rect 12805 11713 12817 11716
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 12897 11747 12955 11753
rect 12897 11713 12909 11747
rect 12943 11744 12955 11747
rect 13004 11744 13032 11772
rect 13446 11744 13452 11756
rect 12943 11716 13032 11744
rect 13188 11716 13452 11744
rect 12943 11713 12955 11716
rect 12897 11707 12955 11713
rect 7156 11648 7196 11676
rect 7190 11636 7196 11648
rect 7248 11639 7256 11685
rect 7469 11679 7527 11685
rect 7469 11645 7481 11679
rect 7515 11645 7527 11679
rect 9490 11676 9496 11688
rect 9403 11648 9496 11676
rect 7469 11639 7527 11645
rect 7248 11636 7254 11639
rect 9490 11636 9496 11648
rect 9548 11676 9554 11688
rect 11606 11676 11612 11688
rect 9548 11648 11612 11676
rect 9548 11636 9554 11648
rect 11606 11636 11612 11648
rect 11664 11636 11670 11688
rect 12710 11676 12716 11688
rect 12671 11648 12716 11676
rect 12710 11636 12716 11648
rect 12768 11636 12774 11688
rect 12989 11679 13047 11685
rect 12989 11645 13001 11679
rect 13035 11676 13047 11679
rect 13188 11676 13216 11716
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 13817 11747 13875 11753
rect 13817 11713 13829 11747
rect 13863 11744 13875 11747
rect 13998 11744 14004 11756
rect 13863 11716 14004 11744
rect 13863 11713 13875 11716
rect 13817 11707 13875 11713
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 15470 11704 15476 11756
rect 15528 11744 15534 11756
rect 15528 11716 16068 11744
rect 15528 11704 15534 11716
rect 13035 11648 13216 11676
rect 13265 11679 13323 11685
rect 13035 11645 13047 11648
rect 12989 11639 13047 11645
rect 13265 11645 13277 11679
rect 13311 11645 13323 11679
rect 13538 11676 13544 11688
rect 13499 11648 13544 11676
rect 13265 11639 13323 11645
rect 4632 11580 5120 11608
rect 7101 11611 7159 11617
rect 4525 11571 4583 11577
rect 7101 11577 7113 11611
rect 7147 11608 7159 11611
rect 7561 11611 7619 11617
rect 7561 11608 7573 11611
rect 7147 11580 7573 11608
rect 7147 11577 7159 11580
rect 7101 11571 7159 11577
rect 7561 11577 7573 11580
rect 7607 11577 7619 11611
rect 7561 11571 7619 11577
rect 4249 11543 4307 11549
rect 4249 11509 4261 11543
rect 4295 11540 4307 11543
rect 4430 11540 4436 11552
rect 4295 11512 4436 11540
rect 4295 11509 4307 11512
rect 4249 11503 4307 11509
rect 4430 11500 4436 11512
rect 4488 11500 4494 11552
rect 4540 11540 4568 11571
rect 11514 11568 11520 11620
rect 11572 11608 11578 11620
rect 13280 11608 13308 11639
rect 13538 11636 13544 11648
rect 13596 11636 13602 11688
rect 13722 11676 13728 11688
rect 13683 11648 13728 11676
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 13906 11676 13912 11688
rect 13867 11648 13912 11676
rect 13906 11636 13912 11648
rect 13964 11636 13970 11688
rect 14090 11676 14096 11688
rect 14051 11648 14096 11676
rect 14090 11636 14096 11648
rect 14148 11636 14154 11688
rect 15580 11685 15608 11716
rect 16040 11688 16068 11716
rect 14553 11679 14611 11685
rect 14553 11676 14565 11679
rect 14200 11648 14565 11676
rect 11572 11580 13308 11608
rect 11572 11568 11578 11580
rect 13354 11568 13360 11620
rect 13412 11608 13418 11620
rect 14200 11608 14228 11648
rect 14553 11645 14565 11648
rect 14599 11645 14611 11679
rect 14553 11639 14611 11645
rect 15562 11679 15620 11685
rect 15562 11645 15574 11679
rect 15608 11645 15620 11679
rect 15562 11639 15620 11645
rect 15933 11679 15991 11685
rect 15933 11645 15945 11679
rect 15979 11645 15991 11679
rect 15933 11639 15991 11645
rect 13412 11580 14228 11608
rect 14277 11611 14335 11617
rect 13412 11568 13418 11580
rect 14277 11577 14289 11611
rect 14323 11608 14335 11611
rect 14369 11611 14427 11617
rect 14369 11608 14381 11611
rect 14323 11580 14381 11608
rect 14323 11577 14335 11580
rect 14277 11571 14335 11577
rect 14369 11577 14381 11580
rect 14415 11577 14427 11611
rect 15654 11608 15660 11620
rect 15567 11580 15660 11608
rect 14369 11571 14427 11577
rect 5077 11543 5135 11549
rect 5077 11540 5089 11543
rect 4540 11512 5089 11540
rect 5077 11509 5089 11512
rect 5123 11509 5135 11543
rect 5077 11503 5135 11509
rect 7377 11543 7435 11549
rect 7377 11509 7389 11543
rect 7423 11540 7435 11543
rect 7742 11540 7748 11552
rect 7423 11512 7748 11540
rect 7423 11509 7435 11512
rect 7377 11503 7435 11509
rect 7742 11500 7748 11512
rect 7800 11500 7806 11552
rect 9674 11540 9680 11552
rect 9635 11512 9680 11540
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 13173 11543 13231 11549
rect 13173 11509 13185 11543
rect 13219 11540 13231 11543
rect 13722 11540 13728 11552
rect 13219 11512 13728 11540
rect 13219 11509 13231 11512
rect 13173 11503 13231 11509
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 14090 11500 14096 11552
rect 14148 11540 14154 11552
rect 14737 11543 14795 11549
rect 14737 11540 14749 11543
rect 14148 11512 14749 11540
rect 14148 11500 14154 11512
rect 14737 11509 14749 11512
rect 14783 11509 14795 11543
rect 14737 11503 14795 11509
rect 14826 11500 14832 11552
rect 14884 11540 14890 11552
rect 15580 11549 15608 11580
rect 15654 11568 15660 11580
rect 15712 11608 15718 11620
rect 15948 11608 15976 11639
rect 16022 11636 16028 11688
rect 16080 11676 16086 11688
rect 16080 11648 16125 11676
rect 16080 11636 16086 11648
rect 16390 11636 16396 11688
rect 16448 11676 16454 11688
rect 16761 11679 16819 11685
rect 16761 11676 16773 11679
rect 16448 11648 16773 11676
rect 16448 11636 16454 11648
rect 16761 11645 16773 11648
rect 16807 11645 16819 11679
rect 16761 11639 16819 11645
rect 15712 11580 17356 11608
rect 15712 11568 15718 11580
rect 15565 11543 15623 11549
rect 15565 11540 15577 11543
rect 14884 11512 15577 11540
rect 14884 11500 14890 11512
rect 15565 11509 15577 11512
rect 15611 11509 15623 11543
rect 15565 11503 15623 11509
rect 1104 11450 17296 11472
rect 1104 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 6571 11450
rect 6623 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 11904 11450
rect 11956 11398 11968 11450
rect 12020 11398 17296 11450
rect 1104 11376 17296 11398
rect 2501 11339 2559 11345
rect 2501 11336 2513 11339
rect 1964 11308 2513 11336
rect 1964 11277 1992 11308
rect 2501 11305 2513 11308
rect 2547 11336 2559 11339
rect 2682 11336 2688 11348
rect 2547 11308 2688 11336
rect 2547 11305 2559 11308
rect 2501 11299 2559 11305
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 5166 11336 5172 11348
rect 5127 11308 5172 11336
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 6822 11336 6828 11348
rect 6783 11308 6828 11336
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7009 11339 7067 11345
rect 7009 11305 7021 11339
rect 7055 11336 7067 11339
rect 7190 11336 7196 11348
rect 7055 11308 7196 11336
rect 7055 11305 7067 11308
rect 7009 11299 7067 11305
rect 1949 11271 2007 11277
rect 1949 11237 1961 11271
rect 1995 11237 2007 11271
rect 1949 11231 2007 11237
rect 4264 11240 5764 11268
rect 1489 11203 1547 11209
rect 1489 11169 1501 11203
rect 1535 11169 1547 11203
rect 2038 11200 2044 11212
rect 1999 11172 2044 11200
rect 1489 11163 1547 11169
rect 1504 11132 1532 11163
rect 2038 11160 2044 11172
rect 2096 11160 2102 11212
rect 4264 11209 4292 11240
rect 5736 11212 5764 11240
rect 4249 11203 4307 11209
rect 4249 11169 4261 11203
rect 4295 11169 4307 11203
rect 4249 11163 4307 11169
rect 4338 11160 4344 11212
rect 4396 11200 4402 11212
rect 5353 11203 5411 11209
rect 4396 11172 4441 11200
rect 4396 11160 4402 11172
rect 5353 11169 5365 11203
rect 5399 11169 5411 11203
rect 5353 11163 5411 11169
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11200 5503 11203
rect 5534 11200 5540 11212
rect 5491 11172 5540 11200
rect 5491 11169 5503 11172
rect 5445 11163 5503 11169
rect 2130 11132 2136 11144
rect 1504 11104 2136 11132
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 4430 11092 4436 11144
rect 4488 11132 4494 11144
rect 4525 11135 4583 11141
rect 4525 11132 4537 11135
rect 4488 11104 4537 11132
rect 4488 11092 4494 11104
rect 4525 11101 4537 11104
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 2501 11067 2559 11073
rect 2501 11033 2513 11067
rect 2547 11064 2559 11067
rect 3050 11064 3056 11076
rect 2547 11036 3056 11064
rect 2547 11033 2559 11036
rect 2501 11027 2559 11033
rect 3050 11024 3056 11036
rect 3108 11024 3114 11076
rect 4430 10956 4436 11008
rect 4488 10996 4494 11008
rect 5368 10996 5396 11163
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 5718 11160 5724 11212
rect 5776 11200 5782 11212
rect 6917 11203 6975 11209
rect 5776 11172 5869 11200
rect 5776 11160 5782 11172
rect 6917 11169 6929 11203
rect 6963 11200 6975 11203
rect 7024 11200 7052 11299
rect 7190 11296 7196 11308
rect 7248 11296 7254 11348
rect 10226 11296 10232 11348
rect 10284 11336 10290 11348
rect 10873 11339 10931 11345
rect 10873 11336 10885 11339
rect 10284 11308 10885 11336
rect 10284 11296 10290 11308
rect 10873 11305 10885 11308
rect 10919 11305 10931 11339
rect 11054 11336 11060 11348
rect 11015 11308 11060 11336
rect 10873 11299 10931 11305
rect 11054 11296 11060 11308
rect 11112 11296 11118 11348
rect 12710 11296 12716 11348
rect 12768 11336 12774 11348
rect 13354 11336 13360 11348
rect 12768 11308 13360 11336
rect 12768 11296 12774 11308
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 13538 11296 13544 11348
rect 13596 11336 13602 11348
rect 14461 11339 14519 11345
rect 14461 11336 14473 11339
rect 13596 11308 14473 11336
rect 13596 11296 13602 11308
rect 14461 11305 14473 11308
rect 14507 11305 14519 11339
rect 15105 11339 15163 11345
rect 14461 11299 14519 11305
rect 14660 11308 14964 11336
rect 7745 11271 7803 11277
rect 7208 11240 7701 11268
rect 7208 11209 7236 11240
rect 6963 11172 7052 11200
rect 7193 11203 7251 11209
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 7193 11169 7205 11203
rect 7239 11169 7251 11203
rect 7193 11163 7251 11169
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 7561 11203 7619 11209
rect 7561 11169 7573 11203
rect 7607 11169 7619 11203
rect 7673 11200 7701 11240
rect 7745 11237 7757 11271
rect 7791 11268 7803 11271
rect 9401 11271 9459 11277
rect 9401 11268 9413 11271
rect 7791 11240 9413 11268
rect 7791 11237 7803 11240
rect 7745 11231 7803 11237
rect 9401 11237 9413 11240
rect 9447 11237 9459 11271
rect 9401 11231 9459 11237
rect 9674 11228 9680 11280
rect 9732 11268 9738 11280
rect 11330 11268 11336 11280
rect 9732 11240 9890 11268
rect 11291 11240 11336 11268
rect 9732 11228 9738 11240
rect 11330 11228 11336 11240
rect 11388 11228 11394 11280
rect 11425 11271 11483 11277
rect 11425 11237 11437 11271
rect 11471 11268 11483 11271
rect 11514 11268 11520 11280
rect 11471 11240 11520 11268
rect 11471 11237 11483 11240
rect 11425 11231 11483 11237
rect 11514 11228 11520 11240
rect 11572 11268 11578 11280
rect 11977 11271 12035 11277
rect 11977 11268 11989 11271
rect 11572 11240 11989 11268
rect 11572 11228 11578 11240
rect 11977 11237 11989 11240
rect 12023 11237 12035 11271
rect 11977 11231 12035 11237
rect 12986 11228 12992 11280
rect 13044 11228 13050 11280
rect 13722 11268 13728 11280
rect 13683 11240 13728 11268
rect 13722 11228 13728 11240
rect 13780 11228 13786 11280
rect 8021 11203 8079 11209
rect 8021 11200 8033 11203
rect 7673 11172 8033 11200
rect 7561 11163 7619 11169
rect 8021 11169 8033 11172
rect 8067 11200 8079 11203
rect 8294 11200 8300 11212
rect 8067 11172 8300 11200
rect 8067 11169 8079 11172
rect 8021 11163 8079 11169
rect 5552 11132 5580 11160
rect 7300 11132 7328 11163
rect 5552 11104 7328 11132
rect 5442 11024 5448 11076
rect 5500 11064 5506 11076
rect 5629 11067 5687 11073
rect 5629 11064 5641 11067
rect 5500 11036 5641 11064
rect 5500 11024 5506 11036
rect 5629 11033 5641 11036
rect 5675 11064 5687 11067
rect 7466 11064 7472 11076
rect 5675 11036 7472 11064
rect 5675 11033 5687 11036
rect 5629 11027 5687 11033
rect 7466 11024 7472 11036
rect 7524 11024 7530 11076
rect 5902 10996 5908 11008
rect 4488 10968 4533 10996
rect 5368 10968 5908 10996
rect 4488 10956 4494 10968
rect 5902 10956 5908 10968
rect 5960 10956 5966 11008
rect 6730 10956 6736 11008
rect 6788 10996 6794 11008
rect 7576 10996 7604 11163
rect 8294 11160 8300 11172
rect 8352 11160 8358 11212
rect 11241 11203 11299 11209
rect 11241 11169 11253 11203
rect 11287 11169 11299 11203
rect 11241 11163 11299 11169
rect 11609 11203 11667 11209
rect 11609 11169 11621 11203
rect 11655 11200 11667 11203
rect 12434 11200 12440 11212
rect 11655 11172 12440 11200
rect 11655 11169 11667 11172
rect 11609 11163 11667 11169
rect 7742 11132 7748 11144
rect 7703 11104 7748 11132
rect 7742 11092 7748 11104
rect 7800 11092 7806 11144
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11132 7987 11135
rect 8110 11132 8116 11144
rect 7975 11104 8116 11132
rect 7975 11101 7987 11104
rect 7929 11095 7987 11101
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 9398 11132 9404 11144
rect 9171 11104 9404 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 9398 11092 9404 11104
rect 9456 11092 9462 11144
rect 11256 11132 11284 11163
rect 12406 11160 12440 11172
rect 12492 11160 12498 11212
rect 14093 11203 14151 11209
rect 14093 11169 14105 11203
rect 14139 11200 14151 11203
rect 14553 11203 14611 11209
rect 14553 11200 14565 11203
rect 14139 11172 14565 11200
rect 14139 11169 14151 11172
rect 14093 11163 14151 11169
rect 14553 11169 14565 11172
rect 14599 11169 14611 11203
rect 14660 11200 14688 11308
rect 14826 11268 14832 11280
rect 14787 11240 14832 11268
rect 14826 11228 14832 11240
rect 14884 11228 14890 11280
rect 14936 11268 14964 11308
rect 15105 11305 15117 11339
rect 15151 11336 15163 11339
rect 16945 11339 17003 11345
rect 15151 11308 15516 11336
rect 15151 11305 15163 11308
rect 15105 11299 15163 11305
rect 15378 11268 15384 11280
rect 14936 11240 15384 11268
rect 15378 11228 15384 11240
rect 15436 11228 15442 11280
rect 15488 11277 15516 11308
rect 16945 11305 16957 11339
rect 16991 11336 17003 11339
rect 17328 11336 17356 11580
rect 16991 11308 17356 11336
rect 16991 11305 17003 11308
rect 16945 11299 17003 11305
rect 15473 11271 15531 11277
rect 15473 11237 15485 11271
rect 15519 11237 15531 11271
rect 15473 11231 15531 11237
rect 16482 11228 16488 11280
rect 16540 11228 16546 11280
rect 14737 11203 14795 11209
rect 14737 11200 14749 11203
rect 14660 11172 14749 11200
rect 14553 11163 14611 11169
rect 14737 11169 14749 11172
rect 14783 11169 14795 11203
rect 14737 11163 14795 11169
rect 14921 11203 14979 11209
rect 14921 11169 14933 11203
rect 14967 11169 14979 11203
rect 14921 11163 14979 11169
rect 12250 11132 12256 11144
rect 11256 11104 12256 11132
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 12406 11132 12434 11160
rect 12406 11104 13952 11132
rect 13924 11064 13952 11104
rect 13998 11092 14004 11144
rect 14056 11132 14062 11144
rect 14461 11135 14519 11141
rect 14056 11104 14228 11132
rect 14056 11092 14062 11104
rect 14093 11067 14151 11073
rect 14093 11064 14105 11067
rect 13924 11036 14105 11064
rect 14093 11033 14105 11036
rect 14139 11033 14151 11067
rect 14200 11064 14228 11104
rect 14461 11101 14473 11135
rect 14507 11132 14519 11135
rect 14936 11132 14964 11163
rect 14507 11104 14964 11132
rect 15197 11135 15255 11141
rect 14507 11101 14519 11104
rect 14461 11095 14519 11101
rect 15197 11101 15209 11135
rect 15243 11101 15255 11135
rect 15197 11095 15255 11101
rect 14366 11064 14372 11076
rect 14200 11036 14372 11064
rect 14093 11027 14151 11033
rect 14366 11024 14372 11036
rect 14424 11064 14430 11076
rect 15212 11064 15240 11095
rect 14424 11036 15240 11064
rect 14424 11024 14430 11036
rect 6788 10968 7604 10996
rect 6788 10956 6794 10968
rect 1104 10906 17296 10928
rect 1104 10854 3680 10906
rect 3732 10854 3744 10906
rect 3796 10854 3808 10906
rect 3860 10854 3872 10906
rect 3924 10854 9078 10906
rect 9130 10854 9142 10906
rect 9194 10854 9206 10906
rect 9258 10854 9270 10906
rect 9322 10854 14475 10906
rect 14527 10854 14539 10906
rect 14591 10854 14603 10906
rect 14655 10854 14667 10906
rect 14719 10854 17296 10906
rect 1104 10832 17296 10854
rect 2130 10792 2136 10804
rect 2091 10764 2136 10792
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 3050 10792 3056 10804
rect 3011 10764 3056 10792
rect 3050 10752 3056 10764
rect 3108 10752 3114 10804
rect 5718 10752 5724 10804
rect 5776 10792 5782 10804
rect 7009 10795 7067 10801
rect 7009 10792 7021 10795
rect 5776 10764 7021 10792
rect 5776 10752 5782 10764
rect 7009 10761 7021 10764
rect 7055 10761 7067 10795
rect 7009 10755 7067 10761
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 11425 10795 11483 10801
rect 11425 10792 11437 10795
rect 11296 10764 11437 10792
rect 11296 10752 11302 10764
rect 11425 10761 11437 10764
rect 11471 10761 11483 10795
rect 11425 10755 11483 10761
rect 12897 10795 12955 10801
rect 12897 10761 12909 10795
rect 12943 10792 12955 10795
rect 12986 10792 12992 10804
rect 12943 10764 12992 10792
rect 12943 10761 12955 10764
rect 12897 10755 12955 10761
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 16393 10795 16451 10801
rect 16393 10761 16405 10795
rect 16439 10792 16451 10795
rect 16482 10792 16488 10804
rect 16439 10764 16488 10792
rect 16439 10761 16451 10764
rect 16393 10755 16451 10761
rect 16482 10752 16488 10764
rect 16540 10752 16546 10804
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10625 1639 10659
rect 1581 10619 1639 10625
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2222 10656 2228 10668
rect 1719 10628 2228 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 1596 10520 1624 10619
rect 2222 10616 2228 10628
rect 2280 10616 2286 10668
rect 3326 10616 3332 10668
rect 3384 10656 3390 10668
rect 4157 10659 4215 10665
rect 4157 10656 4169 10659
rect 3384 10628 4169 10656
rect 3384 10616 3390 10628
rect 4157 10625 4169 10628
rect 4203 10625 4215 10659
rect 4430 10656 4436 10668
rect 4391 10628 4436 10656
rect 4157 10619 4215 10625
rect 2682 10588 2688 10600
rect 2643 10560 2688 10588
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 1670 10520 1676 10532
rect 1596 10492 1676 10520
rect 1670 10480 1676 10492
rect 1728 10480 1734 10532
rect 2866 10520 2872 10532
rect 2827 10492 2872 10520
rect 2866 10480 2872 10492
rect 2924 10480 2930 10532
rect 4172 10520 4200 10619
rect 4430 10616 4436 10628
rect 4488 10616 4494 10668
rect 8570 10616 8576 10668
rect 8628 10656 8634 10668
rect 8665 10659 8723 10665
rect 8665 10656 8677 10659
rect 8628 10628 8677 10656
rect 8628 10616 8634 10628
rect 8665 10625 8677 10628
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10656 8907 10659
rect 9950 10656 9956 10668
rect 8895 10628 9956 10656
rect 8895 10625 8907 10628
rect 8849 10619 8907 10625
rect 9950 10616 9956 10628
rect 10008 10616 10014 10668
rect 14090 10656 14096 10668
rect 14051 10628 14096 10656
rect 14090 10616 14096 10628
rect 14148 10616 14154 10668
rect 15841 10659 15899 10665
rect 15841 10625 15853 10659
rect 15887 10656 15899 10659
rect 16022 10656 16028 10668
rect 15887 10628 16028 10656
rect 15887 10625 15899 10628
rect 15841 10619 15899 10625
rect 16022 10616 16028 10628
rect 16080 10616 16086 10668
rect 6917 10591 6975 10597
rect 6917 10588 6929 10591
rect 5920 10560 6929 10588
rect 4706 10520 4712 10532
rect 4172 10492 4712 10520
rect 4706 10480 4712 10492
rect 4764 10480 4770 10532
rect 5166 10480 5172 10532
rect 5224 10480 5230 10532
rect 5920 10464 5948 10560
rect 6917 10557 6929 10560
rect 6963 10557 6975 10591
rect 10226 10588 10232 10600
rect 10187 10560 10232 10588
rect 6917 10551 6975 10557
rect 10226 10548 10232 10560
rect 10284 10548 10290 10600
rect 11241 10591 11299 10597
rect 11241 10557 11253 10591
rect 11287 10588 11299 10591
rect 11606 10588 11612 10600
rect 11287 10560 11612 10588
rect 11287 10557 11299 10560
rect 11241 10551 11299 10557
rect 11606 10548 11612 10560
rect 11664 10588 11670 10600
rect 13081 10591 13139 10597
rect 13081 10588 13093 10591
rect 11664 10560 13093 10588
rect 11664 10548 11670 10560
rect 13081 10557 13093 10560
rect 13127 10557 13139 10591
rect 13081 10551 13139 10557
rect 13817 10591 13875 10597
rect 13817 10557 13829 10591
rect 13863 10557 13875 10591
rect 16206 10588 16212 10600
rect 16167 10560 16212 10588
rect 13817 10551 13875 10557
rect 13832 10520 13860 10551
rect 16206 10548 16212 10560
rect 16264 10548 16270 10600
rect 13998 10520 14004 10532
rect 13832 10492 14004 10520
rect 13998 10480 14004 10492
rect 14056 10480 14062 10532
rect 14826 10480 14832 10532
rect 14884 10480 14890 10532
rect 1762 10412 1768 10464
rect 1820 10452 1826 10464
rect 1820 10424 1865 10452
rect 1820 10412 1826 10424
rect 2590 10412 2596 10464
rect 2648 10452 2654 10464
rect 3145 10455 3203 10461
rect 3145 10452 3157 10455
rect 2648 10424 3157 10452
rect 2648 10412 2654 10424
rect 3145 10421 3157 10424
rect 3191 10452 3203 10455
rect 3602 10452 3608 10464
rect 3191 10424 3608 10452
rect 3191 10421 3203 10424
rect 3145 10415 3203 10421
rect 3602 10412 3608 10424
rect 3660 10412 3666 10464
rect 5902 10452 5908 10464
rect 5863 10424 5908 10452
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 7374 10452 7380 10464
rect 7064 10424 7380 10452
rect 7064 10412 7070 10424
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 8202 10452 8208 10464
rect 8163 10424 8208 10452
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8573 10455 8631 10461
rect 8573 10421 8585 10455
rect 8619 10452 8631 10455
rect 9122 10452 9128 10464
rect 8619 10424 9128 10452
rect 8619 10421 8631 10424
rect 8573 10415 8631 10421
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 9398 10412 9404 10464
rect 9456 10452 9462 10464
rect 10321 10455 10379 10461
rect 10321 10452 10333 10455
rect 9456 10424 10333 10452
rect 9456 10412 9462 10424
rect 10321 10421 10333 10424
rect 10367 10421 10379 10455
rect 10321 10415 10379 10421
rect 1104 10362 17296 10384
rect 1104 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 6571 10362
rect 6623 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 11904 10362
rect 11956 10310 11968 10362
rect 12020 10310 17296 10362
rect 1104 10288 17296 10310
rect 1486 10248 1492 10260
rect 1447 10220 1492 10248
rect 1486 10208 1492 10220
rect 1544 10208 1550 10260
rect 3602 10248 3608 10260
rect 3563 10220 3608 10248
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 5166 10208 5172 10260
rect 5224 10248 5230 10260
rect 5261 10251 5319 10257
rect 5261 10248 5273 10251
rect 5224 10220 5273 10248
rect 5224 10208 5230 10220
rect 5261 10217 5273 10220
rect 5307 10217 5319 10251
rect 5261 10211 5319 10217
rect 6270 10208 6276 10260
rect 6328 10248 6334 10260
rect 6822 10248 6828 10260
rect 6328 10220 6828 10248
rect 6328 10208 6334 10220
rect 6822 10208 6828 10220
rect 6880 10248 6886 10260
rect 7193 10251 7251 10257
rect 7193 10248 7205 10251
rect 6880 10220 7205 10248
rect 6880 10208 6886 10220
rect 7193 10217 7205 10220
rect 7239 10217 7251 10251
rect 9122 10248 9128 10260
rect 9083 10220 9128 10248
rect 7193 10211 7251 10217
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 9582 10208 9588 10260
rect 9640 10208 9646 10260
rect 14826 10208 14832 10260
rect 14884 10248 14890 10260
rect 14921 10251 14979 10257
rect 14921 10248 14933 10251
rect 14884 10220 14933 10248
rect 14884 10208 14890 10220
rect 14921 10217 14933 10220
rect 14967 10217 14979 10251
rect 14921 10211 14979 10217
rect 8202 10180 8208 10192
rect 3068 10152 4108 10180
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10081 1639 10115
rect 1581 10075 1639 10081
rect 1596 9976 1624 10075
rect 2038 10072 2044 10124
rect 2096 10112 2102 10124
rect 2593 10115 2651 10121
rect 2593 10112 2605 10115
rect 2096 10084 2605 10112
rect 2096 10072 2102 10084
rect 2593 10081 2605 10084
rect 2639 10112 2651 10115
rect 2774 10112 2780 10124
rect 2639 10084 2780 10112
rect 2639 10081 2651 10084
rect 2593 10075 2651 10081
rect 2774 10072 2780 10084
rect 2832 10112 2838 10124
rect 3068 10112 3096 10152
rect 4080 10121 4108 10152
rect 4908 10152 8208 10180
rect 2832 10084 3096 10112
rect 3145 10115 3203 10121
rect 2832 10072 2838 10084
rect 3145 10081 3157 10115
rect 3191 10112 3203 10115
rect 4065 10115 4123 10121
rect 3191 10084 3280 10112
rect 3191 10081 3203 10084
rect 3145 10075 3203 10081
rect 1762 10004 1768 10056
rect 1820 10044 1826 10056
rect 3252 10053 3280 10084
rect 4065 10081 4077 10115
rect 4111 10081 4123 10115
rect 4065 10075 4123 10081
rect 3237 10047 3295 10053
rect 1820 10016 3188 10044
rect 1820 10004 1826 10016
rect 3050 9976 3056 9988
rect 1596 9948 3056 9976
rect 3050 9936 3056 9948
rect 3108 9936 3114 9988
rect 2590 9908 2596 9920
rect 2551 9880 2596 9908
rect 2590 9868 2596 9880
rect 2648 9868 2654 9920
rect 3160 9908 3188 10016
rect 3237 10013 3249 10047
rect 3283 10044 3295 10047
rect 4908 10044 4936 10152
rect 8202 10140 8208 10152
rect 8260 10140 8266 10192
rect 9600 10180 9628 10208
rect 9600 10152 9904 10180
rect 5077 10115 5135 10121
rect 5077 10081 5089 10115
rect 5123 10112 5135 10115
rect 5350 10112 5356 10124
rect 5123 10084 5356 10112
rect 5123 10081 5135 10084
rect 5077 10075 5135 10081
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 5810 10072 5816 10124
rect 5868 10112 5874 10124
rect 6365 10115 6423 10121
rect 6365 10112 6377 10115
rect 5868 10084 6377 10112
rect 5868 10072 5874 10084
rect 6365 10081 6377 10084
rect 6411 10081 6423 10115
rect 6365 10075 6423 10081
rect 6457 10115 6515 10121
rect 6457 10081 6469 10115
rect 6503 10112 6515 10115
rect 7006 10112 7012 10124
rect 6503 10084 7012 10112
rect 6503 10081 6515 10084
rect 6457 10075 6515 10081
rect 6270 10044 6276 10056
rect 3283 10016 4936 10044
rect 6231 10016 6276 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 6270 10004 6276 10016
rect 6328 10004 6334 10056
rect 3605 9979 3663 9985
rect 3605 9945 3617 9979
rect 3651 9976 3663 9979
rect 3881 9979 3939 9985
rect 3881 9976 3893 9979
rect 3651 9948 3893 9976
rect 3651 9945 3663 9948
rect 3605 9939 3663 9945
rect 3881 9945 3893 9948
rect 3927 9945 3939 9979
rect 6380 9976 6408 10075
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 7101 10115 7159 10121
rect 7101 10081 7113 10115
rect 7147 10081 7159 10115
rect 7101 10075 7159 10081
rect 9401 10115 9459 10121
rect 9401 10081 9413 10115
rect 9447 10112 9459 10115
rect 9582 10112 9588 10124
rect 9447 10084 9588 10112
rect 9447 10081 9459 10084
rect 9401 10075 9459 10081
rect 6546 10044 6552 10056
rect 6507 10016 6552 10044
rect 6546 10004 6552 10016
rect 6604 10004 6610 10056
rect 7116 9976 7144 10075
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 9876 10121 9904 10152
rect 9861 10115 9919 10121
rect 9861 10081 9873 10115
rect 9907 10081 9919 10115
rect 9861 10075 9919 10081
rect 14737 10115 14795 10121
rect 14737 10081 14749 10115
rect 14783 10112 14795 10115
rect 16206 10112 16212 10124
rect 14783 10084 16212 10112
rect 14783 10081 14795 10084
rect 14737 10075 14795 10081
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 6380 9948 7144 9976
rect 3881 9939 3939 9945
rect 8294 9936 8300 9988
rect 8352 9976 8358 9988
rect 9398 9976 9404 9988
rect 8352 9948 9404 9976
rect 8352 9936 8358 9948
rect 9398 9936 9404 9948
rect 9456 9976 9462 9988
rect 9585 9979 9643 9985
rect 9585 9976 9597 9979
rect 9456 9948 9597 9976
rect 9456 9936 9462 9948
rect 9585 9945 9597 9948
rect 9631 9945 9643 9979
rect 9585 9939 9643 9945
rect 6089 9911 6147 9917
rect 6089 9908 6101 9911
rect 3160 9880 6101 9908
rect 6089 9877 6101 9880
rect 6135 9877 6147 9911
rect 6089 9871 6147 9877
rect 8846 9868 8852 9920
rect 8904 9908 8910 9920
rect 9493 9911 9551 9917
rect 9493 9908 9505 9911
rect 8904 9880 9505 9908
rect 8904 9868 8910 9880
rect 9493 9877 9505 9880
rect 9539 9877 9551 9911
rect 9674 9908 9680 9920
rect 9635 9880 9680 9908
rect 9493 9871 9551 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 1104 9818 17296 9840
rect 1104 9766 3680 9818
rect 3732 9766 3744 9818
rect 3796 9766 3808 9818
rect 3860 9766 3872 9818
rect 3924 9766 9078 9818
rect 9130 9766 9142 9818
rect 9194 9766 9206 9818
rect 9258 9766 9270 9818
rect 9322 9766 14475 9818
rect 14527 9766 14539 9818
rect 14591 9766 14603 9818
rect 14655 9766 14667 9818
rect 14719 9766 17296 9818
rect 1104 9744 17296 9766
rect 2774 9664 2780 9716
rect 2832 9704 2838 9716
rect 2832 9676 2877 9704
rect 2832 9664 2838 9676
rect 5902 9664 5908 9716
rect 5960 9704 5966 9716
rect 6089 9707 6147 9713
rect 6089 9704 6101 9707
rect 5960 9676 6101 9704
rect 5960 9664 5966 9676
rect 6089 9673 6101 9676
rect 6135 9704 6147 9707
rect 6730 9704 6736 9716
rect 6135 9676 6736 9704
rect 6135 9673 6147 9676
rect 6089 9667 6147 9673
rect 6730 9664 6736 9676
rect 6788 9664 6794 9716
rect 6822 9664 6828 9716
rect 6880 9704 6886 9716
rect 8021 9707 8079 9713
rect 8021 9704 8033 9707
rect 6880 9676 8033 9704
rect 6880 9664 6886 9676
rect 8021 9673 8033 9676
rect 8067 9673 8079 9707
rect 8021 9667 8079 9673
rect 9398 9664 9404 9716
rect 9456 9704 9462 9716
rect 10413 9707 10471 9713
rect 10413 9704 10425 9707
rect 9456 9676 10425 9704
rect 9456 9664 9462 9676
rect 10413 9673 10425 9676
rect 10459 9673 10471 9707
rect 10413 9667 10471 9673
rect 10502 9664 10508 9716
rect 10560 9704 10566 9716
rect 10560 9676 11836 9704
rect 10560 9664 10566 9676
rect 1670 9596 1676 9648
rect 1728 9636 1734 9648
rect 5721 9639 5779 9645
rect 5721 9636 5733 9639
rect 1728 9608 1992 9636
rect 1728 9596 1734 9608
rect 1854 9568 1860 9580
rect 1815 9540 1860 9568
rect 1854 9528 1860 9540
rect 1912 9528 1918 9580
rect 1964 9577 1992 9608
rect 2746 9608 5733 9636
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 1765 9503 1823 9509
rect 1765 9469 1777 9503
rect 1811 9500 1823 9503
rect 2746 9500 2774 9608
rect 5721 9605 5733 9608
rect 5767 9605 5779 9639
rect 5721 9599 5779 9605
rect 5994 9596 6000 9648
rect 6052 9636 6058 9648
rect 6178 9636 6184 9648
rect 6052 9608 6184 9636
rect 6052 9596 6058 9608
rect 6178 9596 6184 9608
rect 6236 9636 6242 9648
rect 6546 9636 6552 9648
rect 6236 9608 6552 9636
rect 6236 9596 6242 9608
rect 6546 9596 6552 9608
rect 6604 9596 6610 9648
rect 6914 9596 6920 9648
rect 6972 9636 6978 9648
rect 7009 9639 7067 9645
rect 7009 9636 7021 9639
rect 6972 9608 7021 9636
rect 6972 9596 6978 9608
rect 7009 9605 7021 9608
rect 7055 9636 7067 9639
rect 7834 9636 7840 9648
rect 7055 9608 7840 9636
rect 7055 9605 7067 9608
rect 7009 9599 7067 9605
rect 7834 9596 7840 9608
rect 7892 9596 7898 9648
rect 8389 9639 8447 9645
rect 8389 9605 8401 9639
rect 8435 9636 8447 9639
rect 10686 9636 10692 9648
rect 8435 9608 10692 9636
rect 8435 9605 8447 9608
rect 8389 9599 8447 9605
rect 10686 9596 10692 9608
rect 10744 9636 10750 9648
rect 11517 9639 11575 9645
rect 11517 9636 11529 9639
rect 10744 9608 11529 9636
rect 10744 9596 10750 9608
rect 11517 9605 11529 9608
rect 11563 9605 11575 9639
rect 11517 9599 11575 9605
rect 11701 9639 11759 9645
rect 11701 9605 11713 9639
rect 11747 9605 11759 9639
rect 11701 9599 11759 9605
rect 4614 9528 4620 9580
rect 4672 9568 4678 9580
rect 7190 9568 7196 9580
rect 4672 9540 7196 9568
rect 4672 9528 4678 9540
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 8113 9571 8171 9577
rect 7300 9540 7696 9568
rect 7300 9512 7328 9540
rect 3970 9500 3976 9512
rect 1811 9472 2774 9500
rect 3931 9472 3976 9500
rect 1811 9469 1823 9472
rect 1765 9463 1823 9469
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 4246 9460 4252 9512
rect 4304 9500 4310 9512
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 4304 9472 4445 9500
rect 4304 9460 4310 9472
rect 4433 9469 4445 9472
rect 4479 9469 4491 9503
rect 5258 9500 5264 9512
rect 5219 9472 5264 9500
rect 4433 9463 4491 9469
rect 5258 9460 5264 9472
rect 5316 9460 5322 9512
rect 5994 9500 6000 9512
rect 5955 9472 6000 9500
rect 5994 9460 6000 9472
rect 6052 9460 6058 9512
rect 6089 9503 6147 9509
rect 6089 9469 6101 9503
rect 6135 9500 6147 9503
rect 6181 9503 6239 9509
rect 6181 9500 6193 9503
rect 6135 9472 6193 9500
rect 6135 9469 6147 9472
rect 6089 9463 6147 9469
rect 6181 9469 6193 9472
rect 6227 9469 6239 9503
rect 6181 9463 6239 9469
rect 6270 9460 6276 9512
rect 6328 9500 6334 9512
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 6328 9472 6837 9500
rect 6328 9460 6334 9472
rect 6825 9469 6837 9472
rect 6871 9500 6883 9503
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 6871 9472 6929 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 6917 9469 6929 9472
rect 6963 9500 6975 9503
rect 7282 9500 7288 9512
rect 6963 9472 7144 9500
rect 7243 9472 7288 9500
rect 6963 9469 6975 9472
rect 6917 9463 6975 9469
rect 2314 9392 2320 9444
rect 2372 9432 2378 9444
rect 2685 9435 2743 9441
rect 2685 9432 2697 9435
rect 2372 9404 2697 9432
rect 2372 9392 2378 9404
rect 2685 9401 2697 9404
rect 2731 9401 2743 9435
rect 3988 9432 4016 9460
rect 5626 9432 5632 9444
rect 3988 9404 5632 9432
rect 2685 9395 2743 9401
rect 5626 9392 5632 9404
rect 5684 9432 5690 9444
rect 6457 9435 6515 9441
rect 6457 9432 6469 9435
rect 5684 9404 6469 9432
rect 5684 9392 5690 9404
rect 6457 9401 6469 9404
rect 6503 9401 6515 9435
rect 6457 9395 6515 9401
rect 6641 9435 6699 9441
rect 6641 9401 6653 9435
rect 6687 9432 6699 9435
rect 6730 9432 6736 9444
rect 6687 9404 6736 9432
rect 6687 9401 6699 9404
rect 6641 9395 6699 9401
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 7116 9432 7144 9472
rect 7282 9460 7288 9472
rect 7340 9460 7346 9512
rect 7558 9500 7564 9512
rect 7519 9472 7564 9500
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 7668 9500 7696 9540
rect 8113 9537 8125 9571
rect 8159 9568 8171 9571
rect 9030 9568 9036 9580
rect 8159 9540 9036 9568
rect 8159 9537 8171 9540
rect 8113 9531 8171 9537
rect 9030 9528 9036 9540
rect 9088 9568 9094 9580
rect 9490 9568 9496 9580
rect 9088 9540 9496 9568
rect 9088 9528 9094 9540
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 11057 9571 11115 9577
rect 11057 9537 11069 9571
rect 11103 9568 11115 9571
rect 11716 9568 11744 9599
rect 11103 9540 11744 9568
rect 11808 9568 11836 9676
rect 12253 9571 12311 9577
rect 12253 9568 12265 9571
rect 11808 9540 12265 9568
rect 11103 9537 11115 9540
rect 11057 9531 11115 9537
rect 12253 9537 12265 9540
rect 12299 9568 12311 9571
rect 12434 9568 12440 9580
rect 12299 9540 12440 9568
rect 12299 9537 12311 9540
rect 12253 9531 12311 9537
rect 12434 9528 12440 9540
rect 12492 9528 12498 9580
rect 12802 9568 12808 9580
rect 12763 9540 12808 9568
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 12897 9571 12955 9577
rect 12897 9537 12909 9571
rect 12943 9568 12955 9571
rect 13170 9568 13176 9580
rect 12943 9540 13176 9568
rect 12943 9537 12955 9540
rect 12897 9531 12955 9537
rect 13170 9528 13176 9540
rect 13228 9528 13234 9580
rect 15013 9571 15071 9577
rect 15013 9537 15025 9571
rect 15059 9537 15071 9571
rect 15013 9531 15071 9537
rect 15197 9571 15255 9577
rect 15197 9537 15209 9571
rect 15243 9568 15255 9571
rect 16666 9568 16672 9580
rect 15243 9540 16672 9568
rect 15243 9537 15255 9540
rect 15197 9531 15255 9537
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 7668 9472 7757 9500
rect 7745 9469 7757 9472
rect 7791 9469 7803 9503
rect 7745 9463 7803 9469
rect 7837 9503 7895 9509
rect 7837 9469 7849 9503
rect 7883 9500 7895 9503
rect 7926 9500 7932 9512
rect 7883 9472 7932 9500
rect 7883 9469 7895 9472
rect 7837 9463 7895 9469
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 8018 9460 8024 9512
rect 8076 9500 8082 9512
rect 9125 9503 9183 9509
rect 8076 9472 8121 9500
rect 8076 9460 8082 9472
rect 9125 9469 9137 9503
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 9140 9432 9168 9463
rect 9214 9460 9220 9512
rect 9272 9500 9278 9512
rect 9398 9500 9404 9512
rect 9272 9472 9317 9500
rect 9359 9472 9404 9500
rect 9272 9460 9278 9472
rect 9398 9460 9404 9472
rect 9456 9460 9462 9512
rect 10413 9503 10471 9509
rect 10413 9469 10425 9503
rect 10459 9500 10471 9503
rect 10505 9503 10563 9509
rect 10505 9500 10517 9503
rect 10459 9472 10517 9500
rect 10459 9469 10471 9472
rect 10413 9463 10471 9469
rect 10505 9469 10517 9472
rect 10551 9469 10563 9503
rect 10686 9500 10692 9512
rect 10647 9472 10692 9500
rect 10505 9463 10563 9469
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 11238 9500 11244 9512
rect 11199 9472 11244 9500
rect 11238 9460 11244 9472
rect 11296 9460 11302 9512
rect 11517 9503 11575 9509
rect 11517 9469 11529 9503
rect 11563 9500 11575 9503
rect 12069 9503 12127 9509
rect 12069 9500 12081 9503
rect 11563 9472 12081 9500
rect 11563 9469 11575 9472
rect 11517 9463 11575 9469
rect 12069 9469 12081 9472
rect 12115 9469 12127 9503
rect 12820 9500 12848 9528
rect 15028 9500 15056 9531
rect 16666 9528 16672 9540
rect 16724 9528 16730 9580
rect 16758 9500 16764 9512
rect 12820 9472 15056 9500
rect 16719 9472 16764 9500
rect 12069 9463 12127 9469
rect 16758 9460 16764 9472
rect 16816 9460 16822 9512
rect 9490 9432 9496 9444
rect 7116 9404 9496 9432
rect 9490 9392 9496 9404
rect 9548 9392 9554 9444
rect 9585 9435 9643 9441
rect 9585 9401 9597 9435
rect 9631 9432 9643 9435
rect 15289 9435 15347 9441
rect 15289 9432 15301 9435
rect 9631 9404 15301 9432
rect 9631 9401 9643 9404
rect 9585 9395 9643 9401
rect 15289 9401 15301 9404
rect 15335 9401 15347 9435
rect 15289 9395 15347 9401
rect 1394 9364 1400 9376
rect 1355 9336 1400 9364
rect 1394 9324 1400 9336
rect 1452 9324 1458 9376
rect 4065 9367 4123 9373
rect 4065 9333 4077 9367
rect 4111 9364 4123 9367
rect 4154 9364 4160 9376
rect 4111 9336 4160 9364
rect 4111 9333 4123 9336
rect 4065 9327 4123 9333
rect 4154 9324 4160 9336
rect 4212 9364 4218 9376
rect 5166 9364 5172 9376
rect 4212 9336 5172 9364
rect 4212 9324 4218 9336
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 5350 9364 5356 9376
rect 5311 9336 5356 9364
rect 5350 9324 5356 9336
rect 5408 9324 5414 9376
rect 6181 9367 6239 9373
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 6914 9364 6920 9376
rect 6227 9336 6920 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 7190 9324 7196 9376
rect 7248 9364 7254 9376
rect 8386 9364 8392 9376
rect 7248 9336 8392 9364
rect 7248 9324 7254 9336
rect 8386 9324 8392 9336
rect 8444 9364 8450 9376
rect 9398 9364 9404 9376
rect 8444 9336 9404 9364
rect 8444 9324 8450 9336
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 10597 9367 10655 9373
rect 10597 9333 10609 9367
rect 10643 9364 10655 9367
rect 11238 9364 11244 9376
rect 10643 9336 11244 9364
rect 10643 9333 10655 9336
rect 10597 9327 10655 9333
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 11425 9367 11483 9373
rect 11425 9333 11437 9367
rect 11471 9364 11483 9367
rect 11606 9364 11612 9376
rect 11471 9336 11612 9364
rect 11471 9333 11483 9336
rect 11425 9327 11483 9333
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 12158 9364 12164 9376
rect 12119 9336 12164 9364
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 12986 9324 12992 9376
rect 13044 9364 13050 9376
rect 13354 9364 13360 9376
rect 13044 9336 13089 9364
rect 13315 9336 13360 9364
rect 13044 9324 13050 9336
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 15470 9324 15476 9376
rect 15528 9364 15534 9376
rect 15657 9367 15715 9373
rect 15657 9364 15669 9367
rect 15528 9336 15669 9364
rect 15528 9324 15534 9336
rect 15657 9333 15669 9336
rect 15703 9333 15715 9367
rect 16574 9364 16580 9376
rect 16535 9336 16580 9364
rect 15657 9327 15715 9333
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 1104 9274 17296 9296
rect 1104 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 6571 9274
rect 6623 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 11904 9274
rect 11956 9222 11968 9274
rect 12020 9222 17296 9274
rect 1104 9200 17296 9222
rect 5074 9160 5080 9172
rect 5035 9132 5080 9160
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 5721 9163 5779 9169
rect 5721 9129 5733 9163
rect 5767 9160 5779 9163
rect 8018 9160 8024 9172
rect 5767 9132 8024 9160
rect 5767 9129 5779 9132
rect 5721 9123 5779 9129
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 8110 9120 8116 9172
rect 8168 9120 8174 9172
rect 8202 9120 8208 9172
rect 8260 9160 8266 9172
rect 8260 9132 9904 9160
rect 8260 9120 8266 9132
rect 5166 9052 5172 9104
rect 5224 9092 5230 9104
rect 5353 9095 5411 9101
rect 5353 9092 5365 9095
rect 5224 9064 5365 9092
rect 5224 9052 5230 9064
rect 5353 9061 5365 9064
rect 5399 9061 5411 9095
rect 5353 9055 5411 9061
rect 6914 9052 6920 9104
rect 6972 9092 6978 9104
rect 8128 9092 8156 9120
rect 6972 9064 8156 9092
rect 8849 9095 8907 9101
rect 6972 9052 6978 9064
rect 8849 9061 8861 9095
rect 8895 9092 8907 9095
rect 8938 9092 8944 9104
rect 8895 9064 8944 9092
rect 8895 9061 8907 9064
rect 8849 9055 8907 9061
rect 8938 9052 8944 9064
rect 8996 9092 9002 9104
rect 9214 9092 9220 9104
rect 8996 9064 9220 9092
rect 8996 9052 9002 9064
rect 9214 9052 9220 9064
rect 9272 9052 9278 9104
rect 9876 9092 9904 9132
rect 9950 9120 9956 9172
rect 10008 9160 10014 9172
rect 11606 9160 11612 9172
rect 10008 9132 10916 9160
rect 11567 9132 11612 9160
rect 10008 9120 10014 9132
rect 9876 9064 10180 9092
rect 2958 9024 2964 9036
rect 2919 8996 2964 9024
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 5537 9027 5595 9033
rect 5537 8993 5549 9027
rect 5583 9024 5595 9027
rect 5718 9024 5724 9036
rect 5583 8996 5724 9024
rect 5583 8993 5595 8996
rect 5537 8987 5595 8993
rect 5718 8984 5724 8996
rect 5776 9024 5782 9036
rect 6086 9024 6092 9036
rect 5776 8996 6092 9024
rect 5776 8984 5782 8996
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 6822 8984 6828 9036
rect 6880 9024 6886 9036
rect 7650 9024 7656 9036
rect 6880 8996 7656 9024
rect 6880 8984 6886 8996
rect 7650 8984 7656 8996
rect 7708 9024 7714 9036
rect 8113 9027 8171 9033
rect 8113 9024 8125 9027
rect 7708 8996 8125 9024
rect 7708 8984 7714 8996
rect 8113 8993 8125 8996
rect 8159 8993 8171 9027
rect 8113 8987 8171 8993
rect 8294 8984 8300 9036
rect 8352 9024 8358 9036
rect 8389 9027 8447 9033
rect 8389 9024 8401 9027
rect 8352 8996 8401 9024
rect 8352 8984 8358 8996
rect 8389 8993 8401 8996
rect 8435 8993 8447 9027
rect 8389 8987 8447 8993
rect 9030 8984 9036 9036
rect 9088 9024 9094 9036
rect 9125 9027 9183 9033
rect 9125 9024 9137 9027
rect 9088 8996 9137 9024
rect 9088 8984 9094 8996
rect 9125 8993 9137 8996
rect 9171 8993 9183 9027
rect 9125 8987 9183 8993
rect 9306 8984 9312 9036
rect 9364 9024 9370 9036
rect 9401 9027 9459 9033
rect 9401 9024 9413 9027
rect 9364 8996 9413 9024
rect 9364 8984 9370 8996
rect 9401 8993 9413 8996
rect 9447 8993 9459 9027
rect 9582 9024 9588 9036
rect 9543 8996 9588 9024
rect 9401 8987 9459 8993
rect 9582 8984 9588 8996
rect 9640 8984 9646 9036
rect 9766 8984 9772 9036
rect 9824 9024 9830 9036
rect 10152 9033 10180 9064
rect 9953 9027 10011 9033
rect 9953 9024 9965 9027
rect 9824 8996 9965 9024
rect 9824 8984 9830 8996
rect 9953 8993 9965 8996
rect 9999 8993 10011 9027
rect 9953 8987 10011 8993
rect 10137 9027 10195 9033
rect 10137 8993 10149 9027
rect 10183 8993 10195 9027
rect 10137 8987 10195 8993
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 9024 10563 9027
rect 10594 9024 10600 9036
rect 10551 8996 10600 9024
rect 10551 8993 10563 8996
rect 10505 8987 10563 8993
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 10781 9027 10839 9033
rect 10781 8993 10793 9027
rect 10827 8993 10839 9027
rect 10781 8987 10839 8993
rect 5074 8956 5080 8968
rect 5035 8928 5080 8956
rect 5074 8916 5080 8928
rect 5132 8916 5138 8968
rect 5166 8916 5172 8968
rect 5224 8956 5230 8968
rect 5224 8928 5269 8956
rect 5224 8916 5230 8928
rect 7374 8916 7380 8968
rect 7432 8956 7438 8968
rect 7558 8956 7564 8968
rect 7432 8928 7564 8956
rect 7432 8916 7438 8928
rect 7558 8916 7564 8928
rect 7616 8956 7622 8968
rect 8202 8956 8208 8968
rect 7616 8928 8208 8956
rect 7616 8916 7622 8928
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 10796 8956 10824 8987
rect 10888 8956 10916 9132
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 11977 9163 12035 9169
rect 11977 9129 11989 9163
rect 12023 9160 12035 9163
rect 12621 9163 12679 9169
rect 12023 9132 12434 9160
rect 12023 9129 12035 9132
rect 11977 9123 12035 9129
rect 10965 9095 11023 9101
rect 10965 9061 10977 9095
rect 11011 9092 11023 9095
rect 12158 9092 12164 9104
rect 11011 9064 12164 9092
rect 11011 9061 11023 9064
rect 10965 9055 11023 9061
rect 12158 9052 12164 9064
rect 12216 9092 12222 9104
rect 12253 9095 12311 9101
rect 12253 9092 12265 9095
rect 12216 9064 12265 9092
rect 12216 9052 12222 9064
rect 12253 9061 12265 9064
rect 12299 9061 12311 9095
rect 12406 9092 12434 9132
rect 12621 9129 12633 9163
rect 12667 9160 12679 9163
rect 12986 9160 12992 9172
rect 12667 9132 12992 9160
rect 12667 9129 12679 9132
rect 12621 9123 12679 9129
rect 12986 9120 12992 9132
rect 13044 9120 13050 9172
rect 14737 9163 14795 9169
rect 14737 9129 14749 9163
rect 14783 9129 14795 9163
rect 16114 9160 16120 9172
rect 14737 9123 14795 9129
rect 15948 9132 16120 9160
rect 12406 9064 14412 9092
rect 12253 9055 12311 9061
rect 12434 9024 12440 9036
rect 11348 8996 11652 9024
rect 12395 8996 12440 9024
rect 10962 8956 10968 8968
rect 9548 8928 10824 8956
rect 10875 8928 10968 8956
rect 9548 8916 9554 8928
rect 10962 8916 10968 8928
rect 11020 8956 11026 8968
rect 11348 8965 11376 8996
rect 11333 8959 11391 8965
rect 11333 8956 11345 8959
rect 11020 8928 11345 8956
rect 11020 8916 11026 8928
rect 11333 8925 11345 8928
rect 11379 8925 11391 8959
rect 11333 8919 11391 8925
rect 11422 8916 11428 8968
rect 11480 8956 11486 8968
rect 11517 8959 11575 8965
rect 11517 8956 11529 8959
rect 11480 8928 11529 8956
rect 11480 8916 11486 8928
rect 11517 8925 11529 8928
rect 11563 8925 11575 8959
rect 11624 8956 11652 8996
rect 12434 8984 12440 8996
rect 12492 9024 12498 9036
rect 12618 9024 12624 9036
rect 12492 8996 12624 9024
rect 12492 8984 12498 8996
rect 12618 8984 12624 8996
rect 12676 9024 12682 9036
rect 13262 9024 13268 9036
rect 12676 8996 13268 9024
rect 12676 8984 12682 8996
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 13372 9033 13400 9064
rect 13357 9027 13415 9033
rect 13357 8993 13369 9027
rect 13403 8993 13415 9027
rect 13357 8987 13415 8993
rect 13909 9027 13967 9033
rect 13909 8993 13921 9027
rect 13955 9024 13967 9027
rect 13998 9024 14004 9036
rect 13955 8996 14004 9024
rect 13955 8993 13967 8996
rect 13909 8987 13967 8993
rect 13998 8984 14004 8996
rect 14056 8984 14062 9036
rect 14384 9033 14412 9064
rect 14369 9027 14427 9033
rect 14369 8993 14381 9027
rect 14415 8993 14427 9027
rect 14369 8987 14427 8993
rect 12802 8956 12808 8968
rect 11624 8928 12808 8956
rect 11517 8919 11575 8925
rect 12802 8916 12808 8928
rect 12860 8956 12866 8968
rect 13078 8956 13084 8968
rect 12860 8928 13084 8956
rect 12860 8916 12866 8928
rect 13078 8916 13084 8928
rect 13136 8916 13142 8968
rect 13817 8959 13875 8965
rect 13817 8925 13829 8959
rect 13863 8956 13875 8959
rect 14752 8956 14780 9123
rect 15948 9101 15976 9132
rect 16114 9120 16120 9132
rect 16172 9160 16178 9172
rect 16485 9163 16543 9169
rect 16485 9160 16497 9163
rect 16172 9132 16497 9160
rect 16172 9120 16178 9132
rect 16485 9129 16497 9132
rect 16531 9129 16543 9163
rect 16485 9123 16543 9129
rect 15933 9095 15991 9101
rect 15933 9061 15945 9095
rect 15979 9061 15991 9095
rect 15933 9055 15991 9061
rect 14918 8984 14924 9036
rect 14976 9024 14982 9036
rect 15013 9027 15071 9033
rect 15013 9024 15025 9027
rect 14976 8996 15025 9024
rect 14976 8984 14982 8996
rect 15013 8993 15025 8996
rect 15059 8993 15071 9027
rect 15470 9024 15476 9036
rect 15431 8996 15476 9024
rect 15013 8987 15071 8993
rect 15470 8984 15476 8996
rect 15528 8984 15534 9036
rect 15838 8984 15844 9036
rect 15896 9024 15902 9036
rect 16025 9027 16083 9033
rect 16025 9024 16037 9027
rect 15896 8996 16037 9024
rect 15896 8984 15902 8996
rect 16025 8993 16037 8996
rect 16071 9024 16083 9027
rect 16761 9027 16819 9033
rect 16761 9024 16773 9027
rect 16071 8996 16773 9024
rect 16071 8993 16083 8996
rect 16025 8987 16083 8993
rect 16761 8993 16773 8996
rect 16807 8993 16819 9027
rect 16761 8987 16819 8993
rect 13863 8928 14780 8956
rect 15488 8956 15516 8984
rect 16117 8959 16175 8965
rect 16117 8956 16129 8959
rect 15488 8928 16129 8956
rect 13863 8925 13875 8928
rect 13817 8919 13875 8925
rect 13924 8900 13952 8928
rect 16117 8925 16129 8928
rect 16163 8925 16175 8959
rect 16117 8919 16175 8925
rect 3234 8848 3240 8900
rect 3292 8888 3298 8900
rect 9861 8891 9919 8897
rect 3292 8860 9812 8888
rect 3292 8848 3298 8860
rect 2222 8780 2228 8832
rect 2280 8820 2286 8832
rect 2869 8823 2927 8829
rect 2869 8820 2881 8823
rect 2280 8792 2881 8820
rect 2280 8780 2286 8792
rect 2869 8789 2881 8792
rect 2915 8789 2927 8823
rect 2869 8783 2927 8789
rect 3970 8780 3976 8832
rect 4028 8820 4034 8832
rect 4617 8823 4675 8829
rect 4617 8820 4629 8823
rect 4028 8792 4629 8820
rect 4028 8780 4034 8792
rect 4617 8789 4629 8792
rect 4663 8789 4675 8823
rect 4617 8783 4675 8789
rect 5810 8780 5816 8832
rect 5868 8820 5874 8832
rect 9309 8823 9367 8829
rect 9309 8820 9321 8823
rect 5868 8792 9321 8820
rect 5868 8780 5874 8792
rect 9309 8789 9321 8792
rect 9355 8820 9367 8823
rect 9674 8820 9680 8832
rect 9355 8792 9680 8820
rect 9355 8789 9367 8792
rect 9309 8783 9367 8789
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 9784 8820 9812 8860
rect 9861 8857 9873 8891
rect 9907 8888 9919 8891
rect 9907 8860 11468 8888
rect 9907 8857 9919 8860
rect 9861 8851 9919 8857
rect 11330 8820 11336 8832
rect 9784 8792 11336 8820
rect 11330 8780 11336 8792
rect 11388 8780 11394 8832
rect 11440 8820 11468 8860
rect 13906 8848 13912 8900
rect 13964 8848 13970 8900
rect 14737 8891 14795 8897
rect 14737 8857 14749 8891
rect 14783 8888 14795 8891
rect 14829 8891 14887 8897
rect 14829 8888 14841 8891
rect 14783 8860 14841 8888
rect 14783 8857 14795 8860
rect 14737 8851 14795 8857
rect 14829 8857 14841 8860
rect 14875 8857 14887 8891
rect 14829 8851 14887 8857
rect 16485 8891 16543 8897
rect 16485 8857 16497 8891
rect 16531 8888 16543 8891
rect 16577 8891 16635 8897
rect 16577 8888 16589 8891
rect 16531 8860 16589 8888
rect 16531 8857 16543 8860
rect 16485 8851 16543 8857
rect 16577 8857 16589 8860
rect 16623 8857 16635 8891
rect 16577 8851 16635 8857
rect 14366 8820 14372 8832
rect 11440 8792 14372 8820
rect 14366 8780 14372 8792
rect 14424 8780 14430 8832
rect 1104 8730 17296 8752
rect 1104 8678 3680 8730
rect 3732 8678 3744 8730
rect 3796 8678 3808 8730
rect 3860 8678 3872 8730
rect 3924 8678 9078 8730
rect 9130 8678 9142 8730
rect 9194 8678 9206 8730
rect 9258 8678 9270 8730
rect 9322 8678 14475 8730
rect 14527 8678 14539 8730
rect 14591 8678 14603 8730
rect 14655 8678 14667 8730
rect 14719 8678 17296 8730
rect 1104 8656 17296 8678
rect 1670 8576 1676 8628
rect 1728 8616 1734 8628
rect 1728 8588 4752 8616
rect 1728 8576 1734 8588
rect 2222 8548 2228 8560
rect 2183 8520 2228 8548
rect 2222 8508 2228 8520
rect 2280 8508 2286 8560
rect 3605 8551 3663 8557
rect 3605 8517 3617 8551
rect 3651 8548 3663 8551
rect 3697 8551 3755 8557
rect 3697 8548 3709 8551
rect 3651 8520 3709 8548
rect 3651 8517 3663 8520
rect 3605 8511 3663 8517
rect 3697 8517 3709 8520
rect 3743 8517 3755 8551
rect 3697 8511 3755 8517
rect 4724 8548 4752 8588
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 5353 8619 5411 8625
rect 5353 8616 5365 8619
rect 5132 8588 5365 8616
rect 5132 8576 5138 8588
rect 5353 8585 5365 8588
rect 5399 8585 5411 8619
rect 10873 8619 10931 8625
rect 10873 8616 10885 8619
rect 5353 8579 5411 8585
rect 5460 8588 10885 8616
rect 5166 8548 5172 8560
rect 4724 8520 5172 8548
rect 1394 8440 1400 8492
rect 1452 8480 1458 8492
rect 1857 8483 1915 8489
rect 1857 8480 1869 8483
rect 1452 8452 1869 8480
rect 1452 8440 1458 8452
rect 1857 8449 1869 8452
rect 1903 8449 1915 8483
rect 1857 8443 1915 8449
rect 2608 8452 3924 8480
rect 2498 8372 2504 8424
rect 2556 8412 2562 8424
rect 2608 8421 2636 8452
rect 3896 8421 3924 8452
rect 4522 8440 4528 8492
rect 4580 8480 4586 8492
rect 4724 8489 4752 8520
rect 5166 8508 5172 8520
rect 5224 8508 5230 8560
rect 4617 8483 4675 8489
rect 4617 8480 4629 8483
rect 4580 8452 4629 8480
rect 4580 8440 4586 8452
rect 4617 8449 4629 8452
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 4709 8483 4767 8489
rect 4709 8449 4721 8483
rect 4755 8449 4767 8483
rect 4709 8443 4767 8449
rect 2593 8415 2651 8421
rect 2593 8412 2605 8415
rect 2556 8384 2605 8412
rect 2556 8372 2562 8384
rect 2593 8381 2605 8384
rect 2639 8381 2651 8415
rect 2593 8375 2651 8381
rect 3145 8415 3203 8421
rect 3145 8381 3157 8415
rect 3191 8412 3203 8415
rect 3237 8415 3295 8421
rect 3237 8412 3249 8415
rect 3191 8384 3249 8412
rect 3191 8381 3203 8384
rect 3145 8375 3203 8381
rect 3237 8381 3249 8384
rect 3283 8412 3295 8415
rect 3881 8415 3939 8421
rect 3283 8384 3832 8412
rect 3283 8381 3295 8384
rect 3237 8375 3295 8381
rect 1394 8344 1400 8356
rect 1355 8316 1400 8344
rect 1394 8304 1400 8316
rect 1452 8304 1458 8356
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 2038 8344 2044 8356
rect 1627 8316 2044 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 2038 8304 2044 8316
rect 2096 8304 2102 8356
rect 2685 8347 2743 8353
rect 2685 8313 2697 8347
rect 2731 8344 2743 8347
rect 2958 8344 2964 8356
rect 2731 8316 2964 8344
rect 2731 8313 2743 8316
rect 2685 8307 2743 8313
rect 2958 8304 2964 8316
rect 3016 8344 3022 8356
rect 3804 8344 3832 8384
rect 3881 8381 3893 8415
rect 3927 8381 3939 8415
rect 3881 8375 3939 8381
rect 5460 8344 5488 8588
rect 10873 8585 10885 8588
rect 10919 8585 10931 8619
rect 10873 8579 10931 8585
rect 5718 8548 5724 8560
rect 5552 8520 5724 8548
rect 5552 8489 5580 8520
rect 5718 8508 5724 8520
rect 5776 8508 5782 8560
rect 6086 8548 6092 8560
rect 6047 8520 6092 8548
rect 6086 8508 6092 8520
rect 6144 8508 6150 8560
rect 8113 8551 8171 8557
rect 8113 8548 8125 8551
rect 7484 8520 8125 8548
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8449 5595 8483
rect 5537 8443 5595 8449
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 5813 8483 5871 8489
rect 5684 8452 5729 8480
rect 5684 8440 5690 8452
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 6273 8483 6331 8489
rect 5859 8452 6224 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 5718 8372 5724 8424
rect 5776 8412 5782 8424
rect 5994 8412 6000 8424
rect 5776 8384 5821 8412
rect 5955 8384 6000 8412
rect 5776 8372 5782 8384
rect 5994 8372 6000 8384
rect 6052 8372 6058 8424
rect 6196 8412 6224 8452
rect 6273 8449 6285 8483
rect 6319 8480 6331 8483
rect 7009 8483 7067 8489
rect 7009 8480 7021 8483
rect 6319 8452 7021 8480
rect 6319 8449 6331 8452
rect 6273 8443 6331 8449
rect 7009 8449 7021 8452
rect 7055 8480 7067 8483
rect 7374 8480 7380 8492
rect 7055 8452 7380 8480
rect 7055 8449 7067 8452
rect 7009 8443 7067 8449
rect 7374 8440 7380 8452
rect 7432 8480 7438 8492
rect 7484 8489 7512 8520
rect 8113 8517 8125 8520
rect 8159 8517 8171 8551
rect 8113 8511 8171 8517
rect 8202 8508 8208 8560
rect 8260 8548 8266 8560
rect 9217 8551 9275 8557
rect 8260 8520 8432 8548
rect 8260 8508 8266 8520
rect 7469 8483 7527 8489
rect 7469 8480 7481 8483
rect 7432 8452 7481 8480
rect 7432 8440 7438 8452
rect 7469 8449 7481 8452
rect 7515 8449 7527 8483
rect 7742 8480 7748 8492
rect 7703 8452 7748 8480
rect 7469 8443 7527 8449
rect 7742 8440 7748 8452
rect 7800 8440 7806 8492
rect 7926 8480 7932 8492
rect 7839 8452 7932 8480
rect 7926 8440 7932 8452
rect 7984 8480 7990 8492
rect 8297 8483 8355 8489
rect 8297 8480 8309 8483
rect 7984 8452 8309 8480
rect 7984 8440 7990 8452
rect 8297 8449 8309 8452
rect 8343 8449 8355 8483
rect 8297 8443 8355 8449
rect 6457 8415 6515 8421
rect 6457 8412 6469 8415
rect 6196 8384 6469 8412
rect 6457 8381 6469 8384
rect 6503 8412 6515 8415
rect 6730 8412 6736 8424
rect 6503 8384 6736 8412
rect 6503 8381 6515 8384
rect 6457 8375 6515 8381
rect 6730 8372 6736 8384
rect 6788 8412 6794 8424
rect 6917 8415 6975 8421
rect 6917 8412 6929 8415
rect 6788 8384 6929 8412
rect 6788 8372 6794 8384
rect 6917 8381 6929 8384
rect 6963 8381 6975 8415
rect 7558 8412 7564 8424
rect 7519 8384 7564 8412
rect 6917 8375 6975 8381
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 7650 8372 7656 8424
rect 7708 8412 7714 8424
rect 7708 8384 7753 8412
rect 7708 8372 7714 8384
rect 7834 8372 7840 8424
rect 7892 8412 7898 8424
rect 8021 8415 8079 8421
rect 8021 8412 8033 8415
rect 7892 8384 8033 8412
rect 7892 8372 7898 8384
rect 8021 8381 8033 8384
rect 8067 8381 8079 8415
rect 8404 8412 8432 8520
rect 9217 8517 9229 8551
rect 9263 8548 9275 8551
rect 9398 8548 9404 8560
rect 9263 8520 9404 8548
rect 9263 8517 9275 8520
rect 9217 8511 9275 8517
rect 9398 8508 9404 8520
rect 9456 8508 9462 8560
rect 9674 8548 9680 8560
rect 9600 8520 9680 8548
rect 8846 8440 8852 8492
rect 8904 8480 8910 8492
rect 9600 8489 9628 8520
rect 9674 8508 9680 8520
rect 9732 8508 9738 8560
rect 10962 8508 10968 8560
rect 11020 8548 11026 8560
rect 13265 8551 13323 8557
rect 13265 8548 13277 8551
rect 11020 8520 11468 8548
rect 11020 8508 11026 8520
rect 9585 8483 9643 8489
rect 8904 8452 9536 8480
rect 8904 8440 8910 8452
rect 9508 8424 9536 8452
rect 9585 8449 9597 8483
rect 9631 8449 9643 8483
rect 11238 8480 11244 8492
rect 11199 8452 11244 8480
rect 9585 8443 9643 8449
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11440 8489 11468 8520
rect 12820 8520 13277 8548
rect 11425 8483 11483 8489
rect 11425 8449 11437 8483
rect 11471 8449 11483 8483
rect 11425 8443 11483 8449
rect 9401 8415 9459 8421
rect 9401 8412 9413 8415
rect 8404 8384 9413 8412
rect 8021 8375 8079 8381
rect 9401 8381 9413 8384
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 9490 8372 9496 8424
rect 9548 8412 9554 8424
rect 9674 8421 9680 8424
rect 9548 8384 9593 8412
rect 9548 8372 9554 8384
rect 9670 8375 9680 8421
rect 9732 8412 9738 8424
rect 10226 8412 10232 8424
rect 9732 8384 10232 8412
rect 9674 8372 9680 8375
rect 9732 8372 9738 8384
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 12820 8421 12848 8520
rect 13265 8517 13277 8520
rect 13311 8517 13323 8551
rect 15562 8548 15568 8560
rect 13265 8511 13323 8517
rect 13648 8520 15568 8548
rect 13078 8480 13084 8492
rect 13039 8452 13084 8480
rect 13078 8440 13084 8452
rect 13136 8440 13142 8492
rect 13648 8480 13676 8520
rect 15562 8508 15568 8520
rect 15620 8508 15626 8560
rect 16574 8480 16580 8492
rect 13188 8452 13676 8480
rect 13740 8452 16580 8480
rect 12805 8415 12863 8421
rect 11348 8384 12434 8412
rect 3016 8316 3648 8344
rect 3804 8316 5488 8344
rect 3016 8304 3022 8316
rect 2225 8279 2283 8285
rect 2225 8245 2237 8279
rect 2271 8276 2283 8279
rect 2314 8276 2320 8288
rect 2271 8248 2320 8276
rect 2271 8245 2283 8248
rect 2225 8239 2283 8245
rect 2314 8236 2320 8248
rect 2372 8236 2378 8288
rect 3620 8285 3648 8316
rect 5810 8304 5816 8356
rect 5868 8344 5874 8356
rect 6273 8347 6331 8353
rect 6273 8344 6285 8347
rect 5868 8316 6285 8344
rect 5868 8304 5874 8316
rect 6273 8313 6285 8316
rect 6319 8313 6331 8347
rect 6273 8307 6331 8313
rect 6641 8347 6699 8353
rect 6641 8313 6653 8347
rect 6687 8313 6699 8347
rect 6641 8307 6699 8313
rect 6825 8347 6883 8353
rect 6825 8313 6837 8347
rect 6871 8344 6883 8347
rect 7576 8344 7604 8372
rect 6871 8316 7604 8344
rect 8297 8347 8355 8353
rect 6871 8313 6883 8316
rect 6825 8307 6883 8313
rect 8297 8313 8309 8347
rect 8343 8344 8355 8347
rect 10502 8344 10508 8356
rect 8343 8316 10508 8344
rect 8343 8313 8355 8316
rect 8297 8307 8355 8313
rect 3605 8279 3663 8285
rect 3605 8245 3617 8279
rect 3651 8245 3663 8279
rect 4154 8276 4160 8288
rect 4115 8248 4160 8276
rect 3605 8239 3663 8245
rect 4154 8236 4160 8248
rect 4212 8236 4218 8288
rect 4525 8279 4583 8285
rect 4525 8245 4537 8279
rect 4571 8276 4583 8279
rect 4614 8276 4620 8288
rect 4571 8248 4620 8276
rect 4571 8245 4583 8248
rect 4525 8239 4583 8245
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 6178 8236 6184 8288
rect 6236 8276 6242 8288
rect 6656 8276 6684 8307
rect 10502 8304 10508 8316
rect 10560 8304 10566 8356
rect 11348 8353 11376 8384
rect 11333 8347 11391 8353
rect 11333 8313 11345 8347
rect 11379 8313 11391 8347
rect 12406 8344 12434 8384
rect 12805 8381 12817 8415
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 12897 8415 12955 8421
rect 12897 8381 12909 8415
rect 12943 8412 12955 8415
rect 13188 8412 13216 8452
rect 12943 8384 13216 8412
rect 12943 8381 12955 8384
rect 12897 8375 12955 8381
rect 13262 8372 13268 8424
rect 13320 8412 13326 8424
rect 13449 8415 13507 8421
rect 13449 8412 13461 8415
rect 13320 8384 13461 8412
rect 13320 8372 13326 8384
rect 13449 8381 13461 8384
rect 13495 8381 13507 8415
rect 13449 8375 13507 8381
rect 13740 8344 13768 8452
rect 16574 8440 16580 8452
rect 16632 8440 16638 8492
rect 13906 8412 13912 8424
rect 13867 8384 13912 8412
rect 13906 8372 13912 8384
rect 13964 8372 13970 8424
rect 16114 8412 16120 8424
rect 16075 8384 16120 8412
rect 16114 8372 16120 8384
rect 16172 8372 16178 8424
rect 14090 8344 14096 8356
rect 12406 8316 13768 8344
rect 14051 8316 14096 8344
rect 11333 8307 11391 8313
rect 14090 8304 14096 8316
rect 14148 8304 14154 8356
rect 15930 8344 15936 8356
rect 15891 8316 15936 8344
rect 15930 8304 15936 8316
rect 15988 8304 15994 8356
rect 6236 8248 6684 8276
rect 6236 8236 6242 8248
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 9674 8276 9680 8288
rect 8812 8248 9680 8276
rect 8812 8236 8818 8248
rect 9674 8236 9680 8248
rect 9732 8236 9738 8288
rect 10686 8236 10692 8288
rect 10744 8276 10750 8288
rect 12437 8279 12495 8285
rect 12437 8276 12449 8279
rect 10744 8248 12449 8276
rect 10744 8236 10750 8248
rect 12437 8245 12449 8248
rect 12483 8245 12495 8279
rect 12437 8239 12495 8245
rect 1104 8186 17296 8208
rect 1104 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 6571 8186
rect 6623 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 11904 8186
rect 11956 8134 11968 8186
rect 12020 8134 17296 8186
rect 1104 8112 17296 8134
rect 6086 8032 6092 8084
rect 6144 8072 6150 8084
rect 7193 8075 7251 8081
rect 7193 8072 7205 8075
rect 6144 8044 7205 8072
rect 6144 8032 6150 8044
rect 7193 8041 7205 8044
rect 7239 8041 7251 8075
rect 7193 8035 7251 8041
rect 7561 8075 7619 8081
rect 7561 8041 7573 8075
rect 7607 8072 7619 8075
rect 12526 8072 12532 8084
rect 7607 8044 12532 8072
rect 7607 8041 7619 8044
rect 7561 8035 7619 8041
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 15933 8075 15991 8081
rect 15933 8041 15945 8075
rect 15979 8041 15991 8075
rect 15933 8035 15991 8041
rect 1857 8007 1915 8013
rect 1857 7973 1869 8007
rect 1903 8004 1915 8007
rect 2314 8004 2320 8016
rect 1903 7976 2320 8004
rect 1903 7973 1915 7976
rect 1857 7967 1915 7973
rect 2314 7964 2320 7976
rect 2372 7964 2378 8016
rect 5626 7964 5632 8016
rect 5684 8004 5690 8016
rect 5813 8007 5871 8013
rect 5813 8004 5825 8007
rect 5684 7976 5825 8004
rect 5684 7964 5690 7976
rect 5813 7973 5825 7976
rect 5859 7973 5871 8007
rect 5813 7967 5871 7973
rect 5997 8007 6055 8013
rect 5997 7973 6009 8007
rect 6043 8004 6055 8007
rect 6730 8004 6736 8016
rect 6043 7976 6736 8004
rect 6043 7973 6055 7976
rect 5997 7967 6055 7973
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1486 7936 1492 7948
rect 1443 7908 1492 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1486 7896 1492 7908
rect 1544 7896 1550 7948
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7936 2007 7939
rect 2498 7936 2504 7948
rect 1995 7908 2504 7936
rect 1995 7905 2007 7908
rect 1949 7899 2007 7905
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 5534 7896 5540 7948
rect 5592 7936 5598 7948
rect 6656 7945 6684 7976
rect 6730 7964 6736 7976
rect 6788 7964 6794 8016
rect 7653 8007 7711 8013
rect 7653 8004 7665 8007
rect 6932 7976 7665 8004
rect 6932 7945 6960 7976
rect 7653 7973 7665 7976
rect 7699 7973 7711 8007
rect 7653 7967 7711 7973
rect 15105 8007 15163 8013
rect 15105 7973 15117 8007
rect 15151 8004 15163 8007
rect 15749 8007 15807 8013
rect 15749 8004 15761 8007
rect 15151 7976 15761 8004
rect 15151 7973 15163 7976
rect 15105 7967 15163 7973
rect 15749 7973 15761 7976
rect 15795 8004 15807 8007
rect 15948 8004 15976 8035
rect 15795 7976 15976 8004
rect 15795 7973 15807 7976
rect 15749 7967 15807 7973
rect 6641 7939 6699 7945
rect 5592 7908 5856 7936
rect 5592 7896 5598 7908
rect 5166 7828 5172 7880
rect 5224 7868 5230 7880
rect 5721 7871 5779 7877
rect 5721 7868 5733 7871
rect 5224 7840 5733 7868
rect 5224 7828 5230 7840
rect 5721 7837 5733 7840
rect 5767 7837 5779 7871
rect 5828 7868 5856 7908
rect 6641 7905 6653 7939
rect 6687 7905 6699 7939
rect 6641 7899 6699 7905
rect 6917 7939 6975 7945
rect 6917 7905 6929 7939
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 7193 7939 7251 7945
rect 7193 7905 7205 7939
rect 7239 7936 7251 7939
rect 7285 7939 7343 7945
rect 7285 7936 7297 7939
rect 7239 7908 7297 7936
rect 7239 7905 7251 7908
rect 7193 7899 7251 7905
rect 7285 7905 7297 7908
rect 7331 7905 7343 7939
rect 7285 7899 7343 7905
rect 7374 7896 7380 7948
rect 7432 7936 7438 7948
rect 7926 7936 7932 7948
rect 7432 7908 7477 7936
rect 7576 7908 7932 7936
rect 7432 7896 7438 7908
rect 5902 7868 5908 7880
rect 5815 7840 5908 7868
rect 5721 7831 5779 7837
rect 5736 7800 5764 7831
rect 5902 7828 5908 7840
rect 5960 7868 5966 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 5960 7840 6745 7868
rect 5960 7828 5966 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 7576 7877 7604 7908
rect 7926 7896 7932 7908
rect 7984 7896 7990 7948
rect 9950 7936 9956 7948
rect 9911 7908 9956 7936
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 15289 7939 15347 7945
rect 15289 7936 15301 7939
rect 12406 7908 15301 7936
rect 7561 7871 7619 7877
rect 6880 7840 6925 7868
rect 6880 7828 6886 7840
rect 7561 7837 7573 7871
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 8110 7828 8116 7880
rect 8168 7868 8174 7880
rect 9309 7871 9367 7877
rect 9309 7868 9321 7871
rect 8168 7840 9321 7868
rect 8168 7828 8174 7840
rect 9309 7837 9321 7840
rect 9355 7837 9367 7871
rect 9309 7831 9367 7837
rect 6178 7800 6184 7812
rect 5736 7772 6184 7800
rect 6178 7760 6184 7772
rect 6236 7760 6242 7812
rect 6273 7803 6331 7809
rect 6273 7769 6285 7803
rect 6319 7800 6331 7803
rect 12406 7800 12434 7908
rect 15289 7905 15301 7908
rect 15335 7905 15347 7939
rect 15838 7936 15844 7948
rect 15799 7908 15844 7936
rect 15289 7899 15347 7905
rect 15304 7868 15332 7899
rect 15838 7896 15844 7908
rect 15896 7896 15902 7948
rect 15930 7896 15936 7948
rect 15988 7936 15994 7948
rect 15988 7908 16033 7936
rect 15988 7896 15994 7908
rect 16301 7871 16359 7877
rect 16301 7868 16313 7871
rect 15304 7840 16313 7868
rect 16301 7837 16313 7840
rect 16347 7837 16359 7871
rect 16301 7831 16359 7837
rect 14918 7800 14924 7812
rect 6319 7772 12434 7800
rect 14879 7772 14924 7800
rect 6319 7769 6331 7772
rect 6273 7763 6331 7769
rect 14918 7760 14924 7772
rect 14976 7760 14982 7812
rect 6457 7735 6515 7741
rect 6457 7701 6469 7735
rect 6503 7732 6515 7735
rect 6914 7732 6920 7744
rect 6503 7704 6920 7732
rect 6503 7701 6515 7704
rect 6457 7695 6515 7701
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 7653 7735 7711 7741
rect 7653 7701 7665 7735
rect 7699 7732 7711 7735
rect 7837 7735 7895 7741
rect 7837 7732 7849 7735
rect 7699 7704 7849 7732
rect 7699 7701 7711 7704
rect 7653 7695 7711 7701
rect 7837 7701 7849 7704
rect 7883 7732 7895 7735
rect 8294 7732 8300 7744
rect 7883 7704 8300 7732
rect 7883 7701 7895 7704
rect 7837 7695 7895 7701
rect 8294 7692 8300 7704
rect 8352 7692 8358 7744
rect 1104 7642 17296 7664
rect 1104 7590 3680 7642
rect 3732 7590 3744 7642
rect 3796 7590 3808 7642
rect 3860 7590 3872 7642
rect 3924 7590 9078 7642
rect 9130 7590 9142 7642
rect 9194 7590 9206 7642
rect 9258 7590 9270 7642
rect 9322 7590 14475 7642
rect 14527 7590 14539 7642
rect 14591 7590 14603 7642
rect 14655 7590 14667 7642
rect 14719 7590 17296 7642
rect 1104 7568 17296 7590
rect 2498 7528 2504 7540
rect 2459 7500 2504 7528
rect 2498 7488 2504 7500
rect 2556 7488 2562 7540
rect 8205 7531 8263 7537
rect 8205 7497 8217 7531
rect 8251 7528 8263 7531
rect 8846 7528 8852 7540
rect 8251 7500 8852 7528
rect 8251 7497 8263 7500
rect 8205 7491 8263 7497
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 8941 7531 8999 7537
rect 8941 7497 8953 7531
rect 8987 7528 8999 7531
rect 10594 7528 10600 7540
rect 8987 7500 10600 7528
rect 8987 7497 8999 7500
rect 8941 7491 8999 7497
rect 1946 7420 1952 7472
rect 2004 7460 2010 7472
rect 2004 7432 5304 7460
rect 2004 7420 2010 7432
rect 3881 7395 3939 7401
rect 3881 7361 3893 7395
rect 3927 7392 3939 7395
rect 4154 7392 4160 7404
rect 3927 7364 4160 7392
rect 3927 7361 3939 7364
rect 3881 7355 3939 7361
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 4249 7327 4307 7333
rect 4249 7293 4261 7327
rect 4295 7324 4307 7327
rect 5074 7324 5080 7336
rect 4295 7296 5080 7324
rect 4295 7293 4307 7296
rect 4249 7287 4307 7293
rect 5074 7284 5080 7296
rect 5132 7284 5138 7336
rect 2498 7216 2504 7268
rect 2556 7256 2562 7268
rect 2593 7259 2651 7265
rect 2593 7256 2605 7259
rect 2556 7228 2605 7256
rect 2556 7216 2562 7228
rect 2593 7225 2605 7228
rect 2639 7225 2651 7259
rect 4341 7259 4399 7265
rect 4341 7256 4353 7259
rect 2593 7219 2651 7225
rect 4264 7228 4353 7256
rect 4264 7197 4292 7228
rect 4341 7225 4353 7228
rect 4387 7256 4399 7259
rect 4982 7256 4988 7268
rect 4387 7228 4988 7256
rect 4387 7225 4399 7228
rect 4341 7219 4399 7225
rect 4982 7216 4988 7228
rect 5040 7216 5046 7268
rect 5169 7259 5227 7265
rect 5169 7225 5181 7259
rect 5215 7225 5227 7259
rect 5276 7256 5304 7432
rect 6086 7420 6092 7472
rect 6144 7460 6150 7472
rect 6549 7463 6607 7469
rect 6549 7460 6561 7463
rect 6144 7432 6561 7460
rect 6144 7420 6150 7432
rect 6549 7429 6561 7432
rect 6595 7429 6607 7463
rect 6549 7423 6607 7429
rect 7834 7420 7840 7472
rect 7892 7460 7898 7472
rect 8956 7460 8984 7491
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 7892 7432 8984 7460
rect 10321 7463 10379 7469
rect 7892 7420 7898 7432
rect 8220 7404 8248 7432
rect 10321 7429 10333 7463
rect 10367 7460 10379 7463
rect 11330 7460 11336 7472
rect 10367 7432 11336 7460
rect 10367 7429 10379 7432
rect 10321 7423 10379 7429
rect 11330 7420 11336 7432
rect 11388 7420 11394 7472
rect 14090 7420 14096 7472
rect 14148 7460 14154 7472
rect 14185 7463 14243 7469
rect 14185 7460 14197 7463
rect 14148 7432 14197 7460
rect 14148 7420 14154 7432
rect 14185 7429 14197 7432
rect 14231 7429 14243 7463
rect 14185 7423 14243 7429
rect 6914 7392 6920 7404
rect 6875 7364 6920 7392
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 7650 7352 7656 7404
rect 7708 7392 7714 7404
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 7708 7364 7941 7392
rect 7708 7352 7714 7364
rect 7929 7361 7941 7364
rect 7975 7392 7987 7395
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 7975 7364 8125 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 8113 7361 8125 7364
rect 8159 7361 8171 7395
rect 8113 7355 8171 7361
rect 8202 7352 8208 7404
rect 8260 7352 8266 7404
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 9861 7395 9919 7401
rect 9861 7392 9873 7395
rect 8352 7364 9873 7392
rect 8352 7352 8358 7364
rect 9861 7361 9873 7364
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 13262 7392 13268 7404
rect 10652 7364 12480 7392
rect 13175 7364 13268 7392
rect 10652 7352 10658 7364
rect 6178 7284 6184 7336
rect 6236 7324 6242 7336
rect 7101 7327 7159 7333
rect 7101 7324 7113 7327
rect 6236 7296 7113 7324
rect 6236 7284 6242 7296
rect 7101 7293 7113 7296
rect 7147 7324 7159 7327
rect 7374 7324 7380 7336
rect 7147 7296 7380 7324
rect 7147 7293 7159 7296
rect 7101 7287 7159 7293
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 8018 7324 8024 7336
rect 7979 7296 8024 7324
rect 8018 7284 8024 7296
rect 8076 7284 8082 7336
rect 8386 7324 8392 7336
rect 8347 7296 8392 7324
rect 8386 7284 8392 7296
rect 8444 7284 8450 7336
rect 10873 7327 10931 7333
rect 8680 7296 10088 7324
rect 7009 7259 7067 7265
rect 7009 7256 7021 7259
rect 5276 7228 7021 7256
rect 5169 7219 5227 7225
rect 7009 7225 7021 7228
rect 7055 7225 7067 7259
rect 8680 7256 8708 7296
rect 7009 7219 7067 7225
rect 8220 7228 8708 7256
rect 4249 7191 4307 7197
rect 4249 7157 4261 7191
rect 4295 7157 4307 7191
rect 4249 7151 4307 7157
rect 4430 7148 4436 7200
rect 4488 7188 4494 7200
rect 4488 7160 4533 7188
rect 4488 7148 4494 7160
rect 4890 7148 4896 7200
rect 4948 7188 4954 7200
rect 5077 7191 5135 7197
rect 5077 7188 5089 7191
rect 4948 7160 5089 7188
rect 4948 7148 4954 7160
rect 5077 7157 5089 7160
rect 5123 7157 5135 7191
rect 5184 7188 5212 7219
rect 8220 7188 8248 7228
rect 8754 7216 8760 7268
rect 8812 7256 8818 7268
rect 8812 7228 8857 7256
rect 8812 7216 8818 7228
rect 8938 7216 8944 7268
rect 8996 7265 9002 7268
rect 8996 7259 9020 7265
rect 9008 7225 9020 7259
rect 8996 7219 9020 7225
rect 9769 7259 9827 7265
rect 9769 7225 9781 7259
rect 9815 7225 9827 7259
rect 9769 7219 9827 7225
rect 8996 7216 9002 7219
rect 5184 7160 8248 7188
rect 5077 7151 5135 7157
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 8573 7191 8631 7197
rect 8573 7188 8585 7191
rect 8352 7160 8585 7188
rect 8352 7148 8358 7160
rect 8573 7157 8585 7160
rect 8619 7157 8631 7191
rect 8573 7151 8631 7157
rect 8846 7148 8852 7200
rect 8904 7188 8910 7200
rect 9125 7191 9183 7197
rect 9125 7188 9137 7191
rect 8904 7160 9137 7188
rect 8904 7148 8910 7160
rect 9125 7157 9137 7160
rect 9171 7188 9183 7191
rect 9582 7188 9588 7200
rect 9171 7160 9588 7188
rect 9171 7157 9183 7160
rect 9125 7151 9183 7157
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 9784 7188 9812 7219
rect 9858 7216 9864 7268
rect 9916 7256 9922 7268
rect 10060 7256 10088 7296
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 11054 7324 11060 7336
rect 10919 7296 11060 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 11425 7327 11483 7333
rect 11425 7293 11437 7327
rect 11471 7324 11483 7327
rect 12066 7324 12072 7336
rect 11471 7296 12072 7324
rect 11471 7293 11483 7296
rect 11425 7287 11483 7293
rect 12066 7284 12072 7296
rect 12124 7284 12130 7336
rect 12452 7333 12480 7364
rect 12437 7327 12495 7333
rect 12437 7293 12449 7327
rect 12483 7293 12495 7327
rect 12618 7324 12624 7336
rect 12579 7296 12624 7324
rect 12437 7287 12495 7293
rect 12618 7284 12624 7296
rect 12676 7284 12682 7336
rect 13188 7333 13216 7364
rect 13262 7352 13268 7364
rect 13320 7392 13326 7404
rect 13817 7395 13875 7401
rect 13817 7392 13829 7395
rect 13320 7364 13829 7392
rect 13320 7352 13326 7364
rect 13817 7361 13829 7364
rect 13863 7361 13875 7395
rect 13817 7355 13875 7361
rect 13173 7327 13231 7333
rect 13173 7293 13185 7327
rect 13219 7293 13231 7327
rect 13173 7287 13231 7293
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7324 13783 7327
rect 13998 7324 14004 7336
rect 13771 7296 14004 7324
rect 13771 7293 13783 7296
rect 13725 7287 13783 7293
rect 13998 7284 14004 7296
rect 14056 7324 14062 7336
rect 14918 7324 14924 7336
rect 14056 7296 14924 7324
rect 14056 7284 14062 7296
rect 14918 7284 14924 7296
rect 14976 7284 14982 7336
rect 10962 7256 10968 7268
rect 9916 7228 9961 7256
rect 10060 7228 10968 7256
rect 9916 7216 9922 7228
rect 10962 7216 10968 7228
rect 11020 7216 11026 7268
rect 13633 7259 13691 7265
rect 13633 7225 13645 7259
rect 13679 7225 13691 7259
rect 13633 7219 13691 7225
rect 9950 7188 9956 7200
rect 9784 7160 9956 7188
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 12802 7188 12808 7200
rect 12763 7160 12808 7188
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 13538 7148 13544 7200
rect 13596 7188 13602 7200
rect 13648 7188 13676 7219
rect 14185 7191 14243 7197
rect 14185 7188 14197 7191
rect 13596 7160 14197 7188
rect 13596 7148 13602 7160
rect 14185 7157 14197 7160
rect 14231 7157 14243 7191
rect 14185 7151 14243 7157
rect 1104 7098 17296 7120
rect 1104 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 6571 7098
rect 6623 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 11904 7098
rect 11956 7046 11968 7098
rect 12020 7046 17296 7098
rect 1104 7024 17296 7046
rect 1949 6987 2007 6993
rect 1949 6953 1961 6987
rect 1995 6984 2007 6987
rect 5445 6987 5503 6993
rect 5445 6984 5457 6987
rect 1995 6956 5457 6984
rect 1995 6953 2007 6956
rect 1949 6947 2007 6953
rect 5445 6953 5457 6956
rect 5491 6953 5503 6987
rect 8294 6984 8300 6996
rect 8255 6956 8300 6984
rect 5445 6947 5503 6953
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 10778 6984 10784 6996
rect 10336 6956 10784 6984
rect 4430 6916 4436 6928
rect 4391 6888 4436 6916
rect 4430 6876 4436 6888
rect 4488 6876 4494 6928
rect 4982 6916 4988 6928
rect 4943 6888 4988 6916
rect 4982 6876 4988 6888
rect 5040 6876 5046 6928
rect 8478 6876 8484 6928
rect 8536 6916 8542 6928
rect 8536 6888 9444 6916
rect 8536 6876 8542 6888
rect 1578 6808 1584 6860
rect 1636 6848 1642 6860
rect 1857 6851 1915 6857
rect 1857 6848 1869 6851
rect 1636 6820 1869 6848
rect 1636 6808 1642 6820
rect 1857 6817 1869 6820
rect 1903 6817 1915 6851
rect 1857 6811 1915 6817
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 3970 6848 3976 6860
rect 3927 6820 3976 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 3970 6808 3976 6820
rect 4028 6808 4034 6860
rect 4154 6808 4160 6860
rect 4212 6848 4218 6860
rect 4525 6851 4583 6857
rect 4525 6848 4537 6851
rect 4212 6820 4537 6848
rect 4212 6808 4218 6820
rect 4525 6817 4537 6820
rect 4571 6817 4583 6851
rect 4525 6811 4583 6817
rect 4890 6808 4896 6860
rect 4948 6848 4954 6860
rect 5077 6851 5135 6857
rect 5077 6848 5089 6851
rect 4948 6820 5089 6848
rect 4948 6808 4954 6820
rect 5077 6817 5089 6820
rect 5123 6848 5135 6851
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 5123 6820 5365 6848
rect 5123 6817 5135 6820
rect 5077 6811 5135 6817
rect 5353 6817 5365 6820
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6848 5687 6851
rect 6270 6848 6276 6860
rect 5675 6820 6276 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 6270 6808 6276 6820
rect 6328 6848 6334 6860
rect 7466 6848 7472 6860
rect 6328 6820 7472 6848
rect 6328 6808 6334 6820
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 7650 6848 7656 6860
rect 7611 6820 7656 6848
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 7745 6851 7803 6857
rect 7745 6817 7757 6851
rect 7791 6848 7803 6851
rect 7834 6848 7840 6860
rect 7791 6820 7840 6848
rect 7791 6817 7803 6820
rect 7745 6811 7803 6817
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 8938 6808 8944 6860
rect 8996 6848 9002 6860
rect 9416 6857 9444 6888
rect 10336 6857 10364 6956
rect 10778 6944 10784 6956
rect 10836 6984 10842 6996
rect 10873 6987 10931 6993
rect 10873 6984 10885 6987
rect 10836 6956 10885 6984
rect 10836 6944 10842 6956
rect 10873 6953 10885 6956
rect 10919 6953 10931 6987
rect 10873 6947 10931 6953
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 13633 6987 13691 6993
rect 13633 6984 13645 6987
rect 12860 6956 13645 6984
rect 12860 6944 12866 6956
rect 13633 6953 13645 6956
rect 13679 6953 13691 6987
rect 13633 6947 13691 6953
rect 15838 6944 15844 6996
rect 15896 6984 15902 6996
rect 16393 6987 16451 6993
rect 16393 6984 16405 6987
rect 15896 6956 16405 6984
rect 15896 6944 15902 6956
rect 16393 6953 16405 6956
rect 16439 6953 16451 6987
rect 16393 6947 16451 6953
rect 10962 6876 10968 6928
rect 11020 6916 11026 6928
rect 12526 6916 12532 6928
rect 11020 6888 11284 6916
rect 12487 6888 12532 6916
rect 11020 6876 11026 6888
rect 9217 6851 9275 6857
rect 9217 6848 9229 6851
rect 8996 6820 9229 6848
rect 8996 6808 9002 6820
rect 9217 6817 9229 6820
rect 9263 6817 9275 6851
rect 9217 6811 9275 6817
rect 9401 6851 9459 6857
rect 9401 6817 9413 6851
rect 9447 6817 9459 6851
rect 9401 6811 9459 6817
rect 9861 6851 9919 6857
rect 9861 6817 9873 6851
rect 9907 6817 9919 6851
rect 9861 6811 9919 6817
rect 10321 6851 10379 6857
rect 10321 6817 10333 6851
rect 10367 6817 10379 6851
rect 10321 6811 10379 6817
rect 10413 6851 10471 6857
rect 10413 6817 10425 6851
rect 10459 6848 10471 6851
rect 11146 6848 11152 6860
rect 10459 6820 10640 6848
rect 11107 6820 11152 6848
rect 10459 6817 10471 6820
rect 10413 6811 10471 6817
rect 1670 6780 1676 6792
rect 1631 6752 1676 6780
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 5718 6740 5724 6792
rect 5776 6780 5782 6792
rect 5905 6783 5963 6789
rect 5905 6780 5917 6783
rect 5776 6752 5917 6780
rect 5776 6740 5782 6752
rect 5905 6749 5917 6752
rect 5951 6749 5963 6783
rect 8018 6780 8024 6792
rect 7979 6752 8024 6780
rect 5905 6743 5963 6749
rect 2498 6672 2504 6724
rect 2556 6712 2562 6724
rect 4341 6715 4399 6721
rect 4341 6712 4353 6715
rect 2556 6684 4353 6712
rect 2556 6672 2562 6684
rect 4341 6681 4353 6684
rect 4387 6681 4399 6715
rect 4341 6675 4399 6681
rect 5074 6672 5080 6724
rect 5132 6712 5138 6724
rect 5169 6715 5227 6721
rect 5169 6712 5181 6715
rect 5132 6684 5181 6712
rect 5132 6672 5138 6684
rect 5169 6681 5181 6684
rect 5215 6681 5227 6715
rect 5920 6712 5948 6743
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6780 8263 6783
rect 8386 6780 8392 6792
rect 8251 6752 8392 6780
rect 8251 6749 8263 6752
rect 8205 6743 8263 6749
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8496 6752 9137 6780
rect 6822 6712 6828 6724
rect 5920 6684 6828 6712
rect 5169 6675 5227 6681
rect 6822 6672 6828 6684
rect 6880 6712 6886 6724
rect 8496 6712 8524 6752
rect 9125 6749 9137 6752
rect 9171 6780 9183 6783
rect 9490 6780 9496 6792
rect 9171 6752 9496 6780
rect 9171 6749 9183 6752
rect 9125 6743 9183 6749
rect 9490 6740 9496 6752
rect 9548 6740 9554 6792
rect 9876 6780 9904 6811
rect 10505 6783 10563 6789
rect 10505 6780 10517 6783
rect 9876 6752 10517 6780
rect 6880 6684 8524 6712
rect 8665 6715 8723 6721
rect 6880 6672 6886 6684
rect 8665 6681 8677 6715
rect 8711 6712 8723 6715
rect 9876 6712 9904 6752
rect 10505 6749 10517 6752
rect 10551 6749 10563 6783
rect 10612 6780 10640 6820
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 11256 6848 11284 6888
rect 12526 6876 12532 6888
rect 12584 6876 12590 6928
rect 12713 6919 12771 6925
rect 12713 6885 12725 6919
rect 12759 6885 12771 6919
rect 12713 6879 12771 6885
rect 13725 6919 13783 6925
rect 13725 6885 13737 6919
rect 13771 6916 13783 6919
rect 13771 6888 13952 6916
rect 13771 6885 13783 6888
rect 13725 6879 13783 6885
rect 11333 6851 11391 6857
rect 11333 6848 11345 6851
rect 11256 6820 11345 6848
rect 11333 6817 11345 6820
rect 11379 6817 11391 6851
rect 12066 6848 12072 6860
rect 12027 6820 12072 6848
rect 11333 6811 11391 6817
rect 12066 6808 12072 6820
rect 12124 6808 12130 6860
rect 12728 6848 12756 6879
rect 12452 6820 12756 6848
rect 11164 6780 11192 6808
rect 10612 6752 11192 6780
rect 10505 6743 10563 6749
rect 10870 6712 10876 6724
rect 8711 6684 9904 6712
rect 10831 6684 10876 6712
rect 8711 6681 8723 6684
rect 8665 6675 8723 6681
rect 10870 6672 10876 6684
rect 10928 6672 10934 6724
rect 12084 6712 12112 6808
rect 12253 6715 12311 6721
rect 12253 6712 12265 6715
rect 12084 6684 12265 6712
rect 12253 6681 12265 6684
rect 12299 6681 12311 6715
rect 12253 6675 12311 6681
rect 2317 6647 2375 6653
rect 2317 6613 2329 6647
rect 2363 6644 2375 6647
rect 2406 6644 2412 6656
rect 2363 6616 2412 6644
rect 2363 6613 2375 6616
rect 2317 6607 2375 6613
rect 2406 6604 2412 6616
rect 2464 6604 2470 6656
rect 5813 6647 5871 6653
rect 5813 6613 5825 6647
rect 5859 6644 5871 6647
rect 5994 6644 6000 6656
rect 5859 6616 6000 6644
rect 5859 6613 5871 6616
rect 5813 6607 5871 6613
rect 5994 6604 6000 6616
rect 6052 6604 6058 6656
rect 7282 6644 7288 6656
rect 7243 6616 7288 6644
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 8018 6644 8024 6656
rect 7432 6616 8024 6644
rect 7432 6604 7438 6616
rect 8018 6604 8024 6616
rect 8076 6604 8082 6656
rect 9582 6644 9588 6656
rect 9543 6616 9588 6644
rect 9582 6604 9588 6616
rect 9640 6604 9646 6656
rect 12452 6644 12480 6820
rect 12526 6740 12532 6792
rect 12584 6780 12590 6792
rect 12805 6783 12863 6789
rect 12805 6780 12817 6783
rect 12584 6752 12817 6780
rect 12584 6740 12590 6752
rect 12805 6749 12817 6752
rect 12851 6780 12863 6783
rect 13078 6780 13084 6792
rect 12851 6752 13084 6780
rect 12851 6749 12863 6752
rect 12805 6743 12863 6749
rect 13078 6740 13084 6752
rect 13136 6780 13142 6792
rect 13817 6783 13875 6789
rect 13817 6780 13829 6783
rect 13136 6752 13829 6780
rect 13136 6740 13142 6752
rect 13817 6749 13829 6752
rect 13863 6749 13875 6783
rect 13924 6780 13952 6888
rect 15838 6808 15844 6860
rect 15896 6848 15902 6860
rect 16301 6851 16359 6857
rect 16301 6848 16313 6851
rect 15896 6820 16313 6848
rect 15896 6808 15902 6820
rect 16301 6817 16313 6820
rect 16347 6817 16359 6851
rect 16942 6848 16948 6860
rect 16903 6820 16948 6848
rect 16301 6811 16359 6817
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 13924 6752 15240 6780
rect 13817 6743 13875 6749
rect 13262 6712 13268 6724
rect 13223 6684 13268 6712
rect 13262 6672 13268 6684
rect 13320 6672 13326 6724
rect 15212 6712 15240 6752
rect 16761 6715 16819 6721
rect 16761 6712 16773 6715
rect 15212 6684 16773 6712
rect 16761 6681 16773 6684
rect 16807 6681 16819 6715
rect 16761 6675 16819 6681
rect 16574 6644 16580 6656
rect 12452 6616 16580 6644
rect 16574 6604 16580 6616
rect 16632 6604 16638 6656
rect 1104 6554 17296 6576
rect 1104 6502 3680 6554
rect 3732 6502 3744 6554
rect 3796 6502 3808 6554
rect 3860 6502 3872 6554
rect 3924 6502 9078 6554
rect 9130 6502 9142 6554
rect 9194 6502 9206 6554
rect 9258 6502 9270 6554
rect 9322 6502 14475 6554
rect 14527 6502 14539 6554
rect 14591 6502 14603 6554
rect 14655 6502 14667 6554
rect 14719 6502 17296 6554
rect 1104 6480 17296 6502
rect 7650 6400 7656 6452
rect 7708 6440 7714 6452
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 7708 6412 7941 6440
rect 7708 6400 7714 6412
rect 7929 6409 7941 6412
rect 7975 6409 7987 6443
rect 10870 6440 10876 6452
rect 10831 6412 10876 6440
rect 7929 6403 7987 6409
rect 10870 6400 10876 6412
rect 10928 6400 10934 6452
rect 11054 6440 11060 6452
rect 11015 6412 11060 6440
rect 11054 6400 11060 6412
rect 11112 6400 11118 6452
rect 15381 6443 15439 6449
rect 15381 6409 15393 6443
rect 15427 6440 15439 6443
rect 15838 6440 15844 6452
rect 15427 6412 15844 6440
rect 15427 6409 15439 6412
rect 15381 6403 15439 6409
rect 15838 6400 15844 6412
rect 15896 6400 15902 6452
rect 5994 6372 6000 6384
rect 5907 6344 6000 6372
rect 5994 6332 6000 6344
rect 6052 6372 6058 6384
rect 6052 6344 7880 6372
rect 6052 6332 6058 6344
rect 1670 6304 1676 6316
rect 1631 6276 1676 6304
rect 1670 6264 1676 6276
rect 1728 6264 1734 6316
rect 5537 6307 5595 6313
rect 5537 6304 5549 6307
rect 1964 6276 5549 6304
rect 1964 6245 1992 6276
rect 5537 6273 5549 6276
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 1949 6239 2007 6245
rect 1949 6205 1961 6239
rect 1995 6205 2007 6239
rect 3145 6239 3203 6245
rect 3145 6236 3157 6239
rect 1949 6199 2007 6205
rect 2746 6208 3157 6236
rect 2498 6128 2504 6180
rect 2556 6168 2562 6180
rect 2746 6168 2774 6208
rect 3145 6205 3157 6208
rect 3191 6205 3203 6239
rect 3145 6199 3203 6205
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 3970 6236 3976 6248
rect 3927 6208 3976 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 5721 6239 5779 6245
rect 5721 6205 5733 6239
rect 5767 6236 5779 6239
rect 5810 6236 5816 6248
rect 5767 6208 5816 6236
rect 5767 6205 5779 6208
rect 5721 6199 5779 6205
rect 5810 6196 5816 6208
rect 5868 6196 5874 6248
rect 6012 6245 6040 6332
rect 7852 6316 7880 6344
rect 7374 6304 7380 6316
rect 7335 6276 7380 6304
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 7834 6264 7840 6316
rect 7892 6304 7898 6316
rect 8021 6307 8079 6313
rect 8021 6304 8033 6307
rect 7892 6276 8033 6304
rect 7892 6264 7898 6276
rect 8021 6273 8033 6276
rect 8067 6273 8079 6307
rect 8021 6267 8079 6273
rect 11330 6264 11336 6316
rect 11388 6304 11394 6316
rect 15473 6307 15531 6313
rect 15473 6304 15485 6307
rect 11388 6276 15485 6304
rect 11388 6264 11394 6276
rect 5997 6239 6055 6245
rect 5997 6205 6009 6239
rect 6043 6205 6055 6239
rect 5997 6199 6055 6205
rect 7193 6239 7251 6245
rect 7193 6205 7205 6239
rect 7239 6236 7251 6239
rect 7282 6236 7288 6248
rect 7239 6208 7288 6236
rect 7239 6205 7251 6208
rect 7193 6199 7251 6205
rect 7282 6196 7288 6208
rect 7340 6196 7346 6248
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 7929 6239 7987 6245
rect 7929 6236 7941 6239
rect 7524 6208 7941 6236
rect 7524 6196 7530 6208
rect 7929 6205 7941 6208
rect 7975 6236 7987 6239
rect 8754 6236 8760 6248
rect 7975 6208 8760 6236
rect 7975 6205 7987 6208
rect 7929 6199 7987 6205
rect 8754 6196 8760 6208
rect 8812 6196 8818 6248
rect 10689 6239 10747 6245
rect 10689 6205 10701 6239
rect 10735 6205 10747 6239
rect 10689 6199 10747 6205
rect 2556 6140 2774 6168
rect 2961 6171 3019 6177
rect 2556 6128 2562 6140
rect 2961 6137 2973 6171
rect 3007 6168 3019 6171
rect 4890 6168 4896 6180
rect 3007 6140 4896 6168
rect 3007 6137 3019 6140
rect 2961 6131 3019 6137
rect 4890 6128 4896 6140
rect 4948 6128 4954 6180
rect 5902 6168 5908 6180
rect 5863 6140 5908 6168
rect 5902 6128 5908 6140
rect 5960 6128 5966 6180
rect 10704 6168 10732 6199
rect 10778 6196 10784 6248
rect 10836 6236 10842 6248
rect 10965 6239 11023 6245
rect 10965 6236 10977 6239
rect 10836 6208 10977 6236
rect 10836 6196 10842 6208
rect 10965 6205 10977 6208
rect 11011 6205 11023 6239
rect 13538 6236 13544 6248
rect 13499 6208 13544 6236
rect 10965 6199 11023 6205
rect 13538 6196 13544 6208
rect 13596 6196 13602 6248
rect 14844 6245 14872 6276
rect 15473 6273 15485 6276
rect 15519 6273 15531 6307
rect 15473 6267 15531 6273
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 15286 6196 15292 6248
rect 15344 6236 15350 6248
rect 15381 6239 15439 6245
rect 15381 6236 15393 6239
rect 15344 6208 15393 6236
rect 15344 6196 15350 6208
rect 15381 6205 15393 6208
rect 15427 6205 15439 6239
rect 15838 6236 15844 6248
rect 15799 6208 15844 6236
rect 15381 6199 15439 6205
rect 15838 6196 15844 6208
rect 15896 6196 15902 6248
rect 11146 6168 11152 6180
rect 10704 6140 11152 6168
rect 11146 6128 11152 6140
rect 11204 6168 11210 6180
rect 13357 6171 13415 6177
rect 13357 6168 13369 6171
rect 11204 6140 13369 6168
rect 11204 6128 11210 6140
rect 13357 6137 13369 6140
rect 13403 6137 13415 6171
rect 13357 6131 13415 6137
rect 1578 6060 1584 6112
rect 1636 6100 1642 6112
rect 1857 6103 1915 6109
rect 1857 6100 1869 6103
rect 1636 6072 1869 6100
rect 1636 6060 1642 6072
rect 1857 6069 1869 6072
rect 1903 6069 1915 6103
rect 2314 6100 2320 6112
rect 2275 6072 2320 6100
rect 1857 6063 1915 6069
rect 2314 6060 2320 6072
rect 2372 6060 2378 6112
rect 6822 6100 6828 6112
rect 6783 6072 6828 6100
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 7098 6060 7104 6112
rect 7156 6100 7162 6112
rect 7285 6103 7343 6109
rect 7285 6100 7297 6103
rect 7156 6072 7297 6100
rect 7156 6060 7162 6072
rect 7285 6069 7297 6072
rect 7331 6069 7343 6103
rect 8294 6100 8300 6112
rect 8255 6072 8300 6100
rect 7285 6063 7343 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 1104 6010 17296 6032
rect 1104 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 6571 6010
rect 6623 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 11904 6010
rect 11956 5958 11968 6010
rect 12020 5958 17296 6010
rect 1104 5936 17296 5958
rect 1578 5896 1584 5908
rect 1539 5868 1584 5896
rect 1578 5856 1584 5868
rect 1636 5856 1642 5908
rect 4798 5896 4804 5908
rect 4632 5868 4804 5896
rect 4246 5828 4252 5840
rect 4207 5800 4252 5828
rect 4246 5788 4252 5800
rect 4304 5788 4310 5840
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 4632 5769 4660 5868
rect 4798 5856 4804 5868
rect 4856 5856 4862 5908
rect 12066 5896 12072 5908
rect 12027 5868 12072 5896
rect 12066 5856 12072 5868
rect 12124 5856 12130 5908
rect 15838 5896 15844 5908
rect 15799 5868 15844 5896
rect 15838 5856 15844 5868
rect 15896 5856 15902 5908
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5729 4675 5763
rect 4798 5760 4804 5772
rect 4759 5732 4804 5760
rect 4617 5723 4675 5729
rect 4798 5720 4804 5732
rect 4856 5720 4862 5772
rect 10226 5760 10232 5772
rect 10187 5732 10232 5760
rect 10226 5720 10232 5732
rect 10284 5720 10290 5772
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 15749 5763 15807 5769
rect 12492 5732 12537 5760
rect 12492 5720 12498 5732
rect 15749 5729 15761 5763
rect 15795 5760 15807 5763
rect 15838 5760 15844 5772
rect 15795 5732 15844 5760
rect 15795 5729 15807 5732
rect 15749 5723 15807 5729
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 11698 5692 11704 5704
rect 11659 5664 11704 5692
rect 11698 5652 11704 5664
rect 11756 5652 11762 5704
rect 12069 5627 12127 5633
rect 12069 5593 12081 5627
rect 12115 5624 12127 5627
rect 12253 5627 12311 5633
rect 12253 5624 12265 5627
rect 12115 5596 12265 5624
rect 12115 5593 12127 5596
rect 12069 5587 12127 5593
rect 12253 5593 12265 5596
rect 12299 5593 12311 5627
rect 12253 5587 12311 5593
rect 10134 5556 10140 5568
rect 10095 5528 10140 5556
rect 10134 5516 10140 5528
rect 10192 5516 10198 5568
rect 1104 5466 17296 5488
rect 1104 5414 3680 5466
rect 3732 5414 3744 5466
rect 3796 5414 3808 5466
rect 3860 5414 3872 5466
rect 3924 5414 9078 5466
rect 9130 5414 9142 5466
rect 9194 5414 9206 5466
rect 9258 5414 9270 5466
rect 9322 5414 14475 5466
rect 14527 5414 14539 5466
rect 14591 5414 14603 5466
rect 14655 5414 14667 5466
rect 14719 5414 17296 5466
rect 1104 5392 17296 5414
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 12529 5355 12587 5361
rect 12529 5352 12541 5355
rect 12492 5324 12541 5352
rect 12492 5312 12498 5324
rect 12529 5321 12541 5324
rect 12575 5321 12587 5355
rect 12529 5315 12587 5321
rect 12713 5355 12771 5361
rect 12713 5321 12725 5355
rect 12759 5352 12771 5355
rect 13725 5355 13783 5361
rect 13725 5352 13737 5355
rect 12759 5324 13737 5352
rect 12759 5321 12771 5324
rect 12713 5315 12771 5321
rect 13725 5321 13737 5324
rect 13771 5321 13783 5355
rect 13725 5315 13783 5321
rect 2406 5284 2412 5296
rect 1780 5256 2412 5284
rect 1780 5157 1808 5256
rect 2406 5244 2412 5256
rect 2464 5244 2470 5296
rect 2777 5287 2835 5293
rect 2777 5253 2789 5287
rect 2823 5284 2835 5287
rect 2869 5287 2927 5293
rect 2869 5284 2881 5287
rect 2823 5256 2881 5284
rect 2823 5253 2835 5256
rect 2777 5247 2835 5253
rect 2869 5253 2881 5256
rect 2915 5253 2927 5287
rect 11057 5287 11115 5293
rect 2869 5247 2927 5253
rect 10060 5256 10916 5284
rect 2332 5188 2774 5216
rect 2332 5157 2360 5188
rect 1765 5151 1823 5157
rect 1765 5117 1777 5151
rect 1811 5117 1823 5151
rect 1765 5111 1823 5117
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5117 2375 5151
rect 2317 5111 2375 5117
rect 2406 5108 2412 5160
rect 2464 5148 2470 5160
rect 2746 5148 2774 5188
rect 4246 5176 4252 5228
rect 4304 5216 4310 5228
rect 4433 5219 4491 5225
rect 4433 5216 4445 5219
rect 4304 5188 4445 5216
rect 4304 5176 4310 5188
rect 4433 5185 4445 5188
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 7101 5219 7159 5225
rect 7101 5185 7113 5219
rect 7147 5216 7159 5219
rect 7374 5216 7380 5228
rect 7147 5188 7380 5216
rect 7147 5185 7159 5188
rect 7101 5179 7159 5185
rect 7374 5176 7380 5188
rect 7432 5216 7438 5228
rect 7929 5219 7987 5225
rect 7929 5216 7941 5219
rect 7432 5188 7941 5216
rect 7432 5176 7438 5188
rect 7929 5185 7941 5188
rect 7975 5216 7987 5219
rect 8110 5216 8116 5228
rect 7975 5188 8116 5216
rect 7975 5185 7987 5188
rect 7929 5179 7987 5185
rect 8110 5176 8116 5188
rect 8168 5216 8174 5228
rect 9125 5219 9183 5225
rect 9125 5216 9137 5219
rect 8168 5188 9137 5216
rect 8168 5176 8174 5188
rect 9125 5185 9137 5188
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 2866 5148 2872 5160
rect 2464 5120 2509 5148
rect 2746 5120 2872 5148
rect 2464 5108 2470 5120
rect 2866 5108 2872 5120
rect 2924 5148 2930 5160
rect 3053 5151 3111 5157
rect 3053 5148 3065 5151
rect 2924 5120 3065 5148
rect 2924 5108 2930 5120
rect 3053 5117 3065 5120
rect 3099 5117 3111 5151
rect 3053 5111 3111 5117
rect 5353 5151 5411 5157
rect 5353 5117 5365 5151
rect 5399 5148 5411 5151
rect 5445 5151 5503 5157
rect 5445 5148 5457 5151
rect 5399 5120 5457 5148
rect 5399 5117 5411 5120
rect 5353 5111 5411 5117
rect 5445 5117 5457 5120
rect 5491 5117 5503 5151
rect 5445 5111 5503 5117
rect 5810 5108 5816 5160
rect 5868 5148 5874 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 5868 5120 6837 5148
rect 5868 5108 5874 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 8205 5151 8263 5157
rect 8205 5117 8217 5151
rect 8251 5148 8263 5151
rect 8294 5148 8300 5160
rect 8251 5120 8300 5148
rect 8251 5117 8263 5120
rect 8205 5111 8263 5117
rect 8294 5108 8300 5120
rect 8352 5108 8358 5160
rect 9398 5148 9404 5160
rect 9359 5120 9404 5148
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 10060 5157 10088 5256
rect 10226 5216 10232 5228
rect 10187 5188 10232 5216
rect 10226 5176 10232 5188
rect 10284 5176 10290 5228
rect 10888 5216 10916 5256
rect 11057 5253 11069 5287
rect 11103 5284 11115 5287
rect 11149 5287 11207 5293
rect 11149 5284 11161 5287
rect 11103 5256 11161 5284
rect 11103 5253 11115 5256
rect 11057 5247 11115 5253
rect 11149 5253 11161 5256
rect 11195 5253 11207 5287
rect 11149 5247 11207 5253
rect 12066 5216 12072 5228
rect 10888 5188 11376 5216
rect 12027 5188 12072 5216
rect 10045 5151 10103 5157
rect 10045 5148 10057 5151
rect 9646 5120 10057 5148
rect 2225 5083 2283 5089
rect 2225 5049 2237 5083
rect 2271 5049 2283 5083
rect 5074 5080 5080 5092
rect 5035 5052 5080 5080
rect 2225 5043 2283 5049
rect 2240 5012 2268 5043
rect 5074 5040 5080 5052
rect 5132 5040 5138 5092
rect 7098 5040 7104 5092
rect 7156 5080 7162 5092
rect 8113 5083 8171 5089
rect 8113 5080 8125 5083
rect 7156 5052 8125 5080
rect 7156 5040 7162 5052
rect 8113 5049 8125 5052
rect 8159 5049 8171 5083
rect 8113 5043 8171 5049
rect 8754 5040 8760 5092
rect 8812 5080 8818 5092
rect 9646 5080 9674 5120
rect 10045 5117 10057 5120
rect 10091 5117 10103 5151
rect 10594 5148 10600 5160
rect 10555 5120 10600 5148
rect 10045 5111 10103 5117
rect 10594 5108 10600 5120
rect 10652 5108 10658 5160
rect 10686 5108 10692 5160
rect 10744 5148 10750 5160
rect 11348 5157 11376 5188
rect 12066 5176 12072 5188
rect 12124 5176 12130 5228
rect 11333 5151 11391 5157
rect 10744 5120 10789 5148
rect 10744 5108 10750 5120
rect 11333 5117 11345 5151
rect 11379 5117 11391 5151
rect 11698 5148 11704 5160
rect 11611 5120 11704 5148
rect 11333 5111 11391 5117
rect 11698 5108 11704 5120
rect 11756 5108 11762 5160
rect 12253 5151 12311 5157
rect 12253 5117 12265 5151
rect 12299 5148 12311 5151
rect 12452 5148 12480 5312
rect 13354 5216 13360 5228
rect 13280 5188 13360 5216
rect 13280 5157 13308 5188
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 13740 5216 13768 5315
rect 15841 5287 15899 5293
rect 15841 5253 15853 5287
rect 15887 5284 15899 5287
rect 15933 5287 15991 5293
rect 15933 5284 15945 5287
rect 15887 5256 15945 5284
rect 15887 5253 15899 5256
rect 15841 5247 15899 5253
rect 15933 5253 15945 5256
rect 15979 5253 15991 5287
rect 15933 5247 15991 5253
rect 14737 5219 14795 5225
rect 13740 5188 14596 5216
rect 14568 5157 14596 5188
rect 14737 5185 14749 5219
rect 14783 5216 14795 5219
rect 15286 5216 15292 5228
rect 14783 5188 15292 5216
rect 14783 5185 14795 5188
rect 14737 5179 14795 5185
rect 14844 5157 14872 5188
rect 15286 5176 15292 5188
rect 15344 5216 15350 5228
rect 15344 5188 16160 5216
rect 15344 5176 15350 5188
rect 12713 5151 12771 5157
rect 12713 5148 12725 5151
rect 12299 5120 12725 5148
rect 12299 5117 12311 5120
rect 12253 5111 12311 5117
rect 12713 5117 12725 5120
rect 12759 5117 12771 5151
rect 12713 5111 12771 5117
rect 13265 5151 13323 5157
rect 13265 5117 13277 5151
rect 13311 5117 13323 5151
rect 13265 5111 13323 5117
rect 13725 5151 13783 5157
rect 13725 5117 13737 5151
rect 13771 5148 13783 5151
rect 13909 5151 13967 5157
rect 13909 5148 13921 5151
rect 13771 5120 13921 5148
rect 13771 5117 13783 5120
rect 13725 5111 13783 5117
rect 13909 5117 13921 5120
rect 13955 5117 13967 5151
rect 13909 5111 13967 5117
rect 14553 5151 14611 5157
rect 14553 5117 14565 5151
rect 14599 5117 14611 5151
rect 14553 5111 14611 5117
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5117 14887 5151
rect 15378 5148 15384 5160
rect 15339 5120 15384 5148
rect 14829 5111 14887 5117
rect 15378 5108 15384 5120
rect 15436 5148 15442 5160
rect 16132 5157 16160 5188
rect 15473 5151 15531 5157
rect 15473 5148 15485 5151
rect 15436 5120 15485 5148
rect 15436 5108 15442 5120
rect 15473 5117 15485 5120
rect 15519 5117 15531 5151
rect 15473 5111 15531 5117
rect 16117 5151 16175 5157
rect 16117 5117 16129 5151
rect 16163 5117 16175 5151
rect 16117 5111 16175 5117
rect 11716 5080 11744 5108
rect 8812 5052 9674 5080
rect 9784 5052 11744 5080
rect 8812 5040 8818 5052
rect 2777 5015 2835 5021
rect 2777 5012 2789 5015
rect 2240 4984 2789 5012
rect 2777 4981 2789 4984
rect 2823 5012 2835 5015
rect 2866 5012 2872 5024
rect 2823 4984 2872 5012
rect 2823 4981 2835 4984
rect 2777 4975 2835 4981
rect 2866 4972 2872 4984
rect 2924 4972 2930 5024
rect 5994 4972 6000 5024
rect 6052 5012 6058 5024
rect 6457 5015 6515 5021
rect 6457 5012 6469 5015
rect 6052 4984 6469 5012
rect 6052 4972 6058 4984
rect 6457 4981 6469 4984
rect 6503 4981 6515 5015
rect 6457 4975 6515 4981
rect 6917 5015 6975 5021
rect 6917 4981 6929 5015
rect 6963 5012 6975 5015
rect 8018 5012 8024 5024
rect 6963 4984 8024 5012
rect 6963 4981 6975 4984
rect 6917 4975 6975 4981
rect 8018 4972 8024 4984
rect 8076 4972 8082 5024
rect 8570 5012 8576 5024
rect 8531 4984 8576 5012
rect 8570 4972 8576 4984
rect 8628 4972 8634 5024
rect 8662 4972 8668 5024
rect 8720 5012 8726 5024
rect 9784 5021 9812 5052
rect 12434 5040 12440 5092
rect 12492 5080 12498 5092
rect 13817 5083 13875 5089
rect 13817 5080 13829 5083
rect 12492 5052 12537 5080
rect 13096 5052 13829 5080
rect 12492 5040 12498 5052
rect 9309 5015 9367 5021
rect 9309 5012 9321 5015
rect 8720 4984 9321 5012
rect 8720 4972 8726 4984
rect 9309 4981 9321 4984
rect 9355 4981 9367 5015
rect 9309 4975 9367 4981
rect 9769 5015 9827 5021
rect 9769 4981 9781 5015
rect 9815 4981 9827 5015
rect 9769 4975 9827 4981
rect 10226 4972 10232 5024
rect 10284 5012 10290 5024
rect 11057 5015 11115 5021
rect 11057 5012 11069 5015
rect 10284 4984 11069 5012
rect 10284 4972 10290 4984
rect 11057 4981 11069 4984
rect 11103 4981 11115 5015
rect 11057 4975 11115 4981
rect 12066 4972 12072 5024
rect 12124 5012 12130 5024
rect 13096 5012 13124 5052
rect 13817 5049 13829 5052
rect 13863 5049 13875 5083
rect 13817 5043 13875 5049
rect 14921 5083 14979 5089
rect 14921 5049 14933 5083
rect 14967 5049 14979 5083
rect 14921 5043 14979 5049
rect 12124 4984 13124 5012
rect 14936 5012 14964 5043
rect 15838 5012 15844 5024
rect 14936 4984 15844 5012
rect 12124 4972 12130 4984
rect 15838 4972 15844 4984
rect 15896 4972 15902 5024
rect 1104 4922 17296 4944
rect 1104 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 6571 4922
rect 6623 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 11904 4922
rect 11956 4870 11968 4922
rect 12020 4870 17296 4922
rect 1104 4848 17296 4870
rect 2774 4808 2780 4820
rect 2240 4780 2780 4808
rect 2240 4749 2268 4780
rect 2774 4768 2780 4780
rect 2832 4808 2838 4820
rect 5074 4808 5080 4820
rect 2832 4780 2877 4808
rect 4724 4780 5080 4808
rect 2832 4768 2838 4780
rect 2225 4743 2283 4749
rect 2225 4709 2237 4743
rect 2271 4709 2283 4743
rect 2866 4740 2872 4752
rect 2827 4712 2872 4740
rect 2225 4703 2283 4709
rect 2866 4700 2872 4712
rect 2924 4700 2930 4752
rect 4246 4700 4252 4752
rect 4304 4740 4310 4752
rect 4617 4743 4675 4749
rect 4617 4740 4629 4743
rect 4304 4712 4629 4740
rect 4304 4700 4310 4712
rect 4617 4709 4629 4712
rect 4663 4709 4675 4743
rect 4617 4703 4675 4709
rect 1765 4675 1823 4681
rect 1765 4641 1777 4675
rect 1811 4641 1823 4675
rect 1765 4635 1823 4641
rect 2317 4675 2375 4681
rect 2317 4641 2329 4675
rect 2363 4672 2375 4675
rect 2958 4672 2964 4684
rect 2363 4644 2964 4672
rect 2363 4641 2375 4644
rect 2317 4635 2375 4641
rect 1780 4604 1808 4635
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 4341 4675 4399 4681
rect 4341 4641 4353 4675
rect 4387 4672 4399 4675
rect 4724 4672 4752 4780
rect 5074 4768 5080 4780
rect 5132 4808 5138 4820
rect 5132 4780 7880 4808
rect 5132 4768 5138 4780
rect 4801 4743 4859 4749
rect 4801 4709 4813 4743
rect 4847 4740 4859 4743
rect 4847 4712 5580 4740
rect 4847 4709 4859 4712
rect 4801 4703 4859 4709
rect 4387 4644 4752 4672
rect 4893 4675 4951 4681
rect 4387 4641 4399 4644
rect 4341 4635 4399 4641
rect 4893 4641 4905 4675
rect 4939 4641 4951 4675
rect 4893 4635 4951 4641
rect 2406 4604 2412 4616
rect 1780 4576 2412 4604
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4604 4491 4607
rect 4908 4604 4936 4635
rect 4479 4576 4936 4604
rect 5552 4604 5580 4712
rect 5644 4681 5672 4780
rect 6656 4749 6684 4780
rect 6641 4743 6699 4749
rect 5736 4712 6040 4740
rect 5629 4675 5687 4681
rect 5629 4641 5641 4675
rect 5675 4641 5687 4675
rect 5629 4635 5687 4641
rect 5736 4604 5764 4712
rect 6012 4684 6040 4712
rect 6641 4709 6653 4743
rect 6687 4709 6699 4743
rect 7745 4743 7803 4749
rect 7745 4740 7757 4743
rect 6641 4703 6699 4709
rect 6932 4712 7757 4740
rect 5813 4675 5871 4681
rect 5813 4641 5825 4675
rect 5859 4641 5871 4675
rect 5994 4672 6000 4684
rect 5955 4644 6000 4672
rect 5813 4635 5871 4641
rect 5552 4576 5764 4604
rect 4479 4573 4491 4576
rect 4433 4567 4491 4573
rect 2777 4539 2835 4545
rect 2777 4505 2789 4539
rect 2823 4536 2835 4539
rect 2961 4539 3019 4545
rect 2961 4536 2973 4539
rect 2823 4508 2973 4536
rect 2823 4505 2835 4508
rect 2777 4499 2835 4505
rect 2961 4505 2973 4508
rect 3007 4505 3019 4539
rect 5828 4536 5856 4635
rect 5994 4632 6000 4644
rect 6052 4632 6058 4684
rect 6932 4681 6960 4712
rect 7745 4709 7757 4712
rect 7791 4709 7803 4743
rect 7745 4703 7803 4709
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4641 6975 4675
rect 6917 4635 6975 4641
rect 7009 4675 7067 4681
rect 7009 4641 7021 4675
rect 7055 4641 7067 4675
rect 7282 4672 7288 4684
rect 7009 4635 7067 4641
rect 7116 4644 7288 4672
rect 6822 4564 6828 4616
rect 6880 4604 6886 4616
rect 7024 4604 7052 4635
rect 6880 4576 7052 4604
rect 6880 4564 6886 4576
rect 7116 4536 7144 4644
rect 7282 4632 7288 4644
rect 7340 4672 7346 4684
rect 7561 4675 7619 4681
rect 7561 4672 7573 4675
rect 7340 4644 7573 4672
rect 7340 4632 7346 4644
rect 7561 4641 7573 4644
rect 7607 4641 7619 4675
rect 7561 4635 7619 4641
rect 7653 4675 7711 4681
rect 7653 4641 7665 4675
rect 7699 4641 7711 4675
rect 7653 4635 7711 4641
rect 7374 4604 7380 4616
rect 7335 4576 7380 4604
rect 7374 4564 7380 4576
rect 7432 4604 7438 4616
rect 7668 4604 7696 4635
rect 7432 4576 7696 4604
rect 7432 4564 7438 4576
rect 5828 4508 7144 4536
rect 7852 4536 7880 4780
rect 14366 4768 14372 4820
rect 14424 4808 14430 4820
rect 14921 4811 14979 4817
rect 14921 4808 14933 4811
rect 14424 4780 14933 4808
rect 14424 4768 14430 4780
rect 14921 4777 14933 4780
rect 14967 4777 14979 4811
rect 14921 4771 14979 4777
rect 15289 4811 15347 4817
rect 15289 4777 15301 4811
rect 15335 4808 15347 4811
rect 15378 4808 15384 4820
rect 15335 4780 15384 4808
rect 15335 4777 15347 4780
rect 15289 4771 15347 4777
rect 15378 4768 15384 4780
rect 15436 4768 15442 4820
rect 16761 4811 16819 4817
rect 16761 4777 16773 4811
rect 16807 4777 16819 4811
rect 16761 4771 16819 4777
rect 8018 4700 8024 4752
rect 8076 4740 8082 4752
rect 16776 4740 16804 4771
rect 8076 4712 16804 4740
rect 8076 4700 8082 4712
rect 8205 4675 8263 4681
rect 8205 4641 8217 4675
rect 8251 4641 8263 4675
rect 8754 4672 8760 4684
rect 8715 4644 8760 4672
rect 8205 4635 8263 4641
rect 8220 4604 8248 4635
rect 8754 4632 8760 4644
rect 8812 4672 8818 4684
rect 9493 4675 9551 4681
rect 8812 4644 9444 4672
rect 8812 4632 8818 4644
rect 8570 4604 8576 4616
rect 8220 4576 8576 4604
rect 8570 4564 8576 4576
rect 8628 4604 8634 4616
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 8628 4576 9137 4604
rect 8628 4564 8634 4576
rect 9125 4573 9137 4576
rect 9171 4573 9183 4607
rect 9416 4604 9444 4644
rect 9493 4641 9505 4675
rect 9539 4672 9551 4675
rect 10134 4672 10140 4684
rect 9539 4644 10140 4672
rect 9539 4641 9551 4644
rect 9493 4635 9551 4641
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 11054 4672 11060 4684
rect 11015 4644 11060 4672
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 16942 4672 16948 4684
rect 16903 4644 16948 4672
rect 16942 4632 16948 4644
rect 17000 4632 17006 4684
rect 10873 4607 10931 4613
rect 10873 4604 10885 4607
rect 9416 4576 10885 4604
rect 9125 4567 9183 4573
rect 10873 4573 10885 4576
rect 10919 4573 10931 4607
rect 10873 4567 10931 4573
rect 12526 4564 12532 4616
rect 12584 4604 12590 4616
rect 14645 4607 14703 4613
rect 14645 4604 14657 4607
rect 12584 4576 14657 4604
rect 12584 4564 12590 4576
rect 14645 4573 14657 4576
rect 14691 4573 14703 4607
rect 14645 4567 14703 4573
rect 14829 4607 14887 4613
rect 14829 4573 14841 4607
rect 14875 4604 14887 4607
rect 15378 4604 15384 4616
rect 14875 4576 15384 4604
rect 14875 4573 14887 4576
rect 14829 4567 14887 4573
rect 15378 4564 15384 4576
rect 15436 4564 15442 4616
rect 12434 4536 12440 4548
rect 7852 4508 12440 4536
rect 2961 4499 3019 4505
rect 12434 4496 12440 4508
rect 12492 4496 12498 4548
rect 4154 4468 4160 4480
rect 4115 4440 4160 4468
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 8570 4428 8576 4480
rect 8628 4468 8634 4480
rect 8757 4471 8815 4477
rect 8757 4468 8769 4471
rect 8628 4440 8769 4468
rect 8628 4428 8634 4440
rect 8757 4437 8769 4440
rect 8803 4468 8815 4471
rect 9493 4471 9551 4477
rect 9493 4468 9505 4471
rect 8803 4440 9505 4468
rect 8803 4437 8815 4440
rect 8757 4431 8815 4437
rect 9493 4437 9505 4440
rect 9539 4437 9551 4471
rect 9493 4431 9551 4437
rect 1104 4378 17296 4400
rect 1104 4326 3680 4378
rect 3732 4326 3744 4378
rect 3796 4326 3808 4378
rect 3860 4326 3872 4378
rect 3924 4326 9078 4378
rect 9130 4326 9142 4378
rect 9194 4326 9206 4378
rect 9258 4326 9270 4378
rect 9322 4326 14475 4378
rect 14527 4326 14539 4378
rect 14591 4326 14603 4378
rect 14655 4326 14667 4378
rect 14719 4326 17296 4378
rect 1104 4304 17296 4326
rect 7009 4267 7067 4273
rect 7009 4233 7021 4267
rect 7055 4264 7067 4267
rect 7374 4264 7380 4276
rect 7055 4236 7380 4264
rect 7055 4233 7067 4236
rect 7009 4227 7067 4233
rect 7374 4224 7380 4236
rect 7432 4224 7438 4276
rect 12069 4199 12127 4205
rect 12069 4165 12081 4199
rect 12115 4165 12127 4199
rect 12069 4159 12127 4165
rect 1394 4128 1400 4140
rect 1355 4100 1400 4128
rect 1394 4088 1400 4100
rect 1452 4088 1458 4140
rect 2038 4088 2044 4140
rect 2096 4128 2102 4140
rect 6641 4131 6699 4137
rect 2096 4100 4660 4128
rect 2096 4088 2102 4100
rect 4154 4060 4160 4072
rect 4115 4032 4160 4060
rect 4154 4020 4160 4032
rect 4212 4020 4218 4072
rect 4632 4060 4660 4100
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 6822 4128 6828 4140
rect 6687 4100 6828 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 12084 4128 12112 4159
rect 12710 4128 12716 4140
rect 6932 4100 12112 4128
rect 12671 4100 12716 4128
rect 6932 4060 6960 4100
rect 12710 4088 12716 4100
rect 12768 4088 12774 4140
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4128 13323 4131
rect 13630 4128 13636 4140
rect 13311 4100 13636 4128
rect 13311 4097 13323 4100
rect 13265 4091 13323 4097
rect 13630 4088 13636 4100
rect 13688 4128 13694 4140
rect 14277 4131 14335 4137
rect 14277 4128 14289 4131
rect 13688 4100 14289 4128
rect 13688 4088 13694 4100
rect 14277 4097 14289 4100
rect 14323 4097 14335 4131
rect 14277 4091 14335 4097
rect 4632 4032 6960 4060
rect 7006 4020 7012 4072
rect 7064 4060 7070 4072
rect 7282 4060 7288 4072
rect 7064 4032 7109 4060
rect 7243 4032 7288 4060
rect 7064 4020 7070 4032
rect 7282 4020 7288 4032
rect 7340 4020 7346 4072
rect 13449 4063 13507 4069
rect 13449 4029 13461 4063
rect 13495 4029 13507 4063
rect 13449 4023 13507 4029
rect 13725 4063 13783 4069
rect 13725 4029 13737 4063
rect 13771 4060 13783 4063
rect 13814 4060 13820 4072
rect 13771 4032 13820 4060
rect 13771 4029 13783 4032
rect 13725 4023 13783 4029
rect 1578 3992 1584 4004
rect 1539 3964 1584 3992
rect 1578 3952 1584 3964
rect 1636 3952 1642 4004
rect 4706 3992 4712 4004
rect 4619 3964 4712 3992
rect 4706 3952 4712 3964
rect 4764 3992 4770 4004
rect 12529 3995 12587 4001
rect 12529 3992 12541 3995
rect 4764 3964 12541 3992
rect 4764 3952 4770 3964
rect 12529 3961 12541 3964
rect 12575 3961 12587 3995
rect 12529 3955 12587 3961
rect 13262 3952 13268 4004
rect 13320 3992 13326 4004
rect 13464 3992 13492 4023
rect 13814 4020 13820 4032
rect 13872 4020 13878 4072
rect 14182 4060 14188 4072
rect 14143 4032 14188 4060
rect 14182 4020 14188 4032
rect 14240 4020 14246 4072
rect 14274 3992 14280 4004
rect 13320 3964 14280 3992
rect 13320 3952 13326 3964
rect 14274 3952 14280 3964
rect 14332 3992 14338 4004
rect 16850 3992 16856 4004
rect 14332 3964 16856 3992
rect 14332 3952 14338 3964
rect 16850 3952 16856 3964
rect 16908 3952 16914 4004
rect 7006 3884 7012 3936
rect 7064 3924 7070 3936
rect 7101 3927 7159 3933
rect 7101 3924 7113 3927
rect 7064 3896 7113 3924
rect 7064 3884 7070 3896
rect 7101 3893 7113 3896
rect 7147 3893 7159 3927
rect 7101 3887 7159 3893
rect 7190 3884 7196 3936
rect 7248 3924 7254 3936
rect 11330 3924 11336 3936
rect 7248 3896 11336 3924
rect 7248 3884 7254 3896
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 13170 3924 13176 3936
rect 12492 3896 12537 3924
rect 13131 3896 13176 3924
rect 12492 3884 12498 3896
rect 13170 3884 13176 3896
rect 13228 3884 13234 3936
rect 14366 3924 14372 3936
rect 14327 3896 14372 3924
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 1104 3834 17296 3856
rect 1104 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 6571 3834
rect 6623 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 11904 3834
rect 11956 3782 11968 3834
rect 12020 3782 17296 3834
rect 1104 3760 17296 3782
rect 3421 3723 3479 3729
rect 3421 3689 3433 3723
rect 3467 3720 3479 3723
rect 9769 3723 9827 3729
rect 3467 3692 8708 3720
rect 3467 3689 3479 3692
rect 3421 3683 3479 3689
rect 2774 3612 2780 3664
rect 2832 3652 2838 3664
rect 3329 3655 3387 3661
rect 3329 3652 3341 3655
rect 2832 3624 3341 3652
rect 2832 3612 2838 3624
rect 3329 3621 3341 3624
rect 3375 3621 3387 3655
rect 3329 3615 3387 3621
rect 5258 3612 5264 3664
rect 5316 3612 5322 3664
rect 6825 3655 6883 3661
rect 6825 3621 6837 3655
rect 6871 3652 6883 3655
rect 7282 3652 7288 3664
rect 6871 3624 7288 3652
rect 6871 3621 6883 3624
rect 6825 3615 6883 3621
rect 7282 3612 7288 3624
rect 7340 3612 7346 3664
rect 8570 3652 8576 3664
rect 8531 3624 8576 3652
rect 8570 3612 8576 3624
rect 8628 3612 8634 3664
rect 1578 3544 1584 3596
rect 1636 3584 1642 3596
rect 3973 3587 4031 3593
rect 3973 3584 3985 3587
rect 1636 3556 3985 3584
rect 1636 3544 1642 3556
rect 3973 3553 3985 3556
rect 4019 3553 4031 3587
rect 6086 3584 6092 3596
rect 6047 3556 6092 3584
rect 3973 3547 4031 3553
rect 3988 3516 4016 3547
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 7009 3587 7067 3593
rect 7009 3553 7021 3587
rect 7055 3584 7067 3587
rect 7466 3584 7472 3596
rect 7055 3556 7472 3584
rect 7055 3553 7067 3556
rect 7009 3547 7067 3553
rect 7466 3544 7472 3556
rect 7524 3584 7530 3596
rect 8389 3587 8447 3593
rect 8389 3584 8401 3587
rect 7524 3556 8401 3584
rect 7524 3544 7530 3556
rect 8389 3553 8401 3556
rect 8435 3553 8447 3587
rect 8680 3584 8708 3692
rect 9769 3689 9781 3723
rect 9815 3720 9827 3723
rect 10318 3720 10324 3732
rect 9815 3692 10324 3720
rect 9815 3689 9827 3692
rect 9769 3683 9827 3689
rect 10318 3680 10324 3692
rect 10376 3680 10382 3732
rect 11054 3720 11060 3732
rect 10520 3692 11060 3720
rect 10520 3661 10548 3692
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 13630 3680 13636 3732
rect 13688 3720 13694 3732
rect 13725 3723 13783 3729
rect 13725 3720 13737 3723
rect 13688 3692 13737 3720
rect 13688 3680 13694 3692
rect 13725 3689 13737 3692
rect 13771 3689 13783 3723
rect 13725 3683 13783 3689
rect 10505 3655 10563 3661
rect 10505 3621 10517 3655
rect 10551 3621 10563 3655
rect 10505 3615 10563 3621
rect 12710 3612 12716 3664
rect 12768 3652 12774 3664
rect 12897 3655 12955 3661
rect 12897 3652 12909 3655
rect 12768 3624 12909 3652
rect 12768 3612 12774 3624
rect 12897 3621 12909 3624
rect 12943 3621 12955 3655
rect 13814 3652 13820 3664
rect 12897 3615 12955 3621
rect 13556 3624 13820 3652
rect 10137 3587 10195 3593
rect 10137 3584 10149 3587
rect 8680 3556 10149 3584
rect 8389 3547 8447 3553
rect 10137 3553 10149 3556
rect 10183 3584 10195 3587
rect 10413 3587 10471 3593
rect 10413 3584 10425 3587
rect 10183 3556 10425 3584
rect 10183 3553 10195 3556
rect 10137 3547 10195 3553
rect 10413 3553 10425 3556
rect 10459 3584 10471 3587
rect 10594 3584 10600 3596
rect 10459 3556 10600 3584
rect 10459 3553 10471 3556
rect 10413 3547 10471 3553
rect 10594 3544 10600 3556
rect 10652 3544 10658 3596
rect 10962 3584 10968 3596
rect 10923 3556 10968 3584
rect 10962 3544 10968 3556
rect 11020 3584 11026 3596
rect 11425 3587 11483 3593
rect 11425 3584 11437 3587
rect 11020 3556 11437 3584
rect 11020 3544 11026 3556
rect 11425 3553 11437 3556
rect 11471 3553 11483 3587
rect 13262 3584 13268 3596
rect 13223 3556 13268 3584
rect 11425 3547 11483 3553
rect 13262 3544 13268 3556
rect 13320 3544 13326 3596
rect 13556 3593 13584 3624
rect 13814 3612 13820 3624
rect 13872 3612 13878 3664
rect 15470 3612 15476 3664
rect 15528 3612 15534 3664
rect 13541 3587 13599 3593
rect 13541 3553 13553 3587
rect 13587 3553 13599 3587
rect 13541 3547 13599 3553
rect 13633 3587 13691 3593
rect 13633 3553 13645 3587
rect 13679 3553 13691 3587
rect 13633 3547 13691 3553
rect 16761 3587 16819 3593
rect 16761 3553 16773 3587
rect 16807 3584 16819 3587
rect 17034 3584 17040 3596
rect 16807 3556 17040 3584
rect 16807 3553 16819 3556
rect 16761 3547 16819 3553
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 3988 3488 5733 3516
rect 5721 3485 5733 3488
rect 5767 3516 5779 3519
rect 5767 3488 5948 3516
rect 5767 3485 5779 3488
rect 5721 3479 5779 3485
rect 5920 3448 5948 3488
rect 5994 3476 6000 3528
rect 6052 3516 6058 3528
rect 7190 3516 7196 3528
rect 6052 3488 7196 3516
rect 6052 3476 6058 3488
rect 7190 3476 7196 3488
rect 7248 3476 7254 3528
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3516 7435 3519
rect 7650 3516 7656 3528
rect 7423 3488 7656 3516
rect 7423 3485 7435 3488
rect 7377 3479 7435 3485
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 7745 3519 7803 3525
rect 7745 3485 7757 3519
rect 7791 3516 7803 3519
rect 8018 3516 8024 3528
rect 7791 3488 8024 3516
rect 7791 3485 7803 3488
rect 7745 3479 7803 3485
rect 8018 3476 8024 3488
rect 8076 3476 8082 3528
rect 9398 3516 9404 3528
rect 9359 3488 9404 3516
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 11054 3516 11060 3528
rect 11015 3488 11060 3516
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13081 3519 13139 3525
rect 13081 3516 13093 3519
rect 13044 3488 13093 3516
rect 13044 3476 13050 3488
rect 13081 3485 13093 3488
rect 13127 3516 13139 3519
rect 13648 3516 13676 3547
rect 13127 3488 13676 3516
rect 14737 3519 14795 3525
rect 13127 3485 13139 3488
rect 13081 3479 13139 3485
rect 14737 3485 14749 3519
rect 14783 3485 14795 3519
rect 15010 3516 15016 3528
rect 14923 3488 15016 3516
rect 14737 3479 14795 3485
rect 9769 3451 9827 3457
rect 5920 3420 9674 3448
rect 7374 3380 7380 3392
rect 7335 3352 7380 3380
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 9646 3380 9674 3420
rect 9769 3417 9781 3451
rect 9815 3448 9827 3451
rect 9953 3451 10011 3457
rect 9953 3448 9965 3451
rect 9815 3420 9965 3448
rect 9815 3417 9827 3420
rect 9769 3411 9827 3417
rect 9953 3417 9965 3420
rect 9999 3417 10011 3451
rect 13722 3448 13728 3460
rect 9953 3411 10011 3417
rect 10060 3420 13728 3448
rect 10060 3380 10088 3420
rect 13722 3408 13728 3420
rect 13780 3448 13786 3460
rect 14752 3448 14780 3479
rect 15010 3476 15016 3488
rect 15068 3516 15074 3528
rect 16776 3516 16804 3547
rect 17034 3544 17040 3556
rect 17092 3544 17098 3596
rect 15068 3488 16804 3516
rect 15068 3476 15074 3488
rect 13780 3420 14780 3448
rect 13780 3408 13786 3420
rect 9646 3352 10088 3380
rect 10134 3340 10140 3392
rect 10192 3380 10198 3392
rect 15470 3380 15476 3392
rect 10192 3352 15476 3380
rect 10192 3340 10198 3352
rect 15470 3340 15476 3352
rect 15528 3340 15534 3392
rect 1104 3290 17296 3312
rect 1104 3238 3680 3290
rect 3732 3238 3744 3290
rect 3796 3238 3808 3290
rect 3860 3238 3872 3290
rect 3924 3238 9078 3290
rect 9130 3238 9142 3290
rect 9194 3238 9206 3290
rect 9258 3238 9270 3290
rect 9322 3238 14475 3290
rect 14527 3238 14539 3290
rect 14591 3238 14603 3290
rect 14655 3238 14667 3290
rect 14719 3238 17296 3290
rect 1104 3216 17296 3238
rect 7374 3136 7380 3188
rect 7432 3176 7438 3188
rect 7469 3179 7527 3185
rect 7469 3176 7481 3179
rect 7432 3148 7481 3176
rect 7432 3136 7438 3148
rect 7469 3145 7481 3148
rect 7515 3145 7527 3179
rect 7469 3139 7527 3145
rect 7650 3136 7656 3188
rect 7708 3176 7714 3188
rect 8113 3179 8171 3185
rect 8113 3176 8125 3179
rect 7708 3148 8125 3176
rect 7708 3136 7714 3148
rect 8113 3145 8125 3148
rect 8159 3145 8171 3179
rect 8113 3139 8171 3145
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 9953 3179 10011 3185
rect 9953 3176 9965 3179
rect 9456 3148 9965 3176
rect 9456 3136 9462 3148
rect 9953 3145 9965 3148
rect 9999 3145 10011 3179
rect 9953 3139 10011 3145
rect 7282 3108 7288 3120
rect 7208 3080 7288 3108
rect 1578 3000 1584 3052
rect 1636 3040 1642 3052
rect 1765 3043 1823 3049
rect 1765 3040 1777 3043
rect 1636 3012 1777 3040
rect 1636 3000 1642 3012
rect 1765 3009 1777 3012
rect 1811 3040 1823 3043
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 1811 3012 2513 3040
rect 1811 3009 1823 3012
rect 1765 3003 1823 3009
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 3142 3000 3148 3052
rect 3200 3040 3206 3052
rect 5994 3040 6000 3052
rect 3200 3012 6000 3040
rect 3200 3000 3206 3012
rect 474 2932 480 2984
rect 532 2972 538 2984
rect 2406 2981 2412 2984
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 532 2944 1409 2972
rect 532 2932 538 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 2271 2975 2329 2981
rect 2271 2972 2283 2975
rect 1903 2944 2283 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 2271 2941 2283 2944
rect 2317 2941 2329 2975
rect 2271 2935 2329 2941
rect 2374 2975 2412 2981
rect 2374 2941 2386 2975
rect 2374 2935 2412 2941
rect 2406 2932 2412 2935
rect 2464 2932 2470 2984
rect 4540 2981 4568 3012
rect 5994 3000 6000 3012
rect 6052 3000 6058 3052
rect 6086 3000 6092 3052
rect 6144 3040 6150 3052
rect 7208 3049 7236 3080
rect 7282 3068 7288 3080
rect 7340 3068 7346 3120
rect 8018 3068 8024 3120
rect 8076 3108 8082 3120
rect 8389 3111 8447 3117
rect 8389 3108 8401 3111
rect 8076 3080 8401 3108
rect 8076 3068 8082 3080
rect 8389 3077 8401 3080
rect 8435 3077 8447 3111
rect 8389 3071 8447 3077
rect 8772 3080 8984 3108
rect 6457 3043 6515 3049
rect 6457 3040 6469 3043
rect 6144 3012 6469 3040
rect 6144 3000 6150 3012
rect 6457 3009 6469 3012
rect 6503 3009 6515 3043
rect 6457 3003 6515 3009
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 8110 3000 8116 3052
rect 8168 3040 8174 3052
rect 8772 3040 8800 3080
rect 8168 3012 8800 3040
rect 8168 3000 8174 3012
rect 8846 3000 8852 3052
rect 8904 3000 8910 3052
rect 8956 3049 8984 3080
rect 8941 3043 8999 3049
rect 8941 3009 8953 3043
rect 8987 3040 8999 3043
rect 9309 3043 9367 3049
rect 9309 3040 9321 3043
rect 8987 3012 9321 3040
rect 8987 3009 8999 3012
rect 8941 3003 8999 3009
rect 9309 3009 9321 3012
rect 9355 3009 9367 3043
rect 9309 3003 9367 3009
rect 9493 3043 9551 3049
rect 9493 3009 9505 3043
rect 9539 3040 9551 3043
rect 9539 3012 9904 3040
rect 9539 3009 9551 3012
rect 9493 3003 9551 3009
rect 4525 2975 4583 2981
rect 4525 2941 4537 2975
rect 4571 2941 4583 2975
rect 7282 2972 7288 2984
rect 7243 2944 7288 2972
rect 4525 2935 4583 2941
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 7466 2972 7472 2984
rect 7427 2944 7472 2972
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 8018 2972 8024 2984
rect 7979 2944 8024 2972
rect 8018 2932 8024 2944
rect 8076 2932 8082 2984
rect 8297 2975 8355 2981
rect 8297 2941 8309 2975
rect 8343 2941 8355 2975
rect 8297 2935 8355 2941
rect 8757 2975 8815 2981
rect 8757 2941 8769 2975
rect 8803 2972 8815 2975
rect 8864 2972 8892 3000
rect 9582 2972 9588 2984
rect 8803 2944 8892 2972
rect 9543 2944 9588 2972
rect 8803 2941 8815 2944
rect 8757 2935 8815 2941
rect 2777 2907 2835 2913
rect 2777 2873 2789 2907
rect 2823 2904 2835 2907
rect 3050 2904 3056 2916
rect 2823 2876 3056 2904
rect 2823 2873 2835 2876
rect 2777 2867 2835 2873
rect 3050 2864 3056 2876
rect 3108 2864 3114 2916
rect 7484 2904 7512 2932
rect 8312 2904 8340 2935
rect 9582 2932 9588 2944
rect 9640 2932 9646 2984
rect 1581 2839 1639 2845
rect 1581 2805 1593 2839
rect 1627 2836 1639 2839
rect 1670 2836 1676 2848
rect 1627 2808 1676 2836
rect 1627 2805 1639 2808
rect 1581 2799 1639 2805
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 3988 2836 4016 2890
rect 7484 2876 8340 2904
rect 8849 2907 8907 2913
rect 8849 2873 8861 2907
rect 8895 2904 8907 2907
rect 9674 2904 9680 2916
rect 8895 2876 9680 2904
rect 8895 2873 8907 2876
rect 8849 2867 8907 2873
rect 9674 2864 9680 2876
rect 9732 2864 9738 2916
rect 9876 2904 9904 3012
rect 9968 2972 9996 3139
rect 10318 3136 10324 3188
rect 10376 3176 10382 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 10376 3148 10609 3176
rect 10376 3136 10382 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 10781 3179 10839 3185
rect 10781 3145 10793 3179
rect 10827 3176 10839 3179
rect 10962 3176 10968 3188
rect 10827 3148 10968 3176
rect 10827 3145 10839 3148
rect 10781 3139 10839 3145
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 13265 3179 13323 3185
rect 13265 3176 13277 3179
rect 12492 3148 12537 3176
rect 13004 3148 13277 3176
rect 12492 3136 12498 3148
rect 11425 3043 11483 3049
rect 11425 3009 11437 3043
rect 11471 3040 11483 3043
rect 12526 3040 12532 3052
rect 11471 3012 12532 3040
rect 11471 3009 11483 3012
rect 11425 3003 11483 3009
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 10045 2975 10103 2981
rect 10045 2972 10057 2975
rect 9968 2944 10057 2972
rect 10045 2941 10057 2944
rect 10091 2941 10103 2975
rect 10594 2972 10600 2984
rect 10555 2944 10600 2972
rect 10045 2935 10103 2941
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 11330 2932 11336 2984
rect 11388 2972 11394 2984
rect 12897 2975 12955 2981
rect 12897 2972 12909 2975
rect 11388 2944 12909 2972
rect 11388 2932 11394 2944
rect 12897 2941 12909 2944
rect 12943 2941 12955 2975
rect 12897 2935 12955 2941
rect 10962 2904 10968 2916
rect 9876 2876 10968 2904
rect 10962 2864 10968 2876
rect 11020 2864 11026 2916
rect 12805 2907 12863 2913
rect 12805 2873 12817 2907
rect 12851 2904 12863 2907
rect 13004 2904 13032 3148
rect 13265 3145 13277 3148
rect 13311 3145 13323 3179
rect 14182 3176 14188 3188
rect 14143 3148 14188 3176
rect 13265 3139 13323 3145
rect 14182 3136 14188 3148
rect 14240 3136 14246 3188
rect 15378 3176 15384 3188
rect 15339 3148 15384 3176
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 16574 3176 16580 3188
rect 16535 3148 16580 3176
rect 16574 3136 16580 3148
rect 16632 3136 16638 3188
rect 16301 3111 16359 3117
rect 16301 3108 16313 3111
rect 13556 3080 16313 3108
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 13170 3040 13176 3052
rect 13127 3012 13176 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 13170 3000 13176 3012
rect 13228 3000 13234 3052
rect 12851 2876 13032 2904
rect 12851 2873 12863 2876
rect 12805 2867 12863 2873
rect 5258 2836 5264 2848
rect 3988 2808 5264 2836
rect 5258 2796 5264 2808
rect 5316 2836 5322 2848
rect 10134 2836 10140 2848
rect 5316 2808 10140 2836
rect 5316 2796 5322 2808
rect 10134 2796 10140 2808
rect 10192 2796 10198 2848
rect 10502 2796 10508 2848
rect 10560 2836 10566 2848
rect 11149 2839 11207 2845
rect 11149 2836 11161 2839
rect 10560 2808 11161 2836
rect 10560 2796 10566 2808
rect 11149 2805 11161 2808
rect 11195 2805 11207 2839
rect 11149 2799 11207 2805
rect 11241 2839 11299 2845
rect 11241 2805 11253 2839
rect 11287 2836 11299 2839
rect 13556 2836 13584 3080
rect 16301 3077 16313 3080
rect 16347 3077 16359 3111
rect 16301 3071 16359 3077
rect 13630 3000 13636 3052
rect 13688 3040 13694 3052
rect 13817 3043 13875 3049
rect 13817 3040 13829 3043
rect 13688 3012 13829 3040
rect 13688 3000 13694 3012
rect 13817 3009 13829 3012
rect 13863 3009 13875 3043
rect 13817 3003 13875 3009
rect 14366 3000 14372 3052
rect 14424 3040 14430 3052
rect 15105 3043 15163 3049
rect 15105 3040 15117 3043
rect 14424 3012 15117 3040
rect 14424 3000 14430 3012
rect 15105 3009 15117 3012
rect 15151 3009 15163 3043
rect 15105 3003 15163 3009
rect 13722 2972 13728 2984
rect 13683 2944 13728 2972
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 14274 2972 14280 2984
rect 14235 2944 14280 2972
rect 14274 2932 14280 2944
rect 14332 2932 14338 2984
rect 15010 2972 15016 2984
rect 14971 2944 15016 2972
rect 15010 2932 15016 2944
rect 15068 2932 15074 2984
rect 15194 2932 15200 2984
rect 15252 2972 15258 2984
rect 15565 2975 15623 2981
rect 15565 2972 15577 2975
rect 15252 2944 15577 2972
rect 15252 2932 15258 2944
rect 15565 2941 15577 2944
rect 15611 2941 15623 2975
rect 16482 2972 16488 2984
rect 16443 2944 16488 2972
rect 15565 2935 15623 2941
rect 16482 2932 16488 2944
rect 16540 2932 16546 2984
rect 16758 2972 16764 2984
rect 16719 2944 16764 2972
rect 16758 2932 16764 2944
rect 16816 2932 16822 2984
rect 13633 2907 13691 2913
rect 13633 2873 13645 2907
rect 13679 2904 13691 2907
rect 13679 2876 14596 2904
rect 13679 2873 13691 2876
rect 13633 2867 13691 2873
rect 14568 2845 14596 2876
rect 11287 2808 13584 2836
rect 14553 2839 14611 2845
rect 11287 2805 11299 2808
rect 11241 2799 11299 2805
rect 14553 2805 14565 2839
rect 14599 2805 14611 2839
rect 14918 2836 14924 2848
rect 14879 2808 14924 2836
rect 14553 2799 14611 2805
rect 14918 2796 14924 2808
rect 14976 2796 14982 2848
rect 1104 2746 17296 2768
rect 1104 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 6571 2746
rect 6623 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 11904 2746
rect 11956 2694 11968 2746
rect 12020 2694 17296 2746
rect 1104 2672 17296 2694
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 2130 2632 2136 2644
rect 1903 2604 2136 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 2130 2592 2136 2604
rect 2188 2592 2194 2644
rect 2225 2635 2283 2641
rect 2225 2601 2237 2635
rect 2271 2632 2283 2635
rect 7098 2632 7104 2644
rect 2271 2604 6914 2632
rect 7059 2604 7104 2632
rect 2271 2601 2283 2604
rect 2225 2595 2283 2601
rect 1578 2564 1584 2576
rect 1539 2536 1584 2564
rect 1578 2524 1584 2536
rect 1636 2524 1642 2576
rect 6886 2564 6914 2604
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 7374 2632 7380 2644
rect 7335 2604 7380 2632
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 8386 2592 8392 2644
rect 8444 2592 8450 2644
rect 9674 2632 9680 2644
rect 9635 2604 9680 2632
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 10410 2592 10416 2644
rect 10468 2632 10474 2644
rect 10597 2635 10655 2641
rect 10597 2632 10609 2635
rect 10468 2604 10609 2632
rect 10468 2592 10474 2604
rect 10597 2601 10609 2604
rect 10643 2601 10655 2635
rect 10597 2595 10655 2601
rect 10689 2635 10747 2641
rect 10689 2601 10701 2635
rect 10735 2632 10747 2635
rect 11054 2632 11060 2644
rect 10735 2604 11060 2632
rect 10735 2601 10747 2604
rect 10689 2595 10747 2601
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 13630 2632 13636 2644
rect 13591 2604 13636 2632
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 14182 2592 14188 2644
rect 14240 2592 14246 2644
rect 14918 2632 14924 2644
rect 14660 2604 14924 2632
rect 8404 2564 8432 2592
rect 2976 2536 5856 2564
rect 6886 2536 8432 2564
rect 8573 2567 8631 2573
rect 1670 2456 1676 2508
rect 1728 2496 1734 2508
rect 1765 2499 1823 2505
rect 1765 2496 1777 2499
rect 1728 2468 1777 2496
rect 1728 2456 1734 2468
rect 1765 2465 1777 2468
rect 1811 2465 1823 2499
rect 2038 2496 2044 2508
rect 1999 2468 2044 2496
rect 1765 2459 1823 2465
rect 2038 2456 2044 2468
rect 2096 2456 2102 2508
rect 2774 2496 2780 2508
rect 2735 2468 2780 2496
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 1394 2360 1400 2372
rect 1355 2332 1400 2360
rect 1394 2320 1400 2332
rect 1452 2320 1458 2372
rect 2976 2369 3004 2536
rect 4154 2496 4160 2508
rect 4115 2468 4160 2496
rect 4154 2456 4160 2468
rect 4212 2456 4218 2508
rect 4798 2456 4804 2508
rect 4856 2496 4862 2508
rect 4893 2499 4951 2505
rect 4893 2496 4905 2499
rect 4856 2468 4905 2496
rect 4856 2456 4862 2468
rect 4893 2465 4905 2468
rect 4939 2496 4951 2499
rect 5442 2496 5448 2508
rect 4939 2468 5448 2496
rect 4939 2465 4951 2468
rect 4893 2459 4951 2465
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 5721 2499 5779 2505
rect 5721 2496 5733 2499
rect 5592 2468 5733 2496
rect 5592 2456 5598 2468
rect 5721 2465 5733 2468
rect 5767 2465 5779 2499
rect 5721 2459 5779 2465
rect 5828 2428 5856 2536
rect 8573 2533 8585 2567
rect 8619 2564 8631 2567
rect 12986 2564 12992 2576
rect 8619 2536 12992 2564
rect 8619 2533 8631 2536
rect 8573 2527 8631 2533
rect 12986 2524 12992 2536
rect 13044 2564 13050 2576
rect 14200 2564 14228 2592
rect 14660 2573 14688 2604
rect 14918 2592 14924 2604
rect 14976 2632 14982 2644
rect 14976 2604 16574 2632
rect 14976 2592 14982 2604
rect 13044 2536 13492 2564
rect 13044 2524 13050 2536
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 7282 2496 7288 2508
rect 6972 2468 7017 2496
rect 7243 2468 7288 2496
rect 6972 2456 6978 2468
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 8294 2456 8300 2508
rect 8352 2496 8358 2508
rect 8389 2499 8447 2505
rect 8389 2496 8401 2499
rect 8352 2468 8401 2496
rect 8352 2456 8358 2468
rect 8389 2465 8401 2468
rect 8435 2465 8447 2499
rect 8389 2459 8447 2465
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 9861 2499 9919 2505
rect 9861 2496 9873 2499
rect 9732 2468 9873 2496
rect 9732 2456 9738 2468
rect 9861 2465 9873 2468
rect 9907 2465 9919 2499
rect 9861 2459 9919 2465
rect 11054 2456 11060 2508
rect 11112 2496 11118 2508
rect 11241 2499 11299 2505
rect 11241 2496 11253 2499
rect 11112 2468 11253 2496
rect 11112 2456 11118 2468
rect 11241 2465 11253 2468
rect 11287 2465 11299 2499
rect 11241 2459 11299 2465
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 13464 2505 13492 2536
rect 13648 2536 14228 2564
rect 14645 2567 14703 2573
rect 13648 2505 13676 2536
rect 14645 2533 14657 2567
rect 14691 2533 14703 2567
rect 16546 2564 16574 2604
rect 16669 2567 16727 2573
rect 16669 2564 16681 2567
rect 16546 2536 16681 2564
rect 14645 2527 14703 2533
rect 16669 2533 16681 2536
rect 16715 2533 16727 2567
rect 16669 2527 16727 2533
rect 12529 2499 12587 2505
rect 12529 2496 12541 2499
rect 12492 2468 12541 2496
rect 12492 2456 12498 2468
rect 12529 2465 12541 2468
rect 12575 2465 12587 2499
rect 12529 2459 12587 2465
rect 13449 2499 13507 2505
rect 13449 2465 13461 2499
rect 13495 2465 13507 2499
rect 13449 2459 13507 2465
rect 13633 2499 13691 2505
rect 13633 2465 13645 2499
rect 13679 2465 13691 2499
rect 13814 2496 13820 2508
rect 13727 2468 13820 2496
rect 13633 2459 13691 2465
rect 13814 2456 13820 2468
rect 13872 2456 13878 2508
rect 13906 2456 13912 2508
rect 13964 2496 13970 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 13964 2468 14197 2496
rect 13964 2456 13970 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 14185 2459 14243 2465
rect 15562 2456 15568 2508
rect 15620 2456 15626 2508
rect 16945 2499 17003 2505
rect 16945 2465 16957 2499
rect 16991 2496 17003 2499
rect 17034 2496 17040 2508
rect 16991 2468 17040 2496
rect 16991 2465 17003 2468
rect 16945 2459 17003 2465
rect 17034 2456 17040 2468
rect 17092 2456 17098 2508
rect 8662 2428 8668 2440
rect 5828 2400 8668 2428
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 12618 2388 12624 2440
rect 12676 2428 12682 2440
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 12676 2400 12817 2428
rect 12676 2388 12682 2400
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 13832 2428 13860 2456
rect 14001 2431 14059 2437
rect 14001 2428 14013 2431
rect 13832 2400 14013 2428
rect 12805 2391 12863 2397
rect 14001 2397 14013 2400
rect 14047 2397 14059 2431
rect 14001 2391 14059 2397
rect 14829 2431 14887 2437
rect 14829 2397 14841 2431
rect 14875 2428 14887 2431
rect 16574 2428 16580 2440
rect 14875 2400 16580 2428
rect 14875 2397 14887 2400
rect 14829 2391 14887 2397
rect 16574 2388 16580 2400
rect 16632 2388 16638 2440
rect 2961 2363 3019 2369
rect 2961 2329 2973 2363
rect 3007 2329 3019 2363
rect 2961 2323 3019 2329
rect 5077 2363 5135 2369
rect 5077 2329 5089 2363
rect 5123 2360 5135 2363
rect 5258 2360 5264 2372
rect 5123 2332 5264 2360
rect 5123 2329 5135 2332
rect 5077 2323 5135 2329
rect 5258 2320 5264 2332
rect 5316 2320 5322 2372
rect 5626 2360 5632 2372
rect 5368 2332 5632 2360
rect 4341 2295 4399 2301
rect 4341 2261 4353 2295
rect 4387 2292 4399 2295
rect 5368 2292 5396 2332
rect 5626 2320 5632 2332
rect 5684 2320 5690 2372
rect 10962 2320 10968 2372
rect 11020 2360 11026 2372
rect 11057 2363 11115 2369
rect 11057 2360 11069 2363
rect 11020 2332 11069 2360
rect 11020 2320 11026 2332
rect 11057 2329 11069 2332
rect 11103 2329 11115 2363
rect 11057 2323 11115 2329
rect 4387 2264 5396 2292
rect 4387 2261 4399 2264
rect 4341 2255 4399 2261
rect 5442 2252 5448 2304
rect 5500 2292 5506 2304
rect 5537 2295 5595 2301
rect 5537 2292 5549 2295
rect 5500 2264 5549 2292
rect 5500 2252 5506 2264
rect 5537 2261 5549 2264
rect 5583 2261 5595 2295
rect 5537 2255 5595 2261
rect 1104 2202 17296 2224
rect 1104 2150 3680 2202
rect 3732 2150 3744 2202
rect 3796 2150 3808 2202
rect 3860 2150 3872 2202
rect 3924 2150 9078 2202
rect 9130 2150 9142 2202
rect 9194 2150 9206 2202
rect 9258 2150 9270 2202
rect 9322 2150 14475 2202
rect 14527 2150 14539 2202
rect 14591 2150 14603 2202
rect 14655 2150 14667 2202
rect 14719 2150 17296 2202
rect 1104 2128 17296 2150
<< via1 >>
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 6571 17926 6623 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 11904 17926 11956 17978
rect 11968 17926 12020 17978
rect 1492 17867 1544 17876
rect 1492 17833 1501 17867
rect 1501 17833 1535 17867
rect 1535 17833 1544 17867
rect 1492 17824 1544 17833
rect 480 17756 532 17808
rect 1584 17731 1636 17740
rect 1584 17697 1593 17731
rect 1593 17697 1627 17731
rect 1627 17697 1636 17731
rect 1584 17688 1636 17697
rect 1860 17731 1912 17740
rect 1860 17697 1869 17731
rect 1869 17697 1903 17731
rect 1903 17697 1912 17731
rect 1860 17688 1912 17697
rect 3240 17731 3292 17740
rect 3240 17697 3249 17731
rect 3249 17697 3283 17731
rect 3283 17697 3292 17731
rect 3240 17688 3292 17697
rect 4252 17731 4304 17740
rect 4252 17697 4253 17731
rect 4253 17697 4287 17731
rect 4287 17697 4304 17731
rect 4252 17688 4304 17697
rect 4620 17688 4672 17740
rect 6000 17731 6052 17740
rect 6000 17697 6009 17731
rect 6009 17697 6043 17731
rect 6043 17697 6052 17731
rect 6000 17688 6052 17697
rect 7380 17688 7432 17740
rect 8300 17688 8352 17740
rect 16028 17756 16080 17808
rect 17040 17756 17092 17808
rect 8852 17688 8904 17740
rect 10140 17731 10192 17740
rect 10140 17697 10149 17731
rect 10149 17697 10183 17731
rect 10183 17697 10192 17731
rect 10140 17688 10192 17697
rect 11520 17688 11572 17740
rect 12348 17731 12400 17740
rect 12348 17697 12357 17731
rect 12357 17697 12391 17731
rect 12391 17697 12400 17731
rect 12348 17688 12400 17697
rect 12900 17731 12952 17740
rect 12900 17697 12909 17731
rect 12909 17697 12943 17731
rect 12943 17697 12952 17731
rect 12900 17688 12952 17697
rect 14280 17688 14332 17740
rect 13452 17620 13504 17672
rect 15384 17620 15436 17672
rect 7564 17552 7616 17604
rect 8576 17552 8628 17604
rect 2044 17527 2096 17536
rect 2044 17493 2053 17527
rect 2053 17493 2087 17527
rect 2087 17493 2096 17527
rect 2044 17484 2096 17493
rect 2228 17484 2280 17536
rect 3240 17484 3292 17536
rect 4436 17527 4488 17536
rect 4436 17493 4445 17527
rect 4445 17493 4479 17527
rect 4479 17493 4488 17527
rect 4436 17484 4488 17493
rect 4528 17484 4580 17536
rect 7104 17484 7156 17536
rect 8944 17527 8996 17536
rect 8944 17493 8953 17527
rect 8953 17493 8987 17527
rect 8987 17493 8996 17527
rect 8944 17484 8996 17493
rect 9864 17484 9916 17536
rect 10416 17484 10468 17536
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 13176 17484 13228 17536
rect 13912 17484 13964 17536
rect 16304 17484 16356 17536
rect 16856 17484 16908 17536
rect 3680 17382 3732 17434
rect 3744 17382 3796 17434
rect 3808 17382 3860 17434
rect 3872 17382 3924 17434
rect 9078 17382 9130 17434
rect 9142 17382 9194 17434
rect 9206 17382 9258 17434
rect 9270 17382 9322 17434
rect 14475 17382 14527 17434
rect 14539 17382 14591 17434
rect 14603 17382 14655 17434
rect 14667 17382 14719 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 2780 17280 2832 17332
rect 2136 17144 2188 17196
rect 4252 17280 4304 17332
rect 15384 17323 15436 17332
rect 15384 17289 15393 17323
rect 15393 17289 15427 17323
rect 15427 17289 15436 17323
rect 15384 17280 15436 17289
rect 16028 17280 16080 17332
rect 1768 17119 1820 17128
rect 1768 17085 1777 17119
rect 1777 17085 1811 17119
rect 1811 17085 1820 17119
rect 1768 17076 1820 17085
rect 2596 17119 2648 17128
rect 2596 17085 2605 17119
rect 2605 17085 2639 17119
rect 2639 17085 2648 17119
rect 2596 17076 2648 17085
rect 2872 17076 2924 17128
rect 3424 17119 3476 17128
rect 3424 17085 3433 17119
rect 3433 17085 3467 17119
rect 3467 17085 3476 17119
rect 3424 17076 3476 17085
rect 4436 17008 4488 17060
rect 6736 17144 6788 17196
rect 7012 17119 7064 17128
rect 1676 16940 1728 16992
rect 3056 16983 3108 16992
rect 3056 16949 3065 16983
rect 3065 16949 3099 16983
rect 3099 16949 3108 16983
rect 3056 16940 3108 16949
rect 3424 16940 3476 16992
rect 6276 16940 6328 16992
rect 7012 17085 7021 17119
rect 7021 17085 7055 17119
rect 7055 17085 7064 17119
rect 7012 17076 7064 17085
rect 8024 17119 8076 17128
rect 8024 17085 8033 17119
rect 8033 17085 8067 17119
rect 8067 17085 8076 17119
rect 8024 17076 8076 17085
rect 10968 17212 11020 17264
rect 15660 17212 15712 17264
rect 13912 17187 13964 17196
rect 13912 17153 13921 17187
rect 13921 17153 13955 17187
rect 13955 17153 13964 17187
rect 13912 17144 13964 17153
rect 10324 17119 10376 17128
rect 10324 17085 10333 17119
rect 10333 17085 10367 17119
rect 10367 17085 10376 17119
rect 10324 17076 10376 17085
rect 10508 17119 10560 17128
rect 10508 17085 10517 17119
rect 10517 17085 10551 17119
rect 10551 17085 10560 17119
rect 10508 17076 10560 17085
rect 11428 17076 11480 17128
rect 13452 17076 13504 17128
rect 15568 17076 15620 17128
rect 15752 17119 15804 17128
rect 15752 17085 15761 17119
rect 15761 17085 15795 17119
rect 15795 17085 15804 17119
rect 15752 17076 15804 17085
rect 17040 17076 17092 17128
rect 7288 17008 7340 17060
rect 8944 17008 8996 17060
rect 6828 16940 6880 16992
rect 11520 17008 11572 17060
rect 12532 17008 12584 17060
rect 14556 17008 14608 17060
rect 16764 17051 16816 17060
rect 16764 17017 16773 17051
rect 16773 17017 16807 17051
rect 16807 17017 16816 17051
rect 16764 17008 16816 17017
rect 10600 16940 10652 16992
rect 12624 16940 12676 16992
rect 15476 16983 15528 16992
rect 15476 16949 15485 16983
rect 15485 16949 15519 16983
rect 15519 16949 15528 16983
rect 15476 16940 15528 16949
rect 15568 16940 15620 16992
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 6571 16838 6623 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 11904 16838 11956 16890
rect 11968 16838 12020 16890
rect 2596 16736 2648 16788
rect 4252 16736 4304 16788
rect 1676 16711 1728 16720
rect 1676 16677 1685 16711
rect 1685 16677 1719 16711
rect 1719 16677 1728 16711
rect 1676 16668 1728 16677
rect 3056 16668 3108 16720
rect 3424 16643 3476 16652
rect 3424 16609 3433 16643
rect 3433 16609 3467 16643
rect 3467 16609 3476 16643
rect 3424 16600 3476 16609
rect 5448 16736 5500 16788
rect 7840 16736 7892 16788
rect 14556 16779 14608 16788
rect 6276 16668 6328 16720
rect 9956 16668 10008 16720
rect 10324 16711 10376 16720
rect 10324 16677 10333 16711
rect 10333 16677 10367 16711
rect 10367 16677 10376 16711
rect 14556 16745 14565 16779
rect 14565 16745 14599 16779
rect 14599 16745 14608 16779
rect 14556 16736 14608 16745
rect 10324 16668 10376 16677
rect 7840 16600 7892 16652
rect 8300 16643 8352 16652
rect 8300 16609 8309 16643
rect 8309 16609 8343 16643
rect 8343 16609 8352 16643
rect 8300 16600 8352 16609
rect 1768 16532 1820 16584
rect 3516 16532 3568 16584
rect 8024 16532 8076 16584
rect 10600 16600 10652 16652
rect 11428 16643 11480 16652
rect 10140 16532 10192 16584
rect 3424 16396 3476 16448
rect 4804 16439 4856 16448
rect 4804 16405 4813 16439
rect 4813 16405 4847 16439
rect 4847 16405 4856 16439
rect 4804 16396 4856 16405
rect 7288 16396 7340 16448
rect 10692 16396 10744 16448
rect 11428 16609 11437 16643
rect 11437 16609 11471 16643
rect 11471 16609 11480 16643
rect 11428 16600 11480 16609
rect 11520 16600 11572 16652
rect 12256 16600 12308 16652
rect 12348 16600 12400 16652
rect 13360 16600 13412 16652
rect 15752 16600 15804 16652
rect 16028 16643 16080 16652
rect 16028 16609 16037 16643
rect 16037 16609 16071 16643
rect 16071 16609 16080 16643
rect 16028 16600 16080 16609
rect 16304 16600 16356 16652
rect 16764 16643 16816 16652
rect 16764 16609 16773 16643
rect 16773 16609 16807 16643
rect 16807 16609 16816 16643
rect 16764 16600 16816 16609
rect 11612 16532 11664 16584
rect 12624 16396 12676 16448
rect 15384 16396 15436 16448
rect 3680 16294 3732 16346
rect 3744 16294 3796 16346
rect 3808 16294 3860 16346
rect 3872 16294 3924 16346
rect 9078 16294 9130 16346
rect 9142 16294 9194 16346
rect 9206 16294 9258 16346
rect 9270 16294 9322 16346
rect 14475 16294 14527 16346
rect 14539 16294 14591 16346
rect 14603 16294 14655 16346
rect 14667 16294 14719 16346
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 3516 15988 3568 16040
rect 7012 16192 7064 16244
rect 16764 16235 16816 16244
rect 16764 16201 16773 16235
rect 16773 16201 16807 16235
rect 16807 16201 16816 16235
rect 16764 16192 16816 16201
rect 7288 16124 7340 16176
rect 6460 15988 6512 16040
rect 6736 16056 6788 16108
rect 7012 16031 7064 16040
rect 4436 15920 4488 15972
rect 4804 15920 4856 15972
rect 7012 15997 7021 16031
rect 7021 15997 7055 16031
rect 7055 15997 7064 16031
rect 7012 15988 7064 15997
rect 7288 16031 7340 16040
rect 7288 15997 7297 16031
rect 7297 15997 7331 16031
rect 7331 15997 7340 16031
rect 10416 16124 10468 16176
rect 10692 16056 10744 16108
rect 13452 16056 13504 16108
rect 16028 16056 16080 16108
rect 7288 15988 7340 15997
rect 9956 16031 10008 16040
rect 9956 15997 9965 16031
rect 9965 15997 9999 16031
rect 9999 15997 10008 16031
rect 9956 15988 10008 15997
rect 10140 16031 10192 16040
rect 10140 15997 10149 16031
rect 10149 15997 10183 16031
rect 10183 15997 10192 16031
rect 10140 15988 10192 15997
rect 10416 15988 10468 16040
rect 12440 16031 12492 16040
rect 4896 15852 4948 15904
rect 8392 15920 8444 15972
rect 8852 15852 8904 15904
rect 9772 15895 9824 15904
rect 9772 15861 9781 15895
rect 9781 15861 9815 15895
rect 9815 15861 9824 15895
rect 9772 15852 9824 15861
rect 10048 15852 10100 15904
rect 10600 15920 10652 15972
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 13452 15920 13504 15972
rect 16028 15920 16080 15972
rect 12900 15852 12952 15904
rect 12992 15852 13044 15904
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 6571 15750 6623 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 11904 15750 11956 15802
rect 11968 15750 12020 15802
rect 3516 15648 3568 15700
rect 10048 15691 10100 15700
rect 10048 15657 10057 15691
rect 10057 15657 10091 15691
rect 10091 15657 10100 15691
rect 10048 15648 10100 15657
rect 2964 15580 3016 15632
rect 2136 15555 2188 15564
rect 2136 15521 2145 15555
rect 2145 15521 2179 15555
rect 2179 15521 2188 15555
rect 2136 15512 2188 15521
rect 3148 15512 3200 15564
rect 3332 15555 3384 15564
rect 3332 15521 3341 15555
rect 3341 15521 3375 15555
rect 3375 15521 3384 15555
rect 3332 15512 3384 15521
rect 4712 15512 4764 15564
rect 8852 15623 8904 15632
rect 8852 15589 8861 15623
rect 8861 15589 8895 15623
rect 8895 15589 8904 15623
rect 8852 15580 8904 15589
rect 10692 15580 10744 15632
rect 7196 15555 7248 15564
rect 7196 15521 7205 15555
rect 7205 15521 7239 15555
rect 7239 15521 7248 15555
rect 7196 15512 7248 15521
rect 7564 15555 7616 15564
rect 7564 15521 7573 15555
rect 7573 15521 7607 15555
rect 7607 15521 7616 15555
rect 7564 15512 7616 15521
rect 8392 15555 8444 15564
rect 8392 15521 8401 15555
rect 8401 15521 8435 15555
rect 8435 15521 8444 15555
rect 8392 15512 8444 15521
rect 9772 15512 9824 15564
rect 10600 15512 10652 15564
rect 11980 15555 12032 15564
rect 11980 15521 11989 15555
rect 11989 15521 12023 15555
rect 12023 15521 12032 15555
rect 11980 15512 12032 15521
rect 4344 15444 4396 15496
rect 7288 15487 7340 15496
rect 7288 15453 7297 15487
rect 7297 15453 7331 15487
rect 7331 15453 7340 15487
rect 7288 15444 7340 15453
rect 7840 15444 7892 15496
rect 8116 15444 8168 15496
rect 3424 15376 3476 15428
rect 4068 15376 4120 15428
rect 12072 15444 12124 15496
rect 9496 15376 9548 15428
rect 12256 15555 12308 15564
rect 12256 15521 12265 15555
rect 12265 15521 12299 15555
rect 12299 15521 12308 15555
rect 12992 15648 13044 15700
rect 13452 15648 13504 15700
rect 16028 15648 16080 15700
rect 12256 15512 12308 15521
rect 12348 15487 12400 15496
rect 12348 15453 12357 15487
rect 12357 15453 12391 15487
rect 12391 15453 12400 15487
rect 12348 15444 12400 15453
rect 12808 15555 12860 15564
rect 12808 15521 12817 15555
rect 12817 15521 12851 15555
rect 12851 15521 12860 15555
rect 12992 15555 13044 15564
rect 12808 15512 12860 15521
rect 12992 15521 13001 15555
rect 13001 15521 13035 15555
rect 13035 15521 13044 15555
rect 12992 15512 13044 15521
rect 13360 15555 13412 15564
rect 13360 15521 13369 15555
rect 13369 15521 13403 15555
rect 13403 15521 13412 15555
rect 13360 15512 13412 15521
rect 15292 15512 15344 15564
rect 15752 15512 15804 15564
rect 16488 15512 16540 15564
rect 12624 15376 12676 15428
rect 1860 15308 1912 15360
rect 4160 15308 4212 15360
rect 8484 15308 8536 15360
rect 12900 15308 12952 15360
rect 13820 15308 13872 15360
rect 3680 15206 3732 15258
rect 3744 15206 3796 15258
rect 3808 15206 3860 15258
rect 3872 15206 3924 15258
rect 9078 15206 9130 15258
rect 9142 15206 9194 15258
rect 9206 15206 9258 15258
rect 9270 15206 9322 15258
rect 14475 15206 14527 15258
rect 14539 15206 14591 15258
rect 14603 15206 14655 15258
rect 14667 15206 14719 15258
rect 3148 15104 3200 15156
rect 4436 15104 4488 15156
rect 7288 15104 7340 15156
rect 3332 15036 3384 15088
rect 4252 15036 4304 15088
rect 6828 15036 6880 15088
rect 10968 15104 11020 15156
rect 12348 15104 12400 15156
rect 12808 15104 12860 15156
rect 14372 15104 14424 15156
rect 15016 15104 15068 15156
rect 15292 15104 15344 15156
rect 3332 14900 3384 14952
rect 3700 14943 3752 14952
rect 3700 14909 3735 14943
rect 3735 14909 3752 14943
rect 3884 14943 3936 14952
rect 3700 14900 3752 14909
rect 3884 14909 3893 14943
rect 3893 14909 3927 14943
rect 3927 14909 3936 14943
rect 3884 14900 3936 14909
rect 1860 14832 1912 14884
rect 3516 14875 3568 14884
rect 3516 14841 3525 14875
rect 3525 14841 3559 14875
rect 3559 14841 3568 14875
rect 3516 14832 3568 14841
rect 2780 14764 2832 14816
rect 4068 14832 4120 14884
rect 3700 14764 3752 14816
rect 4344 14968 4396 15020
rect 5448 14943 5500 14952
rect 5448 14909 5457 14943
rect 5457 14909 5491 14943
rect 5491 14909 5500 14943
rect 5448 14900 5500 14909
rect 7196 14968 7248 15020
rect 9496 15011 9548 15020
rect 7012 14875 7064 14884
rect 7012 14841 7021 14875
rect 7021 14841 7055 14875
rect 7055 14841 7064 14875
rect 7012 14832 7064 14841
rect 8116 14900 8168 14952
rect 8484 14943 8536 14952
rect 8484 14909 8493 14943
rect 8493 14909 8527 14943
rect 8527 14909 8536 14943
rect 8484 14900 8536 14909
rect 8668 14943 8720 14952
rect 8668 14909 8677 14943
rect 8677 14909 8711 14943
rect 8711 14909 8720 14943
rect 8668 14900 8720 14909
rect 8852 14943 8904 14952
rect 8852 14909 8861 14943
rect 8861 14909 8895 14943
rect 8895 14909 8904 14943
rect 8852 14900 8904 14909
rect 9496 14977 9505 15011
rect 9505 14977 9539 15011
rect 9539 14977 9548 15011
rect 9496 14968 9548 14977
rect 13820 14968 13872 15020
rect 14924 15036 14976 15088
rect 15016 15011 15068 15020
rect 15016 14977 15025 15011
rect 15025 14977 15059 15011
rect 15059 14977 15068 15011
rect 15016 14968 15068 14977
rect 7564 14832 7616 14884
rect 10508 14900 10560 14952
rect 10692 14900 10744 14952
rect 10876 14943 10928 14952
rect 10876 14909 10885 14943
rect 10885 14909 10919 14943
rect 10919 14909 10928 14943
rect 10876 14900 10928 14909
rect 10968 14943 11020 14952
rect 10968 14909 10977 14943
rect 10977 14909 11011 14943
rect 11011 14909 11020 14943
rect 10968 14900 11020 14909
rect 12256 14900 12308 14952
rect 5540 14764 5592 14816
rect 6828 14764 6880 14816
rect 10508 14764 10560 14816
rect 12072 14832 12124 14884
rect 14372 14900 14424 14952
rect 14924 14943 14976 14952
rect 14924 14909 14933 14943
rect 14933 14909 14967 14943
rect 14967 14909 14976 14943
rect 15108 14943 15160 14952
rect 14924 14900 14976 14909
rect 15108 14909 15117 14943
rect 15117 14909 15151 14943
rect 15151 14909 15160 14943
rect 15108 14900 15160 14909
rect 15292 14943 15344 14952
rect 15292 14909 15301 14943
rect 15301 14909 15335 14943
rect 15335 14909 15344 14943
rect 15292 14900 15344 14909
rect 15568 14943 15620 14952
rect 15568 14909 15577 14943
rect 15577 14909 15611 14943
rect 15611 14909 15620 14943
rect 15568 14900 15620 14909
rect 16764 14943 16816 14952
rect 16764 14909 16773 14943
rect 16773 14909 16807 14943
rect 16807 14909 16816 14943
rect 16764 14900 16816 14909
rect 10968 14764 11020 14816
rect 12164 14764 12216 14816
rect 15108 14764 15160 14816
rect 16672 14764 16724 14816
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 6571 14662 6623 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 11904 14662 11956 14714
rect 11968 14662 12020 14714
rect 3332 14603 3384 14612
rect 3332 14569 3341 14603
rect 3341 14569 3375 14603
rect 3375 14569 3384 14603
rect 3332 14560 3384 14569
rect 4252 14560 4304 14612
rect 2964 14535 3016 14544
rect 2964 14501 2973 14535
rect 2973 14501 3007 14535
rect 3007 14501 3016 14535
rect 2964 14492 3016 14501
rect 3424 14492 3476 14544
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 3332 14424 3384 14476
rect 4436 14492 4488 14544
rect 3700 14467 3752 14476
rect 3700 14433 3709 14467
rect 3709 14433 3743 14467
rect 3743 14433 3752 14467
rect 3700 14424 3752 14433
rect 3516 14356 3568 14408
rect 4160 14424 4212 14476
rect 4344 14424 4396 14476
rect 5540 14492 5592 14544
rect 5264 14356 5316 14408
rect 7288 14560 7340 14612
rect 10784 14560 10836 14612
rect 7012 14492 7064 14544
rect 12440 14560 12492 14612
rect 7840 14467 7892 14476
rect 7840 14433 7849 14467
rect 7849 14433 7883 14467
rect 7883 14433 7892 14467
rect 7840 14424 7892 14433
rect 10508 14467 10560 14476
rect 10508 14433 10518 14467
rect 10518 14433 10560 14467
rect 10508 14424 10560 14433
rect 10324 14356 10376 14408
rect 10692 14356 10744 14408
rect 11612 14492 11664 14544
rect 12164 14535 12216 14544
rect 12164 14501 12173 14535
rect 12173 14501 12207 14535
rect 12207 14501 12216 14535
rect 12164 14492 12216 14501
rect 12992 14492 13044 14544
rect 12532 14424 12584 14476
rect 12716 14467 12768 14476
rect 12716 14433 12725 14467
rect 12725 14433 12759 14467
rect 12759 14433 12768 14467
rect 12716 14424 12768 14433
rect 12808 14467 12860 14476
rect 12808 14433 12817 14467
rect 12817 14433 12851 14467
rect 12851 14433 12860 14467
rect 14096 14492 14148 14544
rect 15568 14492 15620 14544
rect 12808 14424 12860 14433
rect 15384 14424 15436 14476
rect 8024 14288 8076 14340
rect 9404 14288 9456 14340
rect 10416 14288 10468 14340
rect 10600 14331 10652 14340
rect 10600 14297 10609 14331
rect 10609 14297 10643 14331
rect 10643 14297 10652 14331
rect 10600 14288 10652 14297
rect 14280 14356 14332 14408
rect 13360 14288 13412 14340
rect 1860 14220 1912 14272
rect 3516 14263 3568 14272
rect 3516 14229 3525 14263
rect 3525 14229 3559 14263
rect 3559 14229 3568 14263
rect 3516 14220 3568 14229
rect 5816 14220 5868 14272
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 12624 14220 12676 14272
rect 15292 14220 15344 14272
rect 3680 14118 3732 14170
rect 3744 14118 3796 14170
rect 3808 14118 3860 14170
rect 3872 14118 3924 14170
rect 9078 14118 9130 14170
rect 9142 14118 9194 14170
rect 9206 14118 9258 14170
rect 9270 14118 9322 14170
rect 14475 14118 14527 14170
rect 14539 14118 14591 14170
rect 14603 14118 14655 14170
rect 14667 14118 14719 14170
rect 5264 14059 5316 14068
rect 5264 14025 5273 14059
rect 5273 14025 5307 14059
rect 5307 14025 5316 14059
rect 5264 14016 5316 14025
rect 8116 14059 8168 14068
rect 8116 14025 8125 14059
rect 8125 14025 8159 14059
rect 8159 14025 8168 14059
rect 8116 14016 8168 14025
rect 8852 14059 8904 14068
rect 8852 14025 8861 14059
rect 8861 14025 8895 14059
rect 8895 14025 8904 14059
rect 8852 14016 8904 14025
rect 10416 14016 10468 14068
rect 2320 13948 2372 14000
rect 3516 13812 3568 13864
rect 4712 13812 4764 13864
rect 5908 13855 5960 13864
rect 5908 13821 5917 13855
rect 5917 13821 5951 13855
rect 5951 13821 5960 13855
rect 5908 13812 5960 13821
rect 6000 13855 6052 13864
rect 6000 13821 6009 13855
rect 6009 13821 6043 13855
rect 6043 13821 6052 13855
rect 6000 13812 6052 13821
rect 10324 13948 10376 14000
rect 9956 13923 10008 13932
rect 9956 13889 9965 13923
rect 9965 13889 9999 13923
rect 9999 13889 10008 13923
rect 9956 13880 10008 13889
rect 13360 14016 13412 14068
rect 14096 14059 14148 14068
rect 12624 13923 12676 13932
rect 12624 13889 12633 13923
rect 12633 13889 12667 13923
rect 12667 13889 12676 13923
rect 12624 13880 12676 13889
rect 14096 14025 14105 14059
rect 14105 14025 14139 14059
rect 14139 14025 14148 14059
rect 14096 14016 14148 14025
rect 14372 14016 14424 14068
rect 14372 13880 14424 13932
rect 15292 13923 15344 13932
rect 15292 13889 15301 13923
rect 15301 13889 15335 13923
rect 15335 13889 15344 13923
rect 15292 13880 15344 13889
rect 15660 13880 15712 13932
rect 5540 13787 5592 13796
rect 5540 13753 5549 13787
rect 5549 13753 5583 13787
rect 5583 13753 5592 13787
rect 5540 13744 5592 13753
rect 3424 13676 3476 13728
rect 4068 13676 4120 13728
rect 4436 13676 4488 13728
rect 5816 13744 5868 13796
rect 10048 13855 10100 13864
rect 10048 13821 10057 13855
rect 10057 13821 10091 13855
rect 10091 13821 10100 13855
rect 10324 13855 10376 13864
rect 10048 13812 10100 13821
rect 10324 13821 10333 13855
rect 10333 13821 10367 13855
rect 10367 13821 10376 13855
rect 10324 13812 10376 13821
rect 10784 13812 10836 13864
rect 14924 13855 14976 13864
rect 10968 13744 11020 13796
rect 12900 13744 12952 13796
rect 13360 13744 13412 13796
rect 14924 13821 14933 13855
rect 14933 13821 14967 13855
rect 14967 13821 14976 13855
rect 14924 13812 14976 13821
rect 15384 13744 15436 13796
rect 16304 13744 16356 13796
rect 6000 13676 6052 13728
rect 9956 13676 10008 13728
rect 14280 13676 14332 13728
rect 14740 13676 14792 13728
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 6571 13574 6623 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 11904 13574 11956 13626
rect 11968 13574 12020 13626
rect 4252 13472 4304 13524
rect 5448 13472 5500 13524
rect 5540 13472 5592 13524
rect 3516 13447 3568 13456
rect 3516 13413 3525 13447
rect 3525 13413 3559 13447
rect 3559 13413 3568 13447
rect 3516 13404 3568 13413
rect 4712 13447 4764 13456
rect 2136 13336 2188 13388
rect 4068 13379 4120 13388
rect 1952 13132 2004 13184
rect 3516 13132 3568 13184
rect 4068 13345 4077 13379
rect 4077 13345 4111 13379
rect 4111 13345 4120 13379
rect 4068 13336 4120 13345
rect 4712 13413 4721 13447
rect 4721 13413 4755 13447
rect 4755 13413 4764 13447
rect 4712 13404 4764 13413
rect 4252 13336 4304 13388
rect 4896 13379 4948 13388
rect 4896 13345 4905 13379
rect 4905 13345 4939 13379
rect 4939 13345 4948 13379
rect 4896 13336 4948 13345
rect 6000 13379 6052 13388
rect 6000 13345 6009 13379
rect 6009 13345 6043 13379
rect 6043 13345 6052 13379
rect 6000 13336 6052 13345
rect 6092 13336 6144 13388
rect 4344 13311 4396 13320
rect 4344 13277 4353 13311
rect 4353 13277 4387 13311
rect 4387 13277 4396 13311
rect 4344 13268 4396 13277
rect 3976 13200 4028 13252
rect 7840 13472 7892 13524
rect 12716 13472 12768 13524
rect 13360 13472 13412 13524
rect 16304 13515 16356 13524
rect 16304 13481 16313 13515
rect 16313 13481 16347 13515
rect 16347 13481 16356 13515
rect 16304 13472 16356 13481
rect 12256 13404 12308 13456
rect 13544 13404 13596 13456
rect 15200 13404 15252 13456
rect 6736 13379 6788 13388
rect 6736 13345 6745 13379
rect 6745 13345 6779 13379
rect 6779 13345 6788 13379
rect 6736 13336 6788 13345
rect 7472 13336 7524 13388
rect 7656 13379 7708 13388
rect 7656 13345 7665 13379
rect 7665 13345 7699 13379
rect 7699 13345 7708 13379
rect 7656 13336 7708 13345
rect 11428 13336 11480 13388
rect 6552 13200 6604 13252
rect 4068 13132 4120 13184
rect 4252 13132 4304 13184
rect 4620 13132 4672 13184
rect 4988 13132 5040 13184
rect 5908 13132 5960 13184
rect 6184 13132 6236 13184
rect 6828 13268 6880 13320
rect 12900 13336 12952 13388
rect 13268 13379 13320 13388
rect 13268 13345 13277 13379
rect 13277 13345 13311 13379
rect 13311 13345 13320 13379
rect 13268 13336 13320 13345
rect 14740 13336 14792 13388
rect 15016 13336 15068 13388
rect 15568 13379 15620 13388
rect 15568 13345 15577 13379
rect 15577 13345 15611 13379
rect 15611 13345 15620 13379
rect 15568 13336 15620 13345
rect 16212 13336 16264 13388
rect 16488 13379 16540 13388
rect 16488 13345 16497 13379
rect 16497 13345 16531 13379
rect 16531 13345 16540 13379
rect 16488 13336 16540 13345
rect 13636 13268 13688 13320
rect 15384 13268 15436 13320
rect 7380 13200 7432 13252
rect 12992 13200 13044 13252
rect 7564 13132 7616 13184
rect 11244 13132 11296 13184
rect 12716 13132 12768 13184
rect 3680 13030 3732 13082
rect 3744 13030 3796 13082
rect 3808 13030 3860 13082
rect 3872 13030 3924 13082
rect 9078 13030 9130 13082
rect 9142 13030 9194 13082
rect 9206 13030 9258 13082
rect 9270 13030 9322 13082
rect 14475 13030 14527 13082
rect 14539 13030 14591 13082
rect 14603 13030 14655 13082
rect 14667 13030 14719 13082
rect 3332 12792 3384 12844
rect 3516 12767 3568 12776
rect 3516 12733 3525 12767
rect 3525 12733 3559 12767
rect 3559 12733 3568 12767
rect 3516 12724 3568 12733
rect 3976 12860 4028 12912
rect 4252 12792 4304 12844
rect 4068 12767 4120 12776
rect 4068 12733 4077 12767
rect 4077 12733 4111 12767
rect 4111 12733 4120 12767
rect 4068 12724 4120 12733
rect 4344 12724 4396 12776
rect 7012 12928 7064 12980
rect 10048 12928 10100 12980
rect 11244 12971 11296 12980
rect 11244 12937 11253 12971
rect 11253 12937 11287 12971
rect 11287 12937 11296 12971
rect 11244 12928 11296 12937
rect 11428 12928 11480 12980
rect 12900 12971 12952 12980
rect 12900 12937 12909 12971
rect 12909 12937 12943 12971
rect 12943 12937 12952 12971
rect 12900 12928 12952 12937
rect 14280 12928 14332 12980
rect 14832 12928 14884 12980
rect 15108 12928 15160 12980
rect 4620 12860 4672 12912
rect 6552 12860 6604 12912
rect 6828 12860 6880 12912
rect 4712 12835 4764 12844
rect 4712 12801 4721 12835
rect 4721 12801 4755 12835
rect 4755 12801 4764 12835
rect 4712 12792 4764 12801
rect 6276 12792 6328 12844
rect 6736 12792 6788 12844
rect 4896 12767 4948 12776
rect 4896 12733 4905 12767
rect 4905 12733 4939 12767
rect 4939 12733 4948 12767
rect 4896 12724 4948 12733
rect 5448 12724 5500 12776
rect 11520 12860 11572 12912
rect 8116 12835 8168 12844
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 8116 12792 8168 12801
rect 9312 12792 9364 12844
rect 7196 12767 7248 12776
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 7380 12767 7432 12776
rect 7380 12733 7387 12767
rect 7387 12733 7432 12767
rect 7380 12724 7432 12733
rect 7564 12767 7616 12776
rect 7564 12733 7573 12767
rect 7573 12733 7607 12767
rect 7607 12733 7616 12767
rect 7564 12724 7616 12733
rect 7656 12767 7708 12776
rect 7656 12733 7670 12767
rect 7670 12733 7704 12767
rect 7704 12733 7708 12767
rect 8208 12767 8260 12776
rect 7656 12724 7708 12733
rect 8208 12733 8217 12767
rect 8217 12733 8251 12767
rect 8251 12733 8260 12767
rect 8208 12724 8260 12733
rect 9680 12724 9732 12776
rect 12072 12767 12124 12776
rect 1952 12656 2004 12708
rect 3424 12656 3476 12708
rect 3884 12656 3936 12708
rect 5816 12656 5868 12708
rect 7472 12699 7524 12708
rect 7472 12665 7481 12699
rect 7481 12665 7515 12699
rect 7515 12665 7524 12699
rect 7472 12656 7524 12665
rect 12072 12733 12081 12767
rect 12081 12733 12115 12767
rect 12115 12733 12124 12767
rect 12072 12724 12124 12733
rect 12992 12767 13044 12776
rect 6000 12588 6052 12640
rect 6828 12588 6880 12640
rect 9404 12588 9456 12640
rect 12992 12733 13001 12767
rect 13001 12733 13035 12767
rect 13035 12733 13044 12767
rect 12992 12724 13044 12733
rect 14096 12724 14148 12776
rect 15200 12767 15252 12776
rect 15200 12733 15209 12767
rect 15209 12733 15243 12767
rect 15243 12733 15252 12767
rect 15200 12724 15252 12733
rect 15384 12724 15436 12776
rect 16764 12767 16816 12776
rect 16764 12733 16773 12767
rect 16773 12733 16807 12767
rect 16807 12733 16816 12767
rect 16764 12724 16816 12733
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 6571 12486 6623 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 11904 12486 11956 12538
rect 11968 12486 12020 12538
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 4160 12291 4212 12300
rect 4160 12257 4169 12291
rect 4169 12257 4203 12291
rect 4203 12257 4212 12291
rect 4160 12248 4212 12257
rect 4252 12291 4304 12300
rect 4252 12257 4261 12291
rect 4261 12257 4295 12291
rect 4295 12257 4304 12291
rect 6736 12316 6788 12368
rect 7288 12427 7340 12436
rect 7288 12393 7297 12427
rect 7297 12393 7331 12427
rect 7331 12393 7340 12427
rect 7288 12384 7340 12393
rect 7472 12384 7524 12436
rect 8208 12384 8260 12436
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 12992 12427 13044 12436
rect 12992 12393 13001 12427
rect 13001 12393 13035 12427
rect 13035 12393 13044 12427
rect 12992 12384 13044 12393
rect 13636 12384 13688 12436
rect 4252 12248 4304 12257
rect 6828 12291 6880 12300
rect 6828 12257 6837 12291
rect 6837 12257 6871 12291
rect 6871 12257 6880 12291
rect 6828 12248 6880 12257
rect 7288 12248 7340 12300
rect 9588 12316 9640 12368
rect 11244 12316 11296 12368
rect 3976 12180 4028 12232
rect 4344 12180 4396 12232
rect 5540 12180 5592 12232
rect 6184 12180 6236 12232
rect 7380 12180 7432 12232
rect 8208 12248 8260 12300
rect 9404 12291 9456 12300
rect 9404 12257 9413 12291
rect 9413 12257 9447 12291
rect 9447 12257 9456 12291
rect 9404 12248 9456 12257
rect 9496 12248 9548 12300
rect 13360 12291 13412 12300
rect 13360 12257 13369 12291
rect 13369 12257 13403 12291
rect 13403 12257 13412 12291
rect 13360 12248 13412 12257
rect 14096 12316 14148 12368
rect 15384 12359 15436 12368
rect 15384 12325 15393 12359
rect 15393 12325 15427 12359
rect 15427 12325 15436 12359
rect 15384 12316 15436 12325
rect 15200 12291 15252 12300
rect 7288 12112 7340 12164
rect 9404 12112 9456 12164
rect 11060 12180 11112 12232
rect 14280 12180 14332 12232
rect 15200 12257 15209 12291
rect 15209 12257 15243 12291
rect 15243 12257 15252 12291
rect 15200 12248 15252 12257
rect 15476 12291 15528 12300
rect 15476 12257 15485 12291
rect 15485 12257 15519 12291
rect 15519 12257 15528 12291
rect 15476 12248 15528 12257
rect 15660 12248 15712 12300
rect 1584 12087 1636 12096
rect 1584 12053 1593 12087
rect 1593 12053 1627 12087
rect 1627 12053 1636 12087
rect 1584 12044 1636 12053
rect 4712 12044 4764 12096
rect 7012 12087 7064 12096
rect 7012 12053 7021 12087
rect 7021 12053 7055 12087
rect 7055 12053 7064 12087
rect 7012 12044 7064 12053
rect 7472 12044 7524 12096
rect 11336 12044 11388 12096
rect 12072 12087 12124 12096
rect 12072 12053 12081 12087
rect 12081 12053 12115 12087
rect 12115 12053 12124 12087
rect 12072 12044 12124 12053
rect 13912 12112 13964 12164
rect 13452 12044 13504 12096
rect 13728 12044 13780 12096
rect 3680 11942 3732 11994
rect 3744 11942 3796 11994
rect 3808 11942 3860 11994
rect 3872 11942 3924 11994
rect 9078 11942 9130 11994
rect 9142 11942 9194 11994
rect 9206 11942 9258 11994
rect 9270 11942 9322 11994
rect 14475 11942 14527 11994
rect 14539 11942 14591 11994
rect 14603 11942 14655 11994
rect 14667 11942 14719 11994
rect 4436 11840 4488 11892
rect 8116 11840 8168 11892
rect 13360 11883 13412 11892
rect 5080 11772 5132 11824
rect 12992 11772 13044 11824
rect 13360 11849 13369 11883
rect 13369 11849 13403 11883
rect 13403 11849 13412 11883
rect 13360 11840 13412 11849
rect 15200 11840 15252 11892
rect 4252 11636 4304 11688
rect 4620 11679 4672 11688
rect 4620 11645 4629 11679
rect 4629 11645 4663 11679
rect 4663 11645 4672 11679
rect 4620 11636 4672 11645
rect 4712 11679 4764 11688
rect 4712 11645 4757 11679
rect 4757 11645 4764 11679
rect 4712 11636 4764 11645
rect 4988 11636 5040 11688
rect 5172 11679 5224 11688
rect 5172 11645 5181 11679
rect 5181 11645 5215 11679
rect 5215 11645 5224 11679
rect 5172 11636 5224 11645
rect 6828 11679 6880 11688
rect 6828 11645 6838 11679
rect 6838 11645 6872 11679
rect 6872 11645 6880 11679
rect 7012 11679 7064 11688
rect 6828 11636 6880 11645
rect 7012 11645 7021 11679
rect 7021 11645 7055 11679
rect 7055 11645 7064 11679
rect 7012 11636 7064 11645
rect 7196 11679 7248 11688
rect 12256 11704 12308 11756
rect 7196 11645 7210 11679
rect 7210 11645 7244 11679
rect 7244 11645 7248 11679
rect 7196 11636 7248 11645
rect 9496 11679 9548 11688
rect 9496 11645 9505 11679
rect 9505 11645 9539 11679
rect 9539 11645 9548 11679
rect 9496 11636 9548 11645
rect 11612 11636 11664 11688
rect 12716 11679 12768 11688
rect 12716 11645 12725 11679
rect 12725 11645 12759 11679
rect 12759 11645 12768 11679
rect 12716 11636 12768 11645
rect 13452 11704 13504 11756
rect 14004 11704 14056 11756
rect 15476 11704 15528 11756
rect 13544 11679 13596 11688
rect 4436 11500 4488 11552
rect 11520 11568 11572 11620
rect 13544 11645 13553 11679
rect 13553 11645 13587 11679
rect 13587 11645 13596 11679
rect 13544 11636 13596 11645
rect 13728 11679 13780 11688
rect 13728 11645 13737 11679
rect 13737 11645 13771 11679
rect 13771 11645 13780 11679
rect 13728 11636 13780 11645
rect 13912 11679 13964 11688
rect 13912 11645 13921 11679
rect 13921 11645 13955 11679
rect 13955 11645 13964 11679
rect 13912 11636 13964 11645
rect 14096 11679 14148 11688
rect 14096 11645 14105 11679
rect 14105 11645 14139 11679
rect 14139 11645 14148 11679
rect 14096 11636 14148 11645
rect 13360 11568 13412 11620
rect 7748 11500 7800 11552
rect 9680 11543 9732 11552
rect 9680 11509 9689 11543
rect 9689 11509 9723 11543
rect 9723 11509 9732 11543
rect 9680 11500 9732 11509
rect 13728 11500 13780 11552
rect 14096 11500 14148 11552
rect 14832 11500 14884 11552
rect 15660 11568 15712 11620
rect 16028 11679 16080 11688
rect 16028 11645 16037 11679
rect 16037 11645 16071 11679
rect 16071 11645 16080 11679
rect 16028 11636 16080 11645
rect 16396 11636 16448 11688
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 6571 11398 6623 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 11904 11398 11956 11450
rect 11968 11398 12020 11450
rect 2688 11296 2740 11348
rect 5172 11339 5224 11348
rect 5172 11305 5181 11339
rect 5181 11305 5215 11339
rect 5215 11305 5224 11339
rect 5172 11296 5224 11305
rect 6828 11339 6880 11348
rect 6828 11305 6837 11339
rect 6837 11305 6871 11339
rect 6871 11305 6880 11339
rect 6828 11296 6880 11305
rect 2044 11203 2096 11212
rect 2044 11169 2053 11203
rect 2053 11169 2087 11203
rect 2087 11169 2096 11203
rect 2044 11160 2096 11169
rect 4344 11203 4396 11212
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 2136 11135 2188 11144
rect 2136 11101 2145 11135
rect 2145 11101 2179 11135
rect 2179 11101 2188 11135
rect 2136 11092 2188 11101
rect 4436 11092 4488 11144
rect 3056 11024 3108 11076
rect 4436 10999 4488 11008
rect 4436 10965 4445 10999
rect 4445 10965 4479 10999
rect 4479 10965 4488 10999
rect 5540 11160 5592 11212
rect 5724 11203 5776 11212
rect 5724 11169 5733 11203
rect 5733 11169 5767 11203
rect 5767 11169 5776 11203
rect 5724 11160 5776 11169
rect 7196 11296 7248 11348
rect 10232 11296 10284 11348
rect 11060 11339 11112 11348
rect 11060 11305 11069 11339
rect 11069 11305 11103 11339
rect 11103 11305 11112 11339
rect 11060 11296 11112 11305
rect 12716 11296 12768 11348
rect 13360 11296 13412 11348
rect 13544 11296 13596 11348
rect 9680 11228 9732 11280
rect 11336 11271 11388 11280
rect 11336 11237 11345 11271
rect 11345 11237 11379 11271
rect 11379 11237 11388 11271
rect 11336 11228 11388 11237
rect 11520 11228 11572 11280
rect 12992 11228 13044 11280
rect 13728 11271 13780 11280
rect 13728 11237 13737 11271
rect 13737 11237 13771 11271
rect 13771 11237 13780 11271
rect 13728 11228 13780 11237
rect 5448 11024 5500 11076
rect 7472 11067 7524 11076
rect 7472 11033 7481 11067
rect 7481 11033 7515 11067
rect 7515 11033 7524 11067
rect 7472 11024 7524 11033
rect 4436 10956 4488 10965
rect 5908 10956 5960 11008
rect 6736 10956 6788 11008
rect 8300 11160 8352 11212
rect 7748 11135 7800 11144
rect 7748 11101 7757 11135
rect 7757 11101 7791 11135
rect 7791 11101 7800 11135
rect 7748 11092 7800 11101
rect 8116 11092 8168 11144
rect 9404 11092 9456 11144
rect 12440 11160 12492 11212
rect 14832 11271 14884 11280
rect 14832 11237 14841 11271
rect 14841 11237 14875 11271
rect 14875 11237 14884 11271
rect 14832 11228 14884 11237
rect 15384 11228 15436 11280
rect 16488 11228 16540 11280
rect 12256 11092 12308 11144
rect 14004 11135 14056 11144
rect 14004 11101 14013 11135
rect 14013 11101 14047 11135
rect 14047 11101 14056 11135
rect 14004 11092 14056 11101
rect 14372 11024 14424 11076
rect 3680 10854 3732 10906
rect 3744 10854 3796 10906
rect 3808 10854 3860 10906
rect 3872 10854 3924 10906
rect 9078 10854 9130 10906
rect 9142 10854 9194 10906
rect 9206 10854 9258 10906
rect 9270 10854 9322 10906
rect 14475 10854 14527 10906
rect 14539 10854 14591 10906
rect 14603 10854 14655 10906
rect 14667 10854 14719 10906
rect 2136 10795 2188 10804
rect 2136 10761 2145 10795
rect 2145 10761 2179 10795
rect 2179 10761 2188 10795
rect 2136 10752 2188 10761
rect 3056 10795 3108 10804
rect 3056 10761 3065 10795
rect 3065 10761 3099 10795
rect 3099 10761 3108 10795
rect 3056 10752 3108 10761
rect 5724 10752 5776 10804
rect 11244 10752 11296 10804
rect 12992 10752 13044 10804
rect 16488 10752 16540 10804
rect 2228 10616 2280 10668
rect 3332 10616 3384 10668
rect 4436 10659 4488 10668
rect 2688 10591 2740 10600
rect 2688 10557 2697 10591
rect 2697 10557 2731 10591
rect 2731 10557 2740 10591
rect 2688 10548 2740 10557
rect 1676 10480 1728 10532
rect 2872 10523 2924 10532
rect 2872 10489 2881 10523
rect 2881 10489 2915 10523
rect 2915 10489 2924 10523
rect 2872 10480 2924 10489
rect 4436 10625 4445 10659
rect 4445 10625 4479 10659
rect 4479 10625 4488 10659
rect 4436 10616 4488 10625
rect 8576 10616 8628 10668
rect 9956 10616 10008 10668
rect 14096 10659 14148 10668
rect 14096 10625 14105 10659
rect 14105 10625 14139 10659
rect 14139 10625 14148 10659
rect 14096 10616 14148 10625
rect 16028 10616 16080 10668
rect 4712 10480 4764 10532
rect 5172 10480 5224 10532
rect 10232 10591 10284 10600
rect 10232 10557 10241 10591
rect 10241 10557 10275 10591
rect 10275 10557 10284 10591
rect 10232 10548 10284 10557
rect 11612 10548 11664 10600
rect 16212 10591 16264 10600
rect 16212 10557 16221 10591
rect 16221 10557 16255 10591
rect 16255 10557 16264 10591
rect 16212 10548 16264 10557
rect 14004 10480 14056 10532
rect 14832 10480 14884 10532
rect 1768 10455 1820 10464
rect 1768 10421 1777 10455
rect 1777 10421 1811 10455
rect 1811 10421 1820 10455
rect 1768 10412 1820 10421
rect 2596 10412 2648 10464
rect 3608 10412 3660 10464
rect 5908 10455 5960 10464
rect 5908 10421 5917 10455
rect 5917 10421 5951 10455
rect 5951 10421 5960 10455
rect 5908 10412 5960 10421
rect 7012 10412 7064 10464
rect 7380 10412 7432 10464
rect 8208 10455 8260 10464
rect 8208 10421 8217 10455
rect 8217 10421 8251 10455
rect 8251 10421 8260 10455
rect 8208 10412 8260 10421
rect 9128 10412 9180 10464
rect 9404 10412 9456 10464
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 6571 10310 6623 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 11904 10310 11956 10362
rect 11968 10310 12020 10362
rect 1492 10251 1544 10260
rect 1492 10217 1501 10251
rect 1501 10217 1535 10251
rect 1535 10217 1544 10251
rect 1492 10208 1544 10217
rect 3608 10251 3660 10260
rect 3608 10217 3617 10251
rect 3617 10217 3651 10251
rect 3651 10217 3660 10251
rect 3608 10208 3660 10217
rect 5172 10208 5224 10260
rect 6276 10208 6328 10260
rect 6828 10208 6880 10260
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 9588 10208 9640 10260
rect 14832 10208 14884 10260
rect 2044 10072 2096 10124
rect 2780 10072 2832 10124
rect 1768 10004 1820 10056
rect 3056 9936 3108 9988
rect 2596 9911 2648 9920
rect 2596 9877 2605 9911
rect 2605 9877 2639 9911
rect 2639 9877 2648 9911
rect 2596 9868 2648 9877
rect 8208 10140 8260 10192
rect 5356 10072 5408 10124
rect 5816 10072 5868 10124
rect 6276 10047 6328 10056
rect 6276 10013 6285 10047
rect 6285 10013 6319 10047
rect 6319 10013 6328 10047
rect 6276 10004 6328 10013
rect 7012 10072 7064 10124
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 9588 10072 9640 10124
rect 16212 10072 16264 10124
rect 8300 9936 8352 9988
rect 9404 9936 9456 9988
rect 8852 9868 8904 9920
rect 9680 9911 9732 9920
rect 9680 9877 9689 9911
rect 9689 9877 9723 9911
rect 9723 9877 9732 9911
rect 9680 9868 9732 9877
rect 3680 9766 3732 9818
rect 3744 9766 3796 9818
rect 3808 9766 3860 9818
rect 3872 9766 3924 9818
rect 9078 9766 9130 9818
rect 9142 9766 9194 9818
rect 9206 9766 9258 9818
rect 9270 9766 9322 9818
rect 14475 9766 14527 9818
rect 14539 9766 14591 9818
rect 14603 9766 14655 9818
rect 14667 9766 14719 9818
rect 2780 9707 2832 9716
rect 2780 9673 2789 9707
rect 2789 9673 2823 9707
rect 2823 9673 2832 9707
rect 2780 9664 2832 9673
rect 5908 9664 5960 9716
rect 6736 9664 6788 9716
rect 6828 9664 6880 9716
rect 9404 9664 9456 9716
rect 10508 9664 10560 9716
rect 1676 9596 1728 9648
rect 1860 9571 1912 9580
rect 1860 9537 1869 9571
rect 1869 9537 1903 9571
rect 1903 9537 1912 9571
rect 1860 9528 1912 9537
rect 6000 9596 6052 9648
rect 6184 9596 6236 9648
rect 6552 9596 6604 9648
rect 6920 9596 6972 9648
rect 7840 9596 7892 9648
rect 10692 9596 10744 9648
rect 4620 9528 4672 9580
rect 7196 9571 7248 9580
rect 7196 9537 7205 9571
rect 7205 9537 7239 9571
rect 7239 9537 7248 9571
rect 7196 9528 7248 9537
rect 3976 9503 4028 9512
rect 3976 9469 3985 9503
rect 3985 9469 4019 9503
rect 4019 9469 4028 9503
rect 3976 9460 4028 9469
rect 4252 9460 4304 9512
rect 5264 9503 5316 9512
rect 5264 9469 5273 9503
rect 5273 9469 5307 9503
rect 5307 9469 5316 9503
rect 5264 9460 5316 9469
rect 6000 9503 6052 9512
rect 6000 9469 6009 9503
rect 6009 9469 6043 9503
rect 6043 9469 6052 9503
rect 6000 9460 6052 9469
rect 6276 9460 6328 9512
rect 7288 9503 7340 9512
rect 2320 9392 2372 9444
rect 5632 9392 5684 9444
rect 6736 9392 6788 9444
rect 7288 9469 7297 9503
rect 7297 9469 7331 9503
rect 7331 9469 7340 9503
rect 7288 9460 7340 9469
rect 7564 9503 7616 9512
rect 7564 9469 7573 9503
rect 7573 9469 7607 9503
rect 7607 9469 7616 9503
rect 7564 9460 7616 9469
rect 9036 9528 9088 9580
rect 9496 9528 9548 9580
rect 12440 9528 12492 9580
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 13176 9528 13228 9580
rect 7932 9460 7984 9512
rect 8024 9503 8076 9512
rect 8024 9469 8033 9503
rect 8033 9469 8067 9503
rect 8067 9469 8076 9503
rect 8024 9460 8076 9469
rect 9220 9503 9272 9512
rect 9220 9469 9229 9503
rect 9229 9469 9263 9503
rect 9263 9469 9272 9503
rect 9404 9503 9456 9512
rect 9220 9460 9272 9469
rect 9404 9469 9413 9503
rect 9413 9469 9447 9503
rect 9447 9469 9456 9503
rect 9404 9460 9456 9469
rect 10692 9503 10744 9512
rect 10692 9469 10701 9503
rect 10701 9469 10735 9503
rect 10735 9469 10744 9503
rect 10692 9460 10744 9469
rect 11244 9503 11296 9512
rect 11244 9469 11253 9503
rect 11253 9469 11287 9503
rect 11287 9469 11296 9503
rect 11244 9460 11296 9469
rect 16672 9528 16724 9580
rect 16764 9503 16816 9512
rect 16764 9469 16773 9503
rect 16773 9469 16807 9503
rect 16807 9469 16816 9503
rect 16764 9460 16816 9469
rect 9496 9392 9548 9444
rect 1400 9367 1452 9376
rect 1400 9333 1409 9367
rect 1409 9333 1443 9367
rect 1443 9333 1452 9367
rect 1400 9324 1452 9333
rect 4160 9324 4212 9376
rect 5172 9324 5224 9376
rect 5356 9367 5408 9376
rect 5356 9333 5365 9367
rect 5365 9333 5399 9367
rect 5399 9333 5408 9367
rect 5356 9324 5408 9333
rect 6920 9324 6972 9376
rect 7196 9324 7248 9376
rect 8392 9324 8444 9376
rect 9404 9324 9456 9376
rect 11244 9324 11296 9376
rect 11612 9324 11664 9376
rect 12164 9367 12216 9376
rect 12164 9333 12173 9367
rect 12173 9333 12207 9367
rect 12207 9333 12216 9367
rect 12164 9324 12216 9333
rect 12992 9367 13044 9376
rect 12992 9333 13001 9367
rect 13001 9333 13035 9367
rect 13035 9333 13044 9367
rect 13360 9367 13412 9376
rect 12992 9324 13044 9333
rect 13360 9333 13369 9367
rect 13369 9333 13403 9367
rect 13403 9333 13412 9367
rect 13360 9324 13412 9333
rect 15476 9324 15528 9376
rect 16580 9367 16632 9376
rect 16580 9333 16589 9367
rect 16589 9333 16623 9367
rect 16623 9333 16632 9367
rect 16580 9324 16632 9333
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 6571 9222 6623 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 11904 9222 11956 9274
rect 11968 9222 12020 9274
rect 5080 9163 5132 9172
rect 5080 9129 5089 9163
rect 5089 9129 5123 9163
rect 5123 9129 5132 9163
rect 5080 9120 5132 9129
rect 8024 9120 8076 9172
rect 8116 9120 8168 9172
rect 8208 9120 8260 9172
rect 5172 9052 5224 9104
rect 6920 9052 6972 9104
rect 8944 9052 8996 9104
rect 9220 9052 9272 9104
rect 9956 9120 10008 9172
rect 11612 9163 11664 9172
rect 2964 9027 3016 9036
rect 2964 8993 2973 9027
rect 2973 8993 3007 9027
rect 3007 8993 3016 9027
rect 2964 8984 3016 8993
rect 5724 8984 5776 9036
rect 6092 8984 6144 9036
rect 6828 8984 6880 9036
rect 7656 8984 7708 9036
rect 8300 8984 8352 9036
rect 9036 8984 9088 9036
rect 9312 8984 9364 9036
rect 9588 9027 9640 9036
rect 9588 8993 9597 9027
rect 9597 8993 9631 9027
rect 9631 8993 9640 9027
rect 9588 8984 9640 8993
rect 9772 8984 9824 9036
rect 10600 9027 10652 9036
rect 10600 8993 10609 9027
rect 10609 8993 10643 9027
rect 10643 8993 10652 9027
rect 10600 8984 10652 8993
rect 5080 8959 5132 8968
rect 5080 8925 5089 8959
rect 5089 8925 5123 8959
rect 5123 8925 5132 8959
rect 5080 8916 5132 8925
rect 5172 8959 5224 8968
rect 5172 8925 5181 8959
rect 5181 8925 5215 8959
rect 5215 8925 5224 8959
rect 5172 8916 5224 8925
rect 7380 8916 7432 8968
rect 7564 8916 7616 8968
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 9496 8959 9548 8968
rect 9496 8925 9505 8959
rect 9505 8925 9539 8959
rect 9539 8925 9548 8959
rect 11612 9129 11621 9163
rect 11621 9129 11655 9163
rect 11655 9129 11664 9163
rect 11612 9120 11664 9129
rect 12164 9052 12216 9104
rect 12992 9120 13044 9172
rect 12440 9027 12492 9036
rect 9496 8916 9548 8925
rect 10968 8916 11020 8968
rect 11428 8916 11480 8968
rect 12440 8993 12449 9027
rect 12449 8993 12483 9027
rect 12483 8993 12492 9027
rect 12440 8984 12492 8993
rect 12624 8984 12676 9036
rect 13268 8984 13320 9036
rect 14004 8984 14056 9036
rect 12808 8916 12860 8968
rect 13084 8916 13136 8968
rect 16120 9120 16172 9172
rect 14924 8984 14976 9036
rect 15476 9027 15528 9036
rect 15476 8993 15485 9027
rect 15485 8993 15519 9027
rect 15519 8993 15528 9027
rect 15476 8984 15528 8993
rect 15844 8984 15896 9036
rect 3240 8848 3292 8900
rect 2228 8780 2280 8832
rect 3976 8780 4028 8832
rect 5816 8780 5868 8832
rect 9680 8780 9732 8832
rect 11336 8780 11388 8832
rect 13912 8848 13964 8900
rect 14372 8780 14424 8832
rect 3680 8678 3732 8730
rect 3744 8678 3796 8730
rect 3808 8678 3860 8730
rect 3872 8678 3924 8730
rect 9078 8678 9130 8730
rect 9142 8678 9194 8730
rect 9206 8678 9258 8730
rect 9270 8678 9322 8730
rect 14475 8678 14527 8730
rect 14539 8678 14591 8730
rect 14603 8678 14655 8730
rect 14667 8678 14719 8730
rect 1676 8576 1728 8628
rect 2228 8551 2280 8560
rect 2228 8517 2237 8551
rect 2237 8517 2271 8551
rect 2271 8517 2280 8551
rect 2228 8508 2280 8517
rect 5080 8576 5132 8628
rect 1400 8440 1452 8492
rect 2504 8372 2556 8424
rect 4528 8440 4580 8492
rect 5172 8508 5224 8560
rect 1400 8347 1452 8356
rect 1400 8313 1409 8347
rect 1409 8313 1443 8347
rect 1443 8313 1452 8347
rect 1400 8304 1452 8313
rect 2044 8304 2096 8356
rect 2964 8304 3016 8356
rect 5724 8508 5776 8560
rect 6092 8551 6144 8560
rect 6092 8517 6101 8551
rect 6101 8517 6135 8551
rect 6135 8517 6144 8551
rect 6092 8508 6144 8517
rect 5632 8483 5684 8492
rect 5632 8449 5641 8483
rect 5641 8449 5675 8483
rect 5675 8449 5684 8483
rect 5632 8440 5684 8449
rect 5724 8415 5776 8424
rect 5724 8381 5733 8415
rect 5733 8381 5767 8415
rect 5767 8381 5776 8415
rect 6000 8415 6052 8424
rect 5724 8372 5776 8381
rect 6000 8381 6009 8415
rect 6009 8381 6043 8415
rect 6043 8381 6052 8415
rect 6000 8372 6052 8381
rect 7380 8440 7432 8492
rect 8208 8508 8260 8560
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 7932 8483 7984 8492
rect 7932 8449 7941 8483
rect 7941 8449 7975 8483
rect 7975 8449 7984 8483
rect 7932 8440 7984 8449
rect 6736 8372 6788 8424
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 7656 8415 7708 8424
rect 7656 8381 7665 8415
rect 7665 8381 7699 8415
rect 7699 8381 7708 8415
rect 7656 8372 7708 8381
rect 7840 8372 7892 8424
rect 9404 8508 9456 8560
rect 8852 8440 8904 8492
rect 9680 8508 9732 8560
rect 10968 8508 11020 8560
rect 11244 8483 11296 8492
rect 11244 8449 11253 8483
rect 11253 8449 11287 8483
rect 11287 8449 11296 8483
rect 11244 8440 11296 8449
rect 9496 8415 9548 8424
rect 9496 8381 9505 8415
rect 9505 8381 9539 8415
rect 9539 8381 9548 8415
rect 9496 8372 9548 8381
rect 9680 8415 9732 8424
rect 9680 8381 9682 8415
rect 9682 8381 9716 8415
rect 9716 8381 9732 8415
rect 9680 8372 9732 8381
rect 10232 8372 10284 8424
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 15568 8508 15620 8560
rect 2320 8236 2372 8288
rect 5816 8304 5868 8356
rect 4160 8279 4212 8288
rect 4160 8245 4169 8279
rect 4169 8245 4203 8279
rect 4203 8245 4212 8279
rect 4160 8236 4212 8245
rect 4620 8236 4672 8288
rect 6184 8236 6236 8288
rect 10508 8304 10560 8356
rect 13268 8372 13320 8424
rect 16580 8440 16632 8492
rect 13912 8415 13964 8424
rect 13912 8381 13921 8415
rect 13921 8381 13955 8415
rect 13955 8381 13964 8415
rect 13912 8372 13964 8381
rect 16120 8415 16172 8424
rect 16120 8381 16129 8415
rect 16129 8381 16163 8415
rect 16163 8381 16172 8415
rect 16120 8372 16172 8381
rect 14096 8347 14148 8356
rect 14096 8313 14105 8347
rect 14105 8313 14139 8347
rect 14139 8313 14148 8347
rect 14096 8304 14148 8313
rect 15936 8347 15988 8356
rect 15936 8313 15945 8347
rect 15945 8313 15979 8347
rect 15979 8313 15988 8347
rect 15936 8304 15988 8313
rect 8760 8236 8812 8288
rect 9680 8236 9732 8288
rect 10692 8236 10744 8288
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 6571 8134 6623 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 11904 8134 11956 8186
rect 11968 8134 12020 8186
rect 6092 8032 6144 8084
rect 12532 8032 12584 8084
rect 2320 7964 2372 8016
rect 5632 7964 5684 8016
rect 1492 7896 1544 7948
rect 2504 7896 2556 7948
rect 5540 7896 5592 7948
rect 6736 7964 6788 8016
rect 5172 7828 5224 7880
rect 7380 7939 7432 7948
rect 7380 7905 7389 7939
rect 7389 7905 7423 7939
rect 7423 7905 7432 7939
rect 7932 7939 7984 7948
rect 7380 7896 7432 7905
rect 5908 7828 5960 7880
rect 6828 7871 6880 7880
rect 6828 7837 6837 7871
rect 6837 7837 6871 7871
rect 6871 7837 6880 7871
rect 7932 7905 7941 7939
rect 7941 7905 7975 7939
rect 7975 7905 7984 7939
rect 7932 7896 7984 7905
rect 9956 7939 10008 7948
rect 9956 7905 9965 7939
rect 9965 7905 9999 7939
rect 9999 7905 10008 7939
rect 9956 7896 10008 7905
rect 6828 7828 6880 7837
rect 8116 7828 8168 7880
rect 6184 7760 6236 7812
rect 15844 7939 15896 7948
rect 15844 7905 15853 7939
rect 15853 7905 15887 7939
rect 15887 7905 15896 7939
rect 15844 7896 15896 7905
rect 15936 7939 15988 7948
rect 15936 7905 15945 7939
rect 15945 7905 15979 7939
rect 15979 7905 15988 7939
rect 15936 7896 15988 7905
rect 14924 7803 14976 7812
rect 14924 7769 14933 7803
rect 14933 7769 14967 7803
rect 14967 7769 14976 7803
rect 14924 7760 14976 7769
rect 6920 7692 6972 7744
rect 8300 7692 8352 7744
rect 3680 7590 3732 7642
rect 3744 7590 3796 7642
rect 3808 7590 3860 7642
rect 3872 7590 3924 7642
rect 9078 7590 9130 7642
rect 9142 7590 9194 7642
rect 9206 7590 9258 7642
rect 9270 7590 9322 7642
rect 14475 7590 14527 7642
rect 14539 7590 14591 7642
rect 14603 7590 14655 7642
rect 14667 7590 14719 7642
rect 2504 7531 2556 7540
rect 2504 7497 2513 7531
rect 2513 7497 2547 7531
rect 2547 7497 2556 7531
rect 2504 7488 2556 7497
rect 8852 7488 8904 7540
rect 1952 7420 2004 7472
rect 4160 7352 4212 7404
rect 5080 7284 5132 7336
rect 2504 7216 2556 7268
rect 4988 7216 5040 7268
rect 6092 7420 6144 7472
rect 7840 7420 7892 7472
rect 10600 7488 10652 7540
rect 11336 7420 11388 7472
rect 14096 7420 14148 7472
rect 6920 7395 6972 7404
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 6920 7352 6972 7361
rect 7656 7352 7708 7404
rect 8208 7352 8260 7404
rect 8300 7352 8352 7404
rect 10600 7352 10652 7404
rect 6184 7284 6236 7336
rect 7380 7284 7432 7336
rect 8024 7327 8076 7336
rect 8024 7293 8033 7327
rect 8033 7293 8067 7327
rect 8067 7293 8076 7327
rect 8024 7284 8076 7293
rect 8392 7327 8444 7336
rect 8392 7293 8401 7327
rect 8401 7293 8435 7327
rect 8435 7293 8444 7327
rect 8392 7284 8444 7293
rect 4436 7191 4488 7200
rect 4436 7157 4445 7191
rect 4445 7157 4479 7191
rect 4479 7157 4488 7191
rect 4436 7148 4488 7157
rect 4896 7148 4948 7200
rect 8760 7259 8812 7268
rect 8760 7225 8769 7259
rect 8769 7225 8803 7259
rect 8803 7225 8812 7259
rect 8760 7216 8812 7225
rect 8944 7259 8996 7268
rect 8944 7225 8974 7259
rect 8974 7225 8996 7259
rect 8944 7216 8996 7225
rect 8300 7148 8352 7200
rect 8852 7148 8904 7200
rect 9588 7148 9640 7200
rect 9864 7259 9916 7268
rect 9864 7225 9873 7259
rect 9873 7225 9907 7259
rect 9907 7225 9916 7259
rect 11060 7284 11112 7336
rect 12072 7284 12124 7336
rect 12624 7327 12676 7336
rect 12624 7293 12633 7327
rect 12633 7293 12667 7327
rect 12667 7293 12676 7327
rect 12624 7284 12676 7293
rect 13268 7352 13320 7404
rect 14004 7284 14056 7336
rect 14924 7284 14976 7336
rect 10968 7259 11020 7268
rect 9864 7216 9916 7225
rect 10968 7225 10977 7259
rect 10977 7225 11011 7259
rect 11011 7225 11020 7259
rect 10968 7216 11020 7225
rect 9956 7148 10008 7200
rect 12808 7191 12860 7200
rect 12808 7157 12817 7191
rect 12817 7157 12851 7191
rect 12851 7157 12860 7191
rect 12808 7148 12860 7157
rect 13544 7148 13596 7200
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 6571 7046 6623 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 11904 7046 11956 7098
rect 11968 7046 12020 7098
rect 8300 6987 8352 6996
rect 8300 6953 8309 6987
rect 8309 6953 8343 6987
rect 8343 6953 8352 6987
rect 8300 6944 8352 6953
rect 4436 6919 4488 6928
rect 4436 6885 4445 6919
rect 4445 6885 4479 6919
rect 4479 6885 4488 6919
rect 4436 6876 4488 6885
rect 4988 6919 5040 6928
rect 4988 6885 4997 6919
rect 4997 6885 5031 6919
rect 5031 6885 5040 6919
rect 4988 6876 5040 6885
rect 8484 6876 8536 6928
rect 1584 6808 1636 6860
rect 3976 6808 4028 6860
rect 4160 6808 4212 6860
rect 4896 6808 4948 6860
rect 6276 6808 6328 6860
rect 7472 6851 7524 6860
rect 7472 6817 7481 6851
rect 7481 6817 7515 6851
rect 7515 6817 7524 6851
rect 7472 6808 7524 6817
rect 7656 6851 7708 6860
rect 7656 6817 7665 6851
rect 7665 6817 7699 6851
rect 7699 6817 7708 6851
rect 7656 6808 7708 6817
rect 7840 6808 7892 6860
rect 8944 6808 8996 6860
rect 10784 6944 10836 6996
rect 12808 6944 12860 6996
rect 15844 6944 15896 6996
rect 10968 6876 11020 6928
rect 12532 6919 12584 6928
rect 11152 6851 11204 6860
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 5724 6740 5776 6792
rect 8024 6783 8076 6792
rect 2504 6672 2556 6724
rect 5080 6672 5132 6724
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 8392 6740 8444 6792
rect 6828 6672 6880 6724
rect 9496 6740 9548 6792
rect 11152 6817 11161 6851
rect 11161 6817 11195 6851
rect 11195 6817 11204 6851
rect 11152 6808 11204 6817
rect 12532 6885 12541 6919
rect 12541 6885 12575 6919
rect 12575 6885 12584 6919
rect 12532 6876 12584 6885
rect 12072 6851 12124 6860
rect 12072 6817 12081 6851
rect 12081 6817 12115 6851
rect 12115 6817 12124 6851
rect 12072 6808 12124 6817
rect 10876 6715 10928 6724
rect 10876 6681 10885 6715
rect 10885 6681 10919 6715
rect 10919 6681 10928 6715
rect 10876 6672 10928 6681
rect 2412 6604 2464 6656
rect 6000 6604 6052 6656
rect 7288 6647 7340 6656
rect 7288 6613 7297 6647
rect 7297 6613 7331 6647
rect 7331 6613 7340 6647
rect 7288 6604 7340 6613
rect 7380 6604 7432 6656
rect 8024 6604 8076 6656
rect 9588 6647 9640 6656
rect 9588 6613 9597 6647
rect 9597 6613 9631 6647
rect 9631 6613 9640 6647
rect 9588 6604 9640 6613
rect 12532 6740 12584 6792
rect 13084 6740 13136 6792
rect 15844 6808 15896 6860
rect 16948 6851 17000 6860
rect 16948 6817 16957 6851
rect 16957 6817 16991 6851
rect 16991 6817 17000 6851
rect 16948 6808 17000 6817
rect 13268 6715 13320 6724
rect 13268 6681 13277 6715
rect 13277 6681 13311 6715
rect 13311 6681 13320 6715
rect 13268 6672 13320 6681
rect 16580 6604 16632 6656
rect 3680 6502 3732 6554
rect 3744 6502 3796 6554
rect 3808 6502 3860 6554
rect 3872 6502 3924 6554
rect 9078 6502 9130 6554
rect 9142 6502 9194 6554
rect 9206 6502 9258 6554
rect 9270 6502 9322 6554
rect 14475 6502 14527 6554
rect 14539 6502 14591 6554
rect 14603 6502 14655 6554
rect 14667 6502 14719 6554
rect 7656 6400 7708 6452
rect 10876 6443 10928 6452
rect 10876 6409 10885 6443
rect 10885 6409 10919 6443
rect 10919 6409 10928 6443
rect 10876 6400 10928 6409
rect 11060 6443 11112 6452
rect 11060 6409 11069 6443
rect 11069 6409 11103 6443
rect 11103 6409 11112 6443
rect 11060 6400 11112 6409
rect 15844 6443 15896 6452
rect 15844 6409 15853 6443
rect 15853 6409 15887 6443
rect 15887 6409 15896 6443
rect 15844 6400 15896 6409
rect 6000 6332 6052 6384
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 2504 6128 2556 6180
rect 3976 6196 4028 6248
rect 5816 6196 5868 6248
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 7840 6264 7892 6316
rect 11336 6264 11388 6316
rect 7288 6196 7340 6248
rect 7472 6196 7524 6248
rect 8760 6196 8812 6248
rect 4896 6128 4948 6180
rect 5908 6171 5960 6180
rect 5908 6137 5917 6171
rect 5917 6137 5951 6171
rect 5951 6137 5960 6171
rect 5908 6128 5960 6137
rect 10784 6196 10836 6248
rect 13544 6239 13596 6248
rect 13544 6205 13553 6239
rect 13553 6205 13587 6239
rect 13587 6205 13596 6239
rect 13544 6196 13596 6205
rect 15292 6196 15344 6248
rect 15844 6239 15896 6248
rect 15844 6205 15853 6239
rect 15853 6205 15887 6239
rect 15887 6205 15896 6239
rect 15844 6196 15896 6205
rect 11152 6128 11204 6180
rect 1584 6060 1636 6112
rect 2320 6103 2372 6112
rect 2320 6069 2329 6103
rect 2329 6069 2363 6103
rect 2363 6069 2372 6103
rect 2320 6060 2372 6069
rect 6828 6103 6880 6112
rect 6828 6069 6837 6103
rect 6837 6069 6871 6103
rect 6871 6069 6880 6103
rect 6828 6060 6880 6069
rect 7104 6060 7156 6112
rect 8300 6103 8352 6112
rect 8300 6069 8309 6103
rect 8309 6069 8343 6103
rect 8343 6069 8352 6103
rect 8300 6060 8352 6069
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 6571 5958 6623 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 11904 5958 11956 6010
rect 11968 5958 12020 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 4252 5831 4304 5840
rect 4252 5797 4261 5831
rect 4261 5797 4295 5831
rect 4295 5797 4304 5831
rect 4252 5788 4304 5797
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 4804 5856 4856 5908
rect 12072 5899 12124 5908
rect 12072 5865 12081 5899
rect 12081 5865 12115 5899
rect 12115 5865 12124 5899
rect 12072 5856 12124 5865
rect 15844 5899 15896 5908
rect 15844 5865 15853 5899
rect 15853 5865 15887 5899
rect 15887 5865 15896 5899
rect 15844 5856 15896 5865
rect 4804 5763 4856 5772
rect 4804 5729 4813 5763
rect 4813 5729 4847 5763
rect 4847 5729 4856 5763
rect 4804 5720 4856 5729
rect 10232 5763 10284 5772
rect 10232 5729 10241 5763
rect 10241 5729 10275 5763
rect 10275 5729 10284 5763
rect 10232 5720 10284 5729
rect 12440 5763 12492 5772
rect 12440 5729 12449 5763
rect 12449 5729 12483 5763
rect 12483 5729 12492 5763
rect 12440 5720 12492 5729
rect 15844 5720 15896 5772
rect 11704 5695 11756 5704
rect 11704 5661 11713 5695
rect 11713 5661 11747 5695
rect 11747 5661 11756 5695
rect 11704 5652 11756 5661
rect 10140 5559 10192 5568
rect 10140 5525 10149 5559
rect 10149 5525 10183 5559
rect 10183 5525 10192 5559
rect 10140 5516 10192 5525
rect 3680 5414 3732 5466
rect 3744 5414 3796 5466
rect 3808 5414 3860 5466
rect 3872 5414 3924 5466
rect 9078 5414 9130 5466
rect 9142 5414 9194 5466
rect 9206 5414 9258 5466
rect 9270 5414 9322 5466
rect 14475 5414 14527 5466
rect 14539 5414 14591 5466
rect 14603 5414 14655 5466
rect 14667 5414 14719 5466
rect 12440 5312 12492 5364
rect 2412 5244 2464 5296
rect 2412 5151 2464 5160
rect 2412 5117 2421 5151
rect 2421 5117 2455 5151
rect 2455 5117 2464 5151
rect 4252 5176 4304 5228
rect 7380 5176 7432 5228
rect 8116 5176 8168 5228
rect 2412 5108 2464 5117
rect 2872 5108 2924 5160
rect 5816 5108 5868 5160
rect 8300 5108 8352 5160
rect 9404 5151 9456 5160
rect 9404 5117 9413 5151
rect 9413 5117 9447 5151
rect 9447 5117 9456 5151
rect 9404 5108 9456 5117
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 12072 5219 12124 5228
rect 5080 5083 5132 5092
rect 5080 5049 5089 5083
rect 5089 5049 5123 5083
rect 5123 5049 5132 5083
rect 5080 5040 5132 5049
rect 7104 5040 7156 5092
rect 8760 5040 8812 5092
rect 10600 5151 10652 5160
rect 10600 5117 10609 5151
rect 10609 5117 10643 5151
rect 10643 5117 10652 5151
rect 10600 5108 10652 5117
rect 10692 5151 10744 5160
rect 10692 5117 10701 5151
rect 10701 5117 10735 5151
rect 10735 5117 10744 5151
rect 12072 5185 12081 5219
rect 12081 5185 12115 5219
rect 12115 5185 12124 5219
rect 12072 5176 12124 5185
rect 10692 5108 10744 5117
rect 11704 5151 11756 5160
rect 11704 5117 11713 5151
rect 11713 5117 11747 5151
rect 11747 5117 11756 5151
rect 11704 5108 11756 5117
rect 13360 5219 13412 5228
rect 13360 5185 13369 5219
rect 13369 5185 13403 5219
rect 13403 5185 13412 5219
rect 13360 5176 13412 5185
rect 15292 5176 15344 5228
rect 15384 5151 15436 5160
rect 15384 5117 15393 5151
rect 15393 5117 15427 5151
rect 15427 5117 15436 5151
rect 15384 5108 15436 5117
rect 2872 4972 2924 5024
rect 6000 4972 6052 5024
rect 8024 4972 8076 5024
rect 8576 5015 8628 5024
rect 8576 4981 8585 5015
rect 8585 4981 8619 5015
rect 8619 4981 8628 5015
rect 8576 4972 8628 4981
rect 8668 4972 8720 5024
rect 12440 5083 12492 5092
rect 12440 5049 12449 5083
rect 12449 5049 12483 5083
rect 12483 5049 12492 5083
rect 12440 5040 12492 5049
rect 10232 4972 10284 5024
rect 12072 4972 12124 5024
rect 15844 5015 15896 5024
rect 15844 4981 15853 5015
rect 15853 4981 15887 5015
rect 15887 4981 15896 5015
rect 15844 4972 15896 4981
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 6571 4870 6623 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 11904 4870 11956 4922
rect 11968 4870 12020 4922
rect 2780 4811 2832 4820
rect 2780 4777 2789 4811
rect 2789 4777 2823 4811
rect 2823 4777 2832 4811
rect 2780 4768 2832 4777
rect 2872 4743 2924 4752
rect 2872 4709 2881 4743
rect 2881 4709 2915 4743
rect 2915 4709 2924 4743
rect 2872 4700 2924 4709
rect 4252 4700 4304 4752
rect 2964 4632 3016 4684
rect 5080 4768 5132 4820
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 6000 4675 6052 4684
rect 6000 4641 6009 4675
rect 6009 4641 6043 4675
rect 6043 4641 6052 4675
rect 6000 4632 6052 4641
rect 6828 4564 6880 4616
rect 7288 4632 7340 4684
rect 7380 4607 7432 4616
rect 7380 4573 7389 4607
rect 7389 4573 7423 4607
rect 7423 4573 7432 4607
rect 7380 4564 7432 4573
rect 14372 4768 14424 4820
rect 15384 4768 15436 4820
rect 8024 4700 8076 4752
rect 8760 4675 8812 4684
rect 8760 4641 8769 4675
rect 8769 4641 8803 4675
rect 8803 4641 8812 4675
rect 8760 4632 8812 4641
rect 8576 4564 8628 4616
rect 10140 4632 10192 4684
rect 11060 4675 11112 4684
rect 11060 4641 11069 4675
rect 11069 4641 11103 4675
rect 11103 4641 11112 4675
rect 11060 4632 11112 4641
rect 16948 4675 17000 4684
rect 16948 4641 16957 4675
rect 16957 4641 16991 4675
rect 16991 4641 17000 4675
rect 16948 4632 17000 4641
rect 12532 4564 12584 4616
rect 15384 4564 15436 4616
rect 12440 4496 12492 4548
rect 4160 4471 4212 4480
rect 4160 4437 4169 4471
rect 4169 4437 4203 4471
rect 4203 4437 4212 4471
rect 4160 4428 4212 4437
rect 8576 4428 8628 4480
rect 3680 4326 3732 4378
rect 3744 4326 3796 4378
rect 3808 4326 3860 4378
rect 3872 4326 3924 4378
rect 9078 4326 9130 4378
rect 9142 4326 9194 4378
rect 9206 4326 9258 4378
rect 9270 4326 9322 4378
rect 14475 4326 14527 4378
rect 14539 4326 14591 4378
rect 14603 4326 14655 4378
rect 14667 4326 14719 4378
rect 7380 4224 7432 4276
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 2044 4088 2096 4140
rect 4160 4063 4212 4072
rect 4160 4029 4169 4063
rect 4169 4029 4203 4063
rect 4203 4029 4212 4063
rect 4160 4020 4212 4029
rect 6828 4088 6880 4140
rect 12716 4131 12768 4140
rect 12716 4097 12725 4131
rect 12725 4097 12759 4131
rect 12759 4097 12768 4131
rect 12716 4088 12768 4097
rect 13636 4088 13688 4140
rect 7012 4063 7064 4072
rect 7012 4029 7021 4063
rect 7021 4029 7055 4063
rect 7055 4029 7064 4063
rect 7288 4063 7340 4072
rect 7012 4020 7064 4029
rect 7288 4029 7297 4063
rect 7297 4029 7331 4063
rect 7331 4029 7340 4063
rect 7288 4020 7340 4029
rect 13820 4063 13872 4072
rect 1584 3995 1636 4004
rect 1584 3961 1593 3995
rect 1593 3961 1627 3995
rect 1627 3961 1636 3995
rect 1584 3952 1636 3961
rect 4712 3995 4764 4004
rect 4712 3961 4721 3995
rect 4721 3961 4755 3995
rect 4755 3961 4764 3995
rect 4712 3952 4764 3961
rect 13268 3952 13320 4004
rect 13820 4029 13829 4063
rect 13829 4029 13863 4063
rect 13863 4029 13872 4063
rect 13820 4020 13872 4029
rect 14188 4063 14240 4072
rect 14188 4029 14197 4063
rect 14197 4029 14231 4063
rect 14231 4029 14240 4063
rect 14188 4020 14240 4029
rect 14280 3952 14332 4004
rect 16856 3952 16908 4004
rect 7012 3884 7064 3936
rect 7196 3884 7248 3936
rect 11336 3884 11388 3936
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 13176 3927 13228 3936
rect 12440 3884 12492 3893
rect 13176 3893 13185 3927
rect 13185 3893 13219 3927
rect 13219 3893 13228 3927
rect 13176 3884 13228 3893
rect 14372 3927 14424 3936
rect 14372 3893 14381 3927
rect 14381 3893 14415 3927
rect 14415 3893 14424 3927
rect 14372 3884 14424 3893
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 6571 3782 6623 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 11904 3782 11956 3834
rect 11968 3782 12020 3834
rect 2780 3612 2832 3664
rect 5264 3612 5316 3664
rect 7288 3612 7340 3664
rect 8576 3655 8628 3664
rect 8576 3621 8585 3655
rect 8585 3621 8619 3655
rect 8619 3621 8628 3655
rect 8576 3612 8628 3621
rect 1584 3544 1636 3596
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 7472 3544 7524 3596
rect 10324 3680 10376 3732
rect 11060 3723 11112 3732
rect 11060 3689 11069 3723
rect 11069 3689 11103 3723
rect 11103 3689 11112 3723
rect 11060 3680 11112 3689
rect 13636 3680 13688 3732
rect 12716 3612 12768 3664
rect 10600 3544 10652 3596
rect 10968 3587 11020 3596
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 13268 3587 13320 3596
rect 13268 3553 13277 3587
rect 13277 3553 13311 3587
rect 13311 3553 13320 3587
rect 13268 3544 13320 3553
rect 13820 3612 13872 3664
rect 15476 3612 15528 3664
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 7196 3476 7248 3528
rect 7656 3476 7708 3528
rect 8024 3476 8076 3528
rect 9404 3519 9456 3528
rect 9404 3485 9413 3519
rect 9413 3485 9447 3519
rect 9447 3485 9456 3519
rect 9404 3476 9456 3485
rect 11060 3519 11112 3528
rect 11060 3485 11069 3519
rect 11069 3485 11103 3519
rect 11103 3485 11112 3519
rect 11060 3476 11112 3485
rect 12992 3476 13044 3528
rect 15016 3519 15068 3528
rect 7380 3383 7432 3392
rect 7380 3349 7389 3383
rect 7389 3349 7423 3383
rect 7423 3349 7432 3383
rect 7380 3340 7432 3349
rect 13728 3408 13780 3460
rect 15016 3485 15025 3519
rect 15025 3485 15059 3519
rect 15059 3485 15068 3519
rect 17040 3544 17092 3596
rect 15016 3476 15068 3485
rect 10140 3340 10192 3392
rect 15476 3340 15528 3392
rect 3680 3238 3732 3290
rect 3744 3238 3796 3290
rect 3808 3238 3860 3290
rect 3872 3238 3924 3290
rect 9078 3238 9130 3290
rect 9142 3238 9194 3290
rect 9206 3238 9258 3290
rect 9270 3238 9322 3290
rect 14475 3238 14527 3290
rect 14539 3238 14591 3290
rect 14603 3238 14655 3290
rect 14667 3238 14719 3290
rect 7380 3136 7432 3188
rect 7656 3136 7708 3188
rect 9404 3136 9456 3188
rect 1584 3000 1636 3052
rect 3148 3000 3200 3052
rect 480 2932 532 2984
rect 2412 2975 2464 2984
rect 2412 2941 2420 2975
rect 2420 2941 2464 2975
rect 2412 2932 2464 2941
rect 6000 3000 6052 3052
rect 6092 3000 6144 3052
rect 7288 3068 7340 3120
rect 8024 3068 8076 3120
rect 8116 3000 8168 3052
rect 8852 3000 8904 3052
rect 7288 2975 7340 2984
rect 7288 2941 7297 2975
rect 7297 2941 7331 2975
rect 7331 2941 7340 2975
rect 7288 2932 7340 2941
rect 7472 2975 7524 2984
rect 7472 2941 7481 2975
rect 7481 2941 7515 2975
rect 7515 2941 7524 2975
rect 7472 2932 7524 2941
rect 8024 2975 8076 2984
rect 8024 2941 8033 2975
rect 8033 2941 8067 2975
rect 8067 2941 8076 2975
rect 8024 2932 8076 2941
rect 9588 2975 9640 2984
rect 3056 2864 3108 2916
rect 9588 2941 9597 2975
rect 9597 2941 9631 2975
rect 9631 2941 9640 2975
rect 9588 2932 9640 2941
rect 1676 2796 1728 2848
rect 9680 2864 9732 2916
rect 10324 3136 10376 3188
rect 10968 3136 11020 3188
rect 12440 3179 12492 3188
rect 12440 3145 12449 3179
rect 12449 3145 12483 3179
rect 12483 3145 12492 3179
rect 12440 3136 12492 3145
rect 12532 3000 12584 3052
rect 10600 2975 10652 2984
rect 10600 2941 10609 2975
rect 10609 2941 10643 2975
rect 10643 2941 10652 2975
rect 10600 2932 10652 2941
rect 11336 2932 11388 2984
rect 10968 2864 11020 2916
rect 14188 3179 14240 3188
rect 14188 3145 14197 3179
rect 14197 3145 14231 3179
rect 14231 3145 14240 3179
rect 14188 3136 14240 3145
rect 15384 3179 15436 3188
rect 15384 3145 15393 3179
rect 15393 3145 15427 3179
rect 15427 3145 15436 3179
rect 15384 3136 15436 3145
rect 16580 3179 16632 3188
rect 16580 3145 16589 3179
rect 16589 3145 16623 3179
rect 16623 3145 16632 3179
rect 16580 3136 16632 3145
rect 13176 3000 13228 3052
rect 5264 2796 5316 2848
rect 10140 2796 10192 2848
rect 10508 2796 10560 2848
rect 13636 3000 13688 3052
rect 14372 3000 14424 3052
rect 13728 2975 13780 2984
rect 13728 2941 13737 2975
rect 13737 2941 13771 2975
rect 13771 2941 13780 2975
rect 13728 2932 13780 2941
rect 14280 2975 14332 2984
rect 14280 2941 14289 2975
rect 14289 2941 14323 2975
rect 14323 2941 14332 2975
rect 14280 2932 14332 2941
rect 15016 2975 15068 2984
rect 15016 2941 15025 2975
rect 15025 2941 15059 2975
rect 15059 2941 15068 2975
rect 15016 2932 15068 2941
rect 15200 2932 15252 2984
rect 16488 2975 16540 2984
rect 16488 2941 16497 2975
rect 16497 2941 16531 2975
rect 16531 2941 16540 2975
rect 16488 2932 16540 2941
rect 16764 2975 16816 2984
rect 16764 2941 16773 2975
rect 16773 2941 16807 2975
rect 16807 2941 16816 2975
rect 16764 2932 16816 2941
rect 14924 2839 14976 2848
rect 14924 2805 14933 2839
rect 14933 2805 14967 2839
rect 14967 2805 14976 2839
rect 14924 2796 14976 2805
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 6571 2694 6623 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 11904 2694 11956 2746
rect 11968 2694 12020 2746
rect 2136 2592 2188 2644
rect 7104 2635 7156 2644
rect 1584 2567 1636 2576
rect 1584 2533 1593 2567
rect 1593 2533 1627 2567
rect 1627 2533 1636 2567
rect 1584 2524 1636 2533
rect 7104 2601 7113 2635
rect 7113 2601 7147 2635
rect 7147 2601 7156 2635
rect 7104 2592 7156 2601
rect 7380 2635 7432 2644
rect 7380 2601 7389 2635
rect 7389 2601 7423 2635
rect 7423 2601 7432 2635
rect 7380 2592 7432 2601
rect 8392 2592 8444 2644
rect 9680 2635 9732 2644
rect 9680 2601 9689 2635
rect 9689 2601 9723 2635
rect 9723 2601 9732 2635
rect 9680 2592 9732 2601
rect 10416 2592 10468 2644
rect 11060 2592 11112 2644
rect 13636 2635 13688 2644
rect 13636 2601 13645 2635
rect 13645 2601 13679 2635
rect 13679 2601 13688 2635
rect 13636 2592 13688 2601
rect 14188 2592 14240 2644
rect 14924 2635 14976 2644
rect 1676 2456 1728 2508
rect 2044 2499 2096 2508
rect 2044 2465 2053 2499
rect 2053 2465 2087 2499
rect 2087 2465 2096 2499
rect 2044 2456 2096 2465
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 2780 2456 2832 2465
rect 1400 2363 1452 2372
rect 1400 2329 1409 2363
rect 1409 2329 1443 2363
rect 1443 2329 1452 2363
rect 1400 2320 1452 2329
rect 4160 2499 4212 2508
rect 4160 2465 4169 2499
rect 4169 2465 4203 2499
rect 4203 2465 4212 2499
rect 4160 2456 4212 2465
rect 4804 2456 4856 2508
rect 5448 2456 5500 2508
rect 5540 2456 5592 2508
rect 12992 2524 13044 2576
rect 14924 2601 14933 2635
rect 14933 2601 14967 2635
rect 14967 2601 14976 2635
rect 14924 2592 14976 2601
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 7288 2499 7340 2508
rect 6920 2456 6972 2465
rect 7288 2465 7297 2499
rect 7297 2465 7331 2499
rect 7331 2465 7340 2499
rect 7288 2456 7340 2465
rect 8300 2456 8352 2508
rect 9680 2456 9732 2508
rect 11060 2456 11112 2508
rect 12440 2456 12492 2508
rect 13820 2499 13872 2508
rect 13820 2465 13829 2499
rect 13829 2465 13863 2499
rect 13863 2465 13872 2499
rect 13820 2456 13872 2465
rect 13912 2456 13964 2508
rect 15568 2456 15620 2508
rect 17040 2456 17092 2508
rect 8668 2388 8720 2440
rect 12624 2388 12676 2440
rect 16580 2388 16632 2440
rect 5264 2320 5316 2372
rect 5632 2320 5684 2372
rect 10968 2320 11020 2372
rect 5448 2252 5500 2304
rect 3680 2150 3732 2202
rect 3744 2150 3796 2202
rect 3808 2150 3860 2202
rect 3872 2150 3924 2202
rect 9078 2150 9130 2202
rect 9142 2150 9194 2202
rect 9206 2150 9258 2202
rect 9270 2150 9322 2202
rect 14475 2150 14527 2202
rect 14539 2150 14591 2202
rect 14603 2150 14655 2202
rect 14667 2150 14719 2202
<< metal2 >>
rect 478 19804 534 20604
rect 1858 19804 1914 20604
rect 3238 19804 3294 20604
rect 4618 19804 4674 20604
rect 5998 19804 6054 20604
rect 7378 19804 7434 20604
rect 8758 19804 8814 20604
rect 10138 19804 10194 20604
rect 11518 19804 11574 20604
rect 12898 19804 12954 20604
rect 14278 19804 14334 20604
rect 15658 19804 15714 20604
rect 17038 19804 17094 20604
rect 492 17814 520 19804
rect 1490 18456 1546 18465
rect 1490 18391 1546 18400
rect 1504 17882 1532 18391
rect 1492 17876 1544 17882
rect 1492 17818 1544 17824
rect 480 17808 532 17814
rect 480 17750 532 17756
rect 1872 17746 1900 19804
rect 3252 17746 3280 19804
rect 4632 17746 4660 19804
rect 6012 17746 6040 19804
rect 6353 17980 6649 18000
rect 6409 17978 6433 17980
rect 6489 17978 6513 17980
rect 6569 17978 6593 17980
rect 6431 17926 6433 17978
rect 6495 17926 6507 17978
rect 6569 17926 6571 17978
rect 6409 17924 6433 17926
rect 6489 17924 6513 17926
rect 6569 17924 6593 17926
rect 6353 17904 6649 17924
rect 7392 17746 7420 19804
rect 8772 17762 8800 19804
rect 8772 17746 8892 17762
rect 10152 17746 10180 19804
rect 11532 17746 11560 19804
rect 11750 17980 12046 18000
rect 11806 17978 11830 17980
rect 11886 17978 11910 17980
rect 11966 17978 11990 17980
rect 11828 17926 11830 17978
rect 11892 17926 11904 17978
rect 11966 17926 11968 17978
rect 11806 17924 11830 17926
rect 11886 17924 11910 17926
rect 11966 17924 11990 17926
rect 11750 17904 12046 17924
rect 12912 17746 12940 19804
rect 14292 17746 14320 19804
rect 15566 19136 15622 19145
rect 15566 19071 15622 19080
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 3240 17740 3292 17746
rect 3240 17682 3292 17688
rect 4252 17740 4304 17746
rect 4252 17682 4304 17688
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 6000 17740 6052 17746
rect 6000 17682 6052 17688
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 8300 17740 8352 17746
rect 8772 17740 8904 17746
rect 8772 17734 8852 17740
rect 8300 17682 8352 17688
rect 8852 17682 8904 17688
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 1596 17338 1624 17682
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 2228 17536 2280 17542
rect 2228 17478 2280 17484
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1688 16726 1716 16934
rect 1676 16720 1728 16726
rect 1676 16662 1728 16668
rect 1780 16590 1808 17070
rect 1768 16584 1820 16590
rect 1768 16526 1820 16532
rect 1398 16416 1454 16425
rect 1398 16351 1454 16360
rect 1412 16046 1440 16351
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 1872 14890 1900 15302
rect 1860 14884 1912 14890
rect 1860 14826 1912 14832
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1412 14385 1440 14418
rect 1398 14376 1454 14385
rect 1398 14311 1454 14320
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1398 12336 1454 12345
rect 1398 12271 1400 12280
rect 1452 12271 1454 12280
rect 1400 12242 1452 12248
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1490 10296 1546 10305
rect 1490 10231 1492 10240
rect 1544 10231 1546 10240
rect 1492 10202 1544 10208
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1412 8514 1440 9318
rect 1412 8498 1532 8514
rect 1400 8492 1532 8498
rect 1452 8486 1532 8492
rect 1400 8434 1452 8440
rect 1400 8356 1452 8362
rect 1400 8298 1452 8304
rect 1412 8265 1440 8298
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1504 7954 1532 8486
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1596 6866 1624 12038
rect 1676 10532 1728 10538
rect 1676 10474 1728 10480
rect 1688 9654 1716 10474
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1780 10062 1808 10406
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1688 8634 1716 9590
rect 1872 9586 1900 14214
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 1964 12714 1992 13126
rect 1952 12708 2004 12714
rect 1952 12650 2004 12656
rect 2056 12434 2084 17478
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2148 15570 2176 17138
rect 2136 15564 2188 15570
rect 2136 15506 2188 15512
rect 2148 13394 2176 15506
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 1964 12406 2084 12434
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1688 6798 1716 8570
rect 1964 7478 1992 12406
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 2056 10130 2084 11154
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2148 10810 2176 11086
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2240 10674 2268 17478
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2596 17128 2648 17134
rect 2596 17070 2648 17076
rect 2608 16794 2636 17070
rect 2596 16788 2648 16794
rect 2596 16730 2648 16736
rect 2792 14822 2820 17274
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2884 15065 2912 17070
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 3068 16726 3096 16934
rect 3056 16720 3108 16726
rect 3056 16662 3108 16668
rect 2964 15632 3016 15638
rect 2964 15574 3016 15580
rect 2870 15056 2926 15065
rect 2870 14991 2926 15000
rect 2780 14816 2832 14822
rect 2780 14758 2832 14764
rect 2976 14550 3004 15574
rect 3148 15564 3200 15570
rect 3148 15506 3200 15512
rect 3160 15162 3188 15506
rect 3148 15156 3200 15162
rect 3148 15098 3200 15104
rect 3160 14929 3188 15098
rect 3146 14920 3202 14929
rect 3146 14855 3202 14864
rect 2964 14544 3016 14550
rect 2964 14486 3016 14492
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 2332 9602 2360 13942
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2700 10606 2728 11290
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 3068 10810 3096 11018
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2872 10532 2924 10538
rect 2872 10474 2924 10480
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2608 9926 2636 10406
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2792 9722 2820 10066
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 2148 9574 2360 9602
rect 2044 8356 2096 8362
rect 2044 8298 2096 8304
rect 1952 7472 2004 7478
rect 1952 7414 2004 7420
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1688 6322 1716 6734
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1398 6216 1454 6225
rect 1398 6151 1454 6160
rect 1412 5778 1440 6151
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5914 1624 6054
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1398 4176 1454 4185
rect 2056 4146 2084 8298
rect 1398 4111 1400 4120
rect 1452 4111 1454 4120
rect 2044 4140 2096 4146
rect 1400 4082 1452 4088
rect 2044 4082 2096 4088
rect 1584 4004 1636 4010
rect 1584 3946 1636 3952
rect 1596 3602 1624 3946
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 480 2984 532 2990
rect 480 2926 532 2932
rect 492 800 520 2926
rect 1596 2582 1624 2994
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1584 2576 1636 2582
rect 1584 2518 1636 2524
rect 1688 2514 1716 2790
rect 2148 2650 2176 9574
rect 2320 9444 2372 9450
rect 2320 9386 2372 9392
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2240 8566 2268 8774
rect 2228 8560 2280 8566
rect 2228 8502 2280 8508
rect 2332 8294 2360 9386
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 2332 8022 2360 8230
rect 2320 8016 2372 8022
rect 2320 7958 2372 7964
rect 2516 7954 2544 8366
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2516 7546 2544 7890
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2516 6730 2544 7210
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2332 4740 2360 6054
rect 2424 5302 2452 6598
rect 2516 6186 2544 6666
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 2412 5296 2464 5302
rect 2412 5238 2464 5244
rect 2424 5166 2452 5238
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2332 4712 2452 4740
rect 2424 4622 2452 4712
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2516 4434 2544 6122
rect 2884 5166 2912 10474
rect 3056 9988 3108 9994
rect 3056 9930 3108 9936
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2976 8362 3004 8978
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 2872 5160 2924 5166
rect 2924 5120 3004 5148
rect 2872 5102 2924 5108
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2424 4406 2544 4434
rect 2424 2990 2452 4406
rect 2792 3670 2820 4762
rect 2884 4758 2912 4966
rect 2872 4752 2924 4758
rect 2872 4694 2924 4700
rect 2976 4690 3004 5120
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 3068 3040 3096 9930
rect 3252 8906 3280 17478
rect 3654 17436 3950 17456
rect 3710 17434 3734 17436
rect 3790 17434 3814 17436
rect 3870 17434 3894 17436
rect 3732 17382 3734 17434
rect 3796 17382 3808 17434
rect 3870 17382 3872 17434
rect 3710 17380 3734 17382
rect 3790 17380 3814 17382
rect 3870 17380 3894 17382
rect 3654 17360 3950 17380
rect 4264 17338 4292 17682
rect 7564 17604 7616 17610
rect 7564 17546 7616 17552
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 4528 17536 4580 17542
rect 4528 17478 4580 17484
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 3424 17128 3476 17134
rect 3476 17088 3556 17116
rect 3424 17070 3476 17076
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 3436 16658 3464 16934
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 3436 16454 3464 16594
rect 3528 16590 3556 17088
rect 4264 16794 4292 17274
rect 4448 17066 4476 17478
rect 4436 17060 4488 17066
rect 4436 17002 4488 17008
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 3344 15094 3372 15506
rect 3436 15434 3464 16390
rect 3528 16046 3556 16526
rect 3654 16348 3950 16368
rect 3710 16346 3734 16348
rect 3790 16346 3814 16348
rect 3870 16346 3894 16348
rect 3732 16294 3734 16346
rect 3796 16294 3808 16346
rect 3870 16294 3872 16346
rect 3710 16292 3734 16294
rect 3790 16292 3814 16294
rect 3870 16292 3894 16294
rect 3654 16272 3950 16292
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 4436 15972 4488 15978
rect 4436 15914 4488 15920
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 3424 15428 3476 15434
rect 3424 15370 3476 15376
rect 3332 15088 3384 15094
rect 3332 15030 3384 15036
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3344 14618 3372 14894
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3436 14550 3464 15370
rect 3528 14890 3556 15642
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 3654 15260 3950 15280
rect 3710 15258 3734 15260
rect 3790 15258 3814 15260
rect 3870 15258 3894 15260
rect 3732 15206 3734 15258
rect 3796 15206 3808 15258
rect 3870 15206 3872 15258
rect 3710 15204 3734 15206
rect 3790 15204 3814 15206
rect 3870 15204 3894 15206
rect 3654 15184 3950 15204
rect 3882 15056 3938 15065
rect 3882 14991 3938 15000
rect 3896 14958 3924 14991
rect 3700 14952 3752 14958
rect 3698 14920 3700 14929
rect 3884 14952 3936 14958
rect 3752 14920 3754 14929
rect 3516 14884 3568 14890
rect 3884 14894 3936 14900
rect 4080 14890 4108 15370
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 3698 14855 3754 14864
rect 4068 14884 4120 14890
rect 3516 14826 3568 14832
rect 4068 14826 4120 14832
rect 3424 14544 3476 14550
rect 3424 14486 3476 14492
rect 3332 14476 3384 14482
rect 3332 14418 3384 14424
rect 3344 12850 3372 14418
rect 3528 14414 3556 14826
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3712 14482 3740 14758
rect 3700 14476 3752 14482
rect 3700 14418 3752 14424
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3528 13870 3556 14214
rect 3654 14172 3950 14192
rect 3710 14170 3734 14172
rect 3790 14170 3814 14172
rect 3870 14170 3894 14172
rect 3732 14118 3734 14170
rect 3796 14118 3808 14170
rect 3870 14118 3872 14170
rect 3710 14116 3734 14118
rect 3790 14116 3814 14118
rect 3870 14116 3894 14118
rect 3654 14096 3950 14116
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3424 13728 3476 13734
rect 3424 13670 3476 13676
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3344 10674 3372 12786
rect 3436 12714 3464 13670
rect 3528 13462 3556 13806
rect 4080 13734 4108 14826
rect 4172 14482 4200 15302
rect 4252 15088 4304 15094
rect 4252 15030 4304 15036
rect 4264 14618 4292 15030
rect 4356 15026 4384 15438
rect 4448 15162 4476 15914
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4264 13530 4292 14554
rect 4448 14550 4476 15098
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4344 14476 4396 14482
rect 4344 14418 4396 14424
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 3516 13456 3568 13462
rect 3516 13398 3568 13404
rect 4068 13388 4120 13394
rect 4252 13388 4304 13394
rect 4068 13330 4120 13336
rect 4172 13348 4252 13376
rect 4080 13297 4108 13330
rect 4066 13288 4122 13297
rect 3976 13252 4028 13258
rect 4066 13223 4122 13232
rect 3976 13194 4028 13200
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3528 12782 3556 13126
rect 3654 13084 3950 13104
rect 3710 13082 3734 13084
rect 3790 13082 3814 13084
rect 3870 13082 3894 13084
rect 3732 13030 3734 13082
rect 3796 13030 3808 13082
rect 3870 13030 3872 13082
rect 3710 13028 3734 13030
rect 3790 13028 3814 13030
rect 3870 13028 3894 13030
rect 3654 13008 3950 13028
rect 3988 12918 4016 13194
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 3976 12912 4028 12918
rect 3882 12880 3938 12889
rect 3976 12854 4028 12860
rect 3882 12815 3938 12824
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3896 12714 3924 12815
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3896 12084 3924 12650
rect 3988 12238 4016 12854
rect 4080 12782 4108 13126
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 4172 12306 4200 13348
rect 4252 13330 4304 13336
rect 4356 13326 4384 14418
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4264 12850 4292 13126
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4356 12782 4384 13262
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 3896 12056 4016 12084
rect 3654 11996 3950 12016
rect 3710 11994 3734 11996
rect 3790 11994 3814 11996
rect 3870 11994 3894 11996
rect 3732 11942 3734 11994
rect 3796 11942 3808 11994
rect 3870 11942 3872 11994
rect 3710 11940 3734 11942
rect 3790 11940 3814 11942
rect 3870 11940 3894 11942
rect 3654 11920 3950 11940
rect 3654 10908 3950 10928
rect 3710 10906 3734 10908
rect 3790 10906 3814 10908
rect 3870 10906 3894 10908
rect 3732 10854 3734 10906
rect 3796 10854 3808 10906
rect 3870 10854 3872 10906
rect 3710 10852 3734 10854
rect 3790 10852 3814 10854
rect 3870 10852 3894 10854
rect 3654 10832 3950 10852
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3620 10266 3648 10406
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3654 9820 3950 9840
rect 3710 9818 3734 9820
rect 3790 9818 3814 9820
rect 3870 9818 3894 9820
rect 3732 9766 3734 9818
rect 3796 9766 3808 9818
rect 3870 9766 3872 9818
rect 3710 9764 3734 9766
rect 3790 9764 3814 9766
rect 3870 9764 3894 9766
rect 3654 9744 3950 9764
rect 3988 9518 4016 12056
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 4172 9382 4200 12242
rect 4264 11694 4292 12242
rect 4356 12238 4384 12718
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4448 11898 4476 13670
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4448 11744 4476 11834
rect 4356 11716 4476 11744
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4356 11218 4384 11716
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4448 11150 4476 11494
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4448 10674 4476 10950
rect 4436 10668 4488 10674
rect 4436 10610 4488 10616
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 3240 8900 3292 8906
rect 3240 8842 3292 8848
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3654 8732 3950 8752
rect 3710 8730 3734 8732
rect 3790 8730 3814 8732
rect 3870 8730 3894 8732
rect 3732 8678 3734 8730
rect 3796 8678 3808 8730
rect 3870 8678 3872 8730
rect 3710 8676 3734 8678
rect 3790 8676 3814 8678
rect 3870 8676 3894 8678
rect 3654 8656 3950 8676
rect 3654 7644 3950 7664
rect 3710 7642 3734 7644
rect 3790 7642 3814 7644
rect 3870 7642 3894 7644
rect 3732 7590 3734 7642
rect 3796 7590 3808 7642
rect 3870 7590 3872 7642
rect 3710 7588 3734 7590
rect 3790 7588 3814 7590
rect 3870 7588 3894 7590
rect 3654 7568 3950 7588
rect 3988 6866 4016 8774
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4172 7410 4200 8230
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4172 6866 4200 7346
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 3654 6556 3950 6576
rect 3710 6554 3734 6556
rect 3790 6554 3814 6556
rect 3870 6554 3894 6556
rect 3732 6502 3734 6554
rect 3796 6502 3808 6554
rect 3870 6502 3872 6554
rect 3710 6500 3734 6502
rect 3790 6500 3814 6502
rect 3870 6500 3894 6502
rect 3654 6480 3950 6500
rect 3988 6254 4016 6802
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 4264 5846 4292 9454
rect 4540 8498 4568 17478
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4816 15978 4844 16390
rect 4804 15972 4856 15978
rect 4804 15914 4856 15920
rect 4896 15904 4948 15910
rect 4816 15852 4896 15858
rect 4816 15846 4948 15852
rect 4816 15830 4936 15846
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4724 15065 4752 15506
rect 4710 15056 4766 15065
rect 4632 15014 4710 15042
rect 4632 13190 4660 15014
rect 4710 14991 4766 15000
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 4724 13462 4752 13806
rect 4712 13456 4764 13462
rect 4712 13398 4764 13404
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4632 11694 4660 12854
rect 4724 12850 4752 13398
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4724 11694 4752 12038
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4712 10532 4764 10538
rect 4712 10474 4764 10480
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4632 8294 4660 9522
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4448 6934 4476 7142
rect 4436 6928 4488 6934
rect 4436 6870 4488 6876
rect 4252 5840 4304 5846
rect 4252 5782 4304 5788
rect 3654 5468 3950 5488
rect 3710 5466 3734 5468
rect 3790 5466 3814 5468
rect 3870 5466 3894 5468
rect 3732 5414 3734 5466
rect 3796 5414 3808 5466
rect 3870 5414 3872 5466
rect 3710 5412 3734 5414
rect 3790 5412 3814 5414
rect 3870 5412 3894 5414
rect 3654 5392 3950 5412
rect 4264 5234 4292 5782
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4264 4758 4292 5170
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 3654 4380 3950 4400
rect 3710 4378 3734 4380
rect 3790 4378 3814 4380
rect 3870 4378 3894 4380
rect 3732 4326 3734 4378
rect 3796 4326 3808 4378
rect 3870 4326 3872 4378
rect 3710 4324 3734 4326
rect 3790 4324 3814 4326
rect 3870 4324 3894 4326
rect 3654 4304 3950 4324
rect 4172 4078 4200 4422
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4724 4010 4752 10474
rect 4816 5914 4844 15830
rect 5460 14958 5488 16730
rect 6288 16726 6316 16934
rect 6353 16892 6649 16912
rect 6409 16890 6433 16892
rect 6489 16890 6513 16892
rect 6569 16890 6593 16892
rect 6431 16838 6433 16890
rect 6495 16838 6507 16890
rect 6569 16838 6571 16890
rect 6409 16836 6433 16838
rect 6489 16836 6513 16838
rect 6569 16836 6593 16838
rect 6353 16816 6649 16836
rect 6276 16720 6328 16726
rect 6276 16662 6328 16668
rect 6748 16114 6776 17138
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 6460 16040 6512 16046
rect 6840 15994 6868 16934
rect 7024 16250 7052 17070
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7024 16046 7052 16186
rect 6512 15988 6868 15994
rect 6460 15982 6868 15988
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 6472 15966 6868 15982
rect 6353 15804 6649 15824
rect 6409 15802 6433 15804
rect 6489 15802 6513 15804
rect 6569 15802 6593 15804
rect 6431 15750 6433 15802
rect 6495 15750 6507 15802
rect 6569 15750 6571 15802
rect 6409 15748 6433 15750
rect 6489 15748 6513 15750
rect 6569 15748 6593 15750
rect 6353 15728 6649 15748
rect 6840 15094 6868 15966
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 5448 14952 5500 14958
rect 5368 14912 5448 14940
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5276 14074 5304 14350
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 4908 12782 4936 13330
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 5000 11694 5028 13126
rect 5080 11824 5132 11830
rect 5080 11766 5132 11772
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 5092 9178 5120 11766
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5184 11354 5212 11630
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 5184 10266 5212 10474
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5368 10130 5396 14912
rect 5448 14894 5500 14900
rect 7024 14890 7052 15982
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 5552 14550 5580 14758
rect 6353 14716 6649 14736
rect 6409 14714 6433 14716
rect 6489 14714 6513 14716
rect 6569 14714 6593 14716
rect 6431 14662 6433 14714
rect 6495 14662 6507 14714
rect 6569 14662 6571 14714
rect 6409 14660 6433 14662
rect 6489 14660 6513 14662
rect 6569 14660 6593 14662
rect 6353 14640 6649 14660
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5828 13802 5856 14214
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 6000 13864 6052 13870
rect 6052 13812 6132 13818
rect 6000 13806 6132 13812
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5816 13796 5868 13802
rect 5816 13738 5868 13744
rect 5552 13530 5580 13738
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5460 12782 5488 13466
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5460 11082 5488 12718
rect 5828 12714 5856 13738
rect 5920 13190 5948 13806
rect 6012 13790 6132 13806
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6012 13394 6040 13670
rect 6104 13394 6132 13790
rect 6353 13628 6649 13648
rect 6409 13626 6433 13628
rect 6489 13626 6513 13628
rect 6569 13626 6593 13628
rect 6431 13574 6433 13626
rect 6495 13574 6507 13626
rect 6569 13574 6571 13626
rect 6409 13572 6433 13574
rect 6489 13572 6513 13574
rect 6569 13572 6593 13574
rect 6353 13552 6649 13572
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5920 12889 5948 13126
rect 5906 12880 5962 12889
rect 5906 12815 5962 12824
rect 5816 12708 5868 12714
rect 5816 12650 5868 12656
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 11218 5580 12174
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5736 10810 5764 11154
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5184 9110 5212 9318
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5172 8968 5224 8974
rect 5276 8956 5304 9454
rect 5368 9382 5396 10066
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5224 8928 5304 8956
rect 5172 8910 5224 8916
rect 5092 8634 5120 8910
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5184 8566 5212 8910
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 5184 7886 5212 8502
rect 5644 8498 5672 9386
rect 5736 9042 5764 10746
rect 5828 10130 5856 12650
rect 6012 12646 6040 13330
rect 6552 13252 6604 13258
rect 6552 13194 6604 13200
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 6196 12238 6224 13126
rect 6564 12918 6592 13194
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5920 10470 5948 10950
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5828 8838 5856 10066
rect 5920 9722 5948 10406
rect 6288 10266 6316 12786
rect 6564 12730 6592 12854
rect 6748 12850 6776 13330
rect 6840 13326 6868 14758
rect 7024 14550 7052 14826
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6840 12918 6868 13262
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6564 12702 6776 12730
rect 6353 12540 6649 12560
rect 6409 12538 6433 12540
rect 6489 12538 6513 12540
rect 6569 12538 6593 12540
rect 6431 12486 6433 12538
rect 6495 12486 6507 12538
rect 6569 12486 6571 12538
rect 6409 12484 6433 12486
rect 6489 12484 6513 12486
rect 6569 12484 6593 12486
rect 6353 12464 6649 12484
rect 6748 12374 6776 12702
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6840 12306 6868 12582
rect 7024 12434 7052 12922
rect 6932 12406 7052 12434
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6353 11452 6649 11472
rect 6409 11450 6433 11452
rect 6489 11450 6513 11452
rect 6569 11450 6593 11452
rect 6431 11398 6433 11450
rect 6495 11398 6507 11450
rect 6569 11398 6571 11450
rect 6409 11396 6433 11398
rect 6489 11396 6513 11398
rect 6569 11396 6593 11398
rect 6353 11376 6649 11396
rect 6840 11354 6868 11630
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6353 10364 6649 10384
rect 6409 10362 6433 10364
rect 6489 10362 6513 10364
rect 6569 10362 6593 10364
rect 6431 10310 6433 10362
rect 6495 10310 6507 10362
rect 6569 10310 6571 10362
rect 6409 10308 6433 10310
rect 6489 10308 6513 10310
rect 6569 10308 6593 10310
rect 6353 10288 6649 10308
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6748 10146 6776 10950
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6564 10118 6776 10146
rect 6564 10062 6592 10118
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6012 9518 6040 9590
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5828 8650 5856 8774
rect 5736 8622 5856 8650
rect 5736 8566 5764 8622
rect 6104 8566 6132 8978
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 6092 8560 6144 8566
rect 6092 8502 6144 8508
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5644 8106 5672 8434
rect 5724 8424 5776 8430
rect 6000 8424 6052 8430
rect 5724 8366 5776 8372
rect 5998 8392 6000 8401
rect 6052 8392 6054 8401
rect 5552 8078 5672 8106
rect 5552 7954 5580 8078
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4908 6866 4936 7142
rect 5000 6934 5028 7210
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4908 6186 4936 6802
rect 5092 6730 5120 7278
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 4896 6180 4948 6186
rect 4896 6122 4948 6128
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 3654 3292 3950 3312
rect 3710 3290 3734 3292
rect 3790 3290 3814 3292
rect 3870 3290 3894 3292
rect 3732 3238 3734 3290
rect 3796 3238 3808 3290
rect 3870 3238 3872 3290
rect 3710 3236 3734 3238
rect 3790 3236 3814 3238
rect 3870 3236 3894 3238
rect 3654 3216 3950 3236
rect 3148 3052 3200 3058
rect 3068 3012 3148 3040
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 3068 2922 3096 3012
rect 3148 2994 3200 3000
rect 3056 2916 3108 2922
rect 3056 2858 3108 2864
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 4816 2514 4844 5714
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 5092 4826 5120 5034
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5276 2854 5304 3606
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 1400 2372 1452 2378
rect 1400 2314 1452 2320
rect 1412 800 1440 2314
rect 2056 2145 2084 2450
rect 2042 2136 2098 2145
rect 2042 2071 2098 2080
rect 2792 800 2820 2450
rect 3654 2204 3950 2224
rect 3710 2202 3734 2204
rect 3790 2202 3814 2204
rect 3870 2202 3894 2204
rect 3732 2150 3734 2202
rect 3796 2150 3808 2202
rect 3870 2150 3872 2202
rect 3710 2148 3734 2150
rect 3790 2148 3814 2150
rect 3870 2148 3894 2150
rect 3654 2128 3950 2148
rect 4172 800 4200 2450
rect 5276 2378 5304 2790
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 5460 2310 5488 2450
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5552 800 5580 2450
rect 5644 2378 5672 7958
rect 5736 6798 5764 8366
rect 5816 8356 5868 8362
rect 5998 8327 6054 8336
rect 5816 8298 5868 8304
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5828 6254 5856 8298
rect 6104 8090 6132 8502
rect 6196 8294 6224 9590
rect 6288 9518 6316 9998
rect 6564 9654 6592 9998
rect 6840 9722 6868 10202
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6748 9450 6776 9658
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6353 9276 6649 9296
rect 6409 9274 6433 9276
rect 6489 9274 6513 9276
rect 6569 9274 6593 9276
rect 6431 9222 6433 9274
rect 6495 9222 6507 9274
rect 6569 9222 6571 9274
rect 6409 9220 6433 9222
rect 6489 9220 6513 9222
rect 6569 9220 6593 9222
rect 6353 9200 6649 9220
rect 6748 8922 6776 9386
rect 6840 9042 6868 9658
rect 6932 9654 6960 12406
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7024 11694 7052 12038
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7024 10130 7052 10406
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6932 9110 6960 9318
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6748 8894 6868 8922
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6184 8288 6236 8294
rect 6236 8248 6316 8276
rect 6184 8230 6236 8236
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5828 5166 5856 6190
rect 5920 6186 5948 7822
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 6012 6390 6040 6598
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 5908 6180 5960 6186
rect 5908 6122 5960 6128
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6012 4690 6040 4966
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6104 3602 6132 7414
rect 6196 7342 6224 7754
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6288 6866 6316 8248
rect 6353 8188 6649 8208
rect 6409 8186 6433 8188
rect 6489 8186 6513 8188
rect 6569 8186 6593 8188
rect 6431 8134 6433 8186
rect 6495 8134 6507 8186
rect 6569 8134 6571 8186
rect 6409 8132 6433 8134
rect 6489 8132 6513 8134
rect 6569 8132 6593 8134
rect 6353 8112 6649 8132
rect 6748 8022 6776 8366
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6840 7886 6868 8894
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6353 7100 6649 7120
rect 6409 7098 6433 7100
rect 6489 7098 6513 7100
rect 6569 7098 6593 7100
rect 6431 7046 6433 7098
rect 6495 7046 6507 7098
rect 6569 7046 6571 7098
rect 6409 7044 6433 7046
rect 6489 7044 6513 7046
rect 6569 7044 6593 7046
rect 6353 7024 6649 7044
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6840 6730 6868 7822
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 7410 6960 7686
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 7116 6118 7144 17478
rect 7288 17060 7340 17066
rect 7288 17002 7340 17008
rect 7300 16454 7328 17002
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7300 16182 7328 16390
rect 7288 16176 7340 16182
rect 7288 16118 7340 16124
rect 7300 16046 7328 16118
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7576 15570 7604 17546
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 7852 16658 7880 16730
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 8036 16590 8064 17070
rect 8312 16658 8340 17682
rect 8576 17604 8628 17610
rect 8576 17546 8628 17552
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7208 15026 7236 15506
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 7300 15162 7328 15438
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7300 14618 7328 15098
rect 7576 14890 7604 15506
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7852 14482 7880 15438
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 7852 13530 7880 14418
rect 8036 14346 8064 16526
rect 8392 15972 8444 15978
rect 8392 15914 8444 15920
rect 8404 15570 8432 15914
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 8128 14958 8156 15438
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8496 14958 8524 15302
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8024 14340 8076 14346
rect 8024 14282 8076 14288
rect 8128 14074 8156 14894
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7380 13252 7432 13258
rect 7380 13194 7432 13200
rect 7194 12880 7250 12889
rect 7194 12815 7250 12824
rect 7208 12782 7236 12815
rect 7392 12782 7420 13194
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7484 12714 7512 13330
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7576 12782 7604 13126
rect 7668 12782 7696 13330
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7484 12442 7512 12650
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7300 12306 7328 12378
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7208 11354 7236 11630
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7208 9382 7236 9522
rect 7300 9518 7328 12106
rect 7392 10470 7420 12174
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7484 11082 7512 12038
rect 8128 11898 8156 12786
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8220 12442 8248 12718
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8220 12306 8248 12378
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7760 11150 7788 11494
rect 8128 11150 8156 11834
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7392 8974 7420 10406
rect 8220 10198 8248 10406
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8312 9994 8340 11154
rect 8588 10674 8616 17546
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 10416 17536 10468 17542
rect 10416 17478 10468 17484
rect 8956 17066 8984 17478
rect 9052 17436 9348 17456
rect 9108 17434 9132 17436
rect 9188 17434 9212 17436
rect 9268 17434 9292 17436
rect 9130 17382 9132 17434
rect 9194 17382 9206 17434
rect 9268 17382 9270 17434
rect 9108 17380 9132 17382
rect 9188 17380 9212 17382
rect 9268 17380 9292 17382
rect 9052 17360 9348 17380
rect 8944 17060 8996 17066
rect 8944 17002 8996 17008
rect 9052 16348 9348 16368
rect 9108 16346 9132 16348
rect 9188 16346 9212 16348
rect 9268 16346 9292 16348
rect 9130 16294 9132 16346
rect 9194 16294 9206 16346
rect 9268 16294 9270 16346
rect 9108 16292 9132 16294
rect 9188 16292 9212 16294
rect 9268 16292 9292 16294
rect 9052 16272 9348 16292
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 8864 15638 8892 15846
rect 8852 15632 8904 15638
rect 8772 15592 8852 15620
rect 8668 14952 8720 14958
rect 8772 14906 8800 15592
rect 8852 15574 8904 15580
rect 9784 15570 9812 15846
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9052 15260 9348 15280
rect 9108 15258 9132 15260
rect 9188 15258 9212 15260
rect 9268 15258 9292 15260
rect 9130 15206 9132 15258
rect 9194 15206 9206 15258
rect 9268 15206 9270 15258
rect 9108 15204 9132 15206
rect 9188 15204 9212 15206
rect 9268 15204 9292 15206
rect 9052 15184 9348 15204
rect 9508 15026 9536 15370
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 8720 14900 8800 14906
rect 8668 14894 8800 14900
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 8680 14878 8800 14894
rect 8864 14074 8892 14894
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9052 14172 9348 14192
rect 9108 14170 9132 14172
rect 9188 14170 9212 14172
rect 9268 14170 9292 14172
rect 9130 14118 9132 14170
rect 9194 14118 9206 14170
rect 9268 14118 9270 14170
rect 9108 14116 9132 14118
rect 9188 14116 9212 14118
rect 9268 14116 9292 14118
rect 9052 14096 9348 14116
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 9052 13084 9348 13104
rect 9108 13082 9132 13084
rect 9188 13082 9212 13084
rect 9268 13082 9292 13084
rect 9130 13030 9132 13082
rect 9194 13030 9206 13082
rect 9268 13030 9270 13082
rect 9108 13028 9132 13030
rect 9188 13028 9212 13030
rect 9268 13028 9292 13030
rect 9052 13008 9348 13028
rect 9312 12844 9364 12850
rect 9416 12832 9444 14282
rect 9364 12804 9444 12832
rect 9312 12786 9364 12792
rect 9324 12152 9352 12786
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9416 12306 9444 12582
rect 9692 12442 9720 12718
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 9404 12164 9456 12170
rect 9324 12124 9404 12152
rect 9404 12106 9456 12112
rect 9052 11996 9348 12016
rect 9108 11994 9132 11996
rect 9188 11994 9212 11996
rect 9268 11994 9292 11996
rect 9130 11942 9132 11994
rect 9194 11942 9206 11994
rect 9268 11942 9270 11994
rect 9108 11940 9132 11942
rect 9188 11940 9212 11942
rect 9268 11940 9292 11942
rect 9052 11920 9348 11940
rect 9416 11150 9444 12106
rect 9508 11694 9536 12242
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9052 10908 9348 10928
rect 9108 10906 9132 10908
rect 9188 10906 9212 10908
rect 9268 10906 9292 10908
rect 9130 10854 9132 10906
rect 9194 10854 9206 10906
rect 9268 10854 9270 10906
rect 9108 10852 9132 10854
rect 9188 10852 9212 10854
rect 9268 10852 9292 10854
rect 9052 10832 9348 10852
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9140 10266 9168 10406
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9416 9994 9444 10406
rect 9600 10282 9628 12310
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9692 11286 9720 11494
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9508 10266 9628 10282
rect 9508 10260 9640 10266
rect 9508 10254 9588 10260
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 9404 9988 9456 9994
rect 9404 9930 9456 9936
rect 7840 9648 7892 9654
rect 7840 9590 7892 9596
rect 7564 9512 7616 9518
rect 7562 9480 7564 9489
rect 7616 9480 7618 9489
rect 7562 9415 7618 9424
rect 7746 9480 7802 9489
rect 7746 9415 7802 9424
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7392 7954 7420 8434
rect 7576 8430 7604 8910
rect 7668 8430 7696 8978
rect 7760 8498 7788 9415
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7852 8430 7880 9590
rect 7944 9574 8156 9602
rect 7944 9518 7972 9574
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 8036 9178 8064 9454
rect 8128 9178 8156 9574
rect 8312 9489 8340 9930
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8298 9480 8354 9489
rect 8298 9415 8354 9424
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7564 8424 7616 8430
rect 7656 8424 7708 8430
rect 7564 8366 7616 8372
rect 7654 8392 7656 8401
rect 7840 8424 7892 8430
rect 7708 8392 7710 8401
rect 7840 8366 7892 8372
rect 7654 8327 7710 8336
rect 7944 7954 7972 8434
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7392 6662 7420 7278
rect 7668 6866 7696 7346
rect 7852 6866 7880 7414
rect 8036 7342 8064 9114
rect 8128 8242 8156 9114
rect 8220 8974 8248 9114
rect 8312 9042 8340 9415
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8220 8566 8248 8910
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8128 8214 8248 8242
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7300 6254 7328 6598
rect 7392 6322 7420 6598
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 6353 6012 6649 6032
rect 6409 6010 6433 6012
rect 6489 6010 6513 6012
rect 6569 6010 6593 6012
rect 6431 5958 6433 6010
rect 6495 5958 6507 6010
rect 6569 5958 6571 6010
rect 6409 5956 6433 5958
rect 6489 5956 6513 5958
rect 6569 5956 6593 5958
rect 6353 5936 6649 5956
rect 6353 4924 6649 4944
rect 6409 4922 6433 4924
rect 6489 4922 6513 4924
rect 6569 4922 6593 4924
rect 6431 4870 6433 4922
rect 6495 4870 6507 4922
rect 6569 4870 6571 4922
rect 6409 4868 6433 4870
rect 6489 4868 6513 4870
rect 6569 4868 6593 4870
rect 6353 4848 6649 4868
rect 6840 4622 6868 6054
rect 7392 5234 7420 6258
rect 7484 6254 7512 6802
rect 7668 6458 7696 6802
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7852 6322 7880 6802
rect 8024 6792 8076 6798
rect 8128 6780 8156 7822
rect 8220 7410 8248 8214
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 7410 8340 7686
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8404 7342 8432 9318
rect 8864 8498 8892 9862
rect 9052 9820 9348 9840
rect 9108 9818 9132 9820
rect 9188 9818 9212 9820
rect 9268 9818 9292 9820
rect 9130 9766 9132 9818
rect 9194 9766 9206 9818
rect 9268 9766 9270 9818
rect 9108 9764 9132 9766
rect 9188 9764 9212 9766
rect 9268 9764 9292 9766
rect 9052 9744 9348 9764
rect 9416 9722 9444 9930
rect 9404 9716 9456 9722
rect 9324 9664 9404 9674
rect 9324 9658 9456 9664
rect 9324 9646 9444 9658
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8392 7336 8444 7342
rect 8444 7296 8524 7324
rect 8392 7278 8444 7284
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8312 7002 8340 7142
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8496 6934 8524 7296
rect 8772 7274 8800 8230
rect 8852 7540 8904 7546
rect 8956 7528 8984 9046
rect 9048 9042 9076 9522
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9232 9110 9260 9454
rect 9220 9104 9272 9110
rect 9220 9046 9272 9052
rect 9324 9042 9352 9646
rect 9416 9593 9444 9646
rect 9508 9586 9536 10254
rect 9588 10202 9640 10208
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9416 9382 9444 9454
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9508 8974 9536 9386
rect 9600 9042 9628 10066
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9692 9024 9720 9862
rect 9772 9036 9824 9042
rect 9692 8996 9772 9024
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9052 8732 9348 8752
rect 9108 8730 9132 8732
rect 9188 8730 9212 8732
rect 9268 8730 9292 8732
rect 9130 8678 9132 8730
rect 9194 8678 9206 8730
rect 9268 8678 9270 8730
rect 9108 8676 9132 8678
rect 9188 8676 9212 8678
rect 9268 8676 9292 8678
rect 9052 8656 9348 8676
rect 9404 8560 9456 8566
rect 9404 8502 9456 8508
rect 9052 7644 9348 7664
rect 9108 7642 9132 7644
rect 9188 7642 9212 7644
rect 9268 7642 9292 7644
rect 9130 7590 9132 7642
rect 9194 7590 9206 7642
rect 9268 7590 9270 7642
rect 9108 7588 9132 7590
rect 9188 7588 9212 7590
rect 9268 7588 9292 7590
rect 9052 7568 9348 7588
rect 8904 7500 8984 7528
rect 8852 7482 8904 7488
rect 8956 7274 8984 7500
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8944 7268 8996 7274
rect 8944 7210 8996 7216
rect 8484 6928 8536 6934
rect 8484 6870 8536 6876
rect 8076 6752 8156 6780
rect 8392 6792 8444 6798
rect 8024 6734 8076 6740
rect 8392 6734 8444 6740
rect 8036 6662 8064 6734
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6840 4146 6868 4558
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 7024 3942 7052 4014
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 6353 3836 6649 3856
rect 6409 3834 6433 3836
rect 6489 3834 6513 3836
rect 6569 3834 6593 3836
rect 6431 3782 6433 3834
rect 6495 3782 6507 3834
rect 6569 3782 6571 3834
rect 6409 3780 6433 3782
rect 6489 3780 6513 3782
rect 6569 3780 6593 3782
rect 6353 3760 6649 3780
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6012 3058 6040 3470
rect 6104 3058 6132 3538
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 6353 2748 6649 2768
rect 6409 2746 6433 2748
rect 6489 2746 6513 2748
rect 6569 2746 6593 2748
rect 6431 2694 6433 2746
rect 6495 2694 6507 2746
rect 6569 2694 6571 2746
rect 6409 2692 6433 2694
rect 6489 2692 6513 2694
rect 6569 2692 6593 2694
rect 6353 2672 6649 2692
rect 7116 2650 7144 5034
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 8036 4758 8064 4966
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7300 4078 7328 4626
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7392 4282 7420 4558
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7208 3534 7236 3878
rect 7300 3670 7328 4014
rect 7288 3664 7340 3670
rect 7288 3606 7340 3612
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 7300 3126 7328 3606
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7392 3194 7420 3334
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7300 2514 7328 2926
rect 7392 2650 7420 3130
rect 7484 2990 7512 3538
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7668 3194 7696 3470
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 8036 3126 8064 3470
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 8036 2990 8064 3062
rect 8128 3058 8156 5170
rect 8312 5166 8340 6054
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 8404 2650 8432 6734
rect 8772 6254 8800 7210
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8588 4622 8616 4966
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8588 3670 8616 4422
rect 8576 3664 8628 3670
rect 8576 3606 8628 3612
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 5632 2372 5684 2378
rect 5632 2314 5684 2320
rect 6932 800 6960 2450
rect 8312 800 8340 2450
rect 8680 2446 8708 4966
rect 8772 4690 8800 5034
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 8864 3058 8892 7142
rect 8956 6866 8984 7210
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 9052 6556 9348 6576
rect 9108 6554 9132 6556
rect 9188 6554 9212 6556
rect 9268 6554 9292 6556
rect 9130 6502 9132 6554
rect 9194 6502 9206 6554
rect 9268 6502 9270 6554
rect 9108 6500 9132 6502
rect 9188 6500 9212 6502
rect 9268 6500 9292 6502
rect 9052 6480 9348 6500
rect 9052 5468 9348 5488
rect 9108 5466 9132 5468
rect 9188 5466 9212 5468
rect 9268 5466 9292 5468
rect 9130 5414 9132 5466
rect 9194 5414 9206 5466
rect 9268 5414 9270 5466
rect 9108 5412 9132 5414
rect 9188 5412 9212 5414
rect 9268 5412 9292 5414
rect 9052 5392 9348 5412
rect 9416 5166 9444 8502
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9508 6798 9536 8366
rect 9600 7206 9628 8978
rect 9692 8838 9720 8996
rect 9772 8978 9824 8984
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9692 8566 9720 8774
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9692 8294 9720 8366
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9876 7274 9904 17478
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10336 16726 10364 17070
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 9968 16046 9996 16662
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10152 16046 10180 16526
rect 10428 16182 10456 17478
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10416 16176 10468 16182
rect 10416 16118 10468 16124
rect 10428 16046 10456 16118
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 10060 15706 10088 15846
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10520 14958 10548 17070
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10612 16658 10640 16934
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10704 16114 10732 16390
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10600 15972 10652 15978
rect 10600 15914 10652 15920
rect 10612 15570 10640 15914
rect 10704 15638 10732 16050
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10508 14952 10560 14958
rect 10508 14894 10560 14900
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10520 14482 10548 14758
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9968 13734 9996 13874
rect 10060 13870 10088 14214
rect 10336 14006 10364 14350
rect 10612 14346 10640 15506
rect 10980 15162 11008 17206
rect 11428 17128 11480 17134
rect 11428 17070 11480 17076
rect 11440 16658 11468 17070
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 11532 16658 11560 17002
rect 11750 16892 12046 16912
rect 11806 16890 11830 16892
rect 11886 16890 11910 16892
rect 11966 16890 11990 16892
rect 11828 16838 11830 16890
rect 11892 16838 11904 16890
rect 11966 16838 11968 16890
rect 11806 16836 11830 16838
rect 11886 16836 11910 16838
rect 11966 16836 11990 16838
rect 11750 16816 12046 16836
rect 12360 16658 12388 17682
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 12544 17066 12572 17478
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 10980 14958 11008 15098
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 10704 14414 10732 14894
rect 10784 14612 10836 14618
rect 10888 14600 10916 14894
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10836 14572 10916 14600
rect 10784 14554 10836 14560
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10416 14340 10468 14346
rect 10416 14282 10468 14288
rect 10600 14340 10652 14346
rect 10600 14282 10652 14288
rect 10428 14074 10456 14282
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10324 14000 10376 14006
rect 10324 13942 10376 13948
rect 10336 13870 10364 13942
rect 10796 13870 10824 14554
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 10060 12986 10088 13806
rect 10980 13802 11008 14758
rect 11624 14550 11652 16526
rect 11750 15804 12046 15824
rect 11806 15802 11830 15804
rect 11886 15802 11910 15804
rect 11966 15802 11990 15804
rect 11828 15750 11830 15802
rect 11892 15750 11904 15802
rect 11966 15750 11968 15802
rect 11806 15748 11830 15750
rect 11886 15748 11910 15750
rect 11966 15748 11990 15750
rect 11750 15728 12046 15748
rect 11992 15570 12204 15586
rect 12268 15570 12296 16594
rect 12636 16454 12664 16934
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12440 16040 12492 16046
rect 12492 16000 12572 16028
rect 12440 15982 12492 15988
rect 11980 15564 12204 15570
rect 12032 15558 12204 15564
rect 11980 15506 12032 15512
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 12176 15450 12204 15558
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12348 15496 12400 15502
rect 12084 14890 12112 15438
rect 12176 15422 12296 15450
rect 12348 15438 12400 15444
rect 12268 14958 12296 15422
rect 12360 15162 12388 15438
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 11750 14716 12046 14736
rect 11806 14714 11830 14716
rect 11886 14714 11910 14716
rect 11966 14714 11990 14716
rect 11828 14662 11830 14714
rect 11892 14662 11904 14714
rect 11966 14662 11968 14714
rect 11806 14660 11830 14662
rect 11886 14660 11910 14662
rect 11966 14660 11990 14662
rect 11750 14640 12046 14660
rect 12176 14550 12204 14758
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11256 12986 11284 13126
rect 11440 12986 11468 13330
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11072 11354 11100 12174
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9968 9178 9996 10610
rect 10244 10606 10272 11290
rect 11256 10810 11284 12310
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11348 11286 11376 12038
rect 11532 11626 11560 12854
rect 11624 11694 11652 14486
rect 11750 13628 12046 13648
rect 11806 13626 11830 13628
rect 11886 13626 11910 13628
rect 11966 13626 11990 13628
rect 11828 13574 11830 13626
rect 11892 13574 11904 13626
rect 11966 13574 11968 13626
rect 11806 13572 11830 13574
rect 11886 13572 11910 13574
rect 11966 13572 11990 13574
rect 11750 13552 12046 13572
rect 12268 13462 12296 14894
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 11750 12540 12046 12560
rect 11806 12538 11830 12540
rect 11886 12538 11910 12540
rect 11966 12538 11990 12540
rect 11828 12486 11830 12538
rect 11892 12486 11904 12538
rect 11966 12486 11968 12538
rect 11806 12484 11830 12486
rect 11886 12484 11910 12486
rect 11966 12484 11990 12486
rect 11750 12464 12046 12484
rect 12084 12102 12112 12718
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 12268 11762 12296 13398
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11532 11286 11560 11562
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11624 10606 11652 11630
rect 11750 11452 12046 11472
rect 11806 11450 11830 11452
rect 11886 11450 11910 11452
rect 11966 11450 11990 11452
rect 11828 11398 11830 11450
rect 11892 11398 11904 11450
rect 11966 11398 11968 11450
rect 11806 11396 11830 11398
rect 11886 11396 11910 11398
rect 11966 11396 11990 11398
rect 11750 11376 12046 11396
rect 12268 11150 12296 11698
rect 12452 11218 12480 14554
rect 12544 14482 12572 16000
rect 12636 15434 12664 16390
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12532 14476 12584 14482
rect 12636 14464 12664 15370
rect 12820 15162 12848 15506
rect 12912 15366 12940 15846
rect 13004 15706 13032 15846
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 13004 15570 13032 15642
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12820 14482 12848 15098
rect 13004 14550 13032 15506
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 12716 14476 12768 14482
rect 12636 14436 12716 14464
rect 12532 14418 12584 14424
rect 12716 14418 12768 14424
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12636 13938 12664 14214
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12728 13530 12756 14418
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12820 13376 12848 14418
rect 12900 13796 12952 13802
rect 13004 13784 13032 14486
rect 12952 13756 13032 13784
rect 12900 13738 12952 13744
rect 12900 13388 12952 13394
rect 12820 13348 12900 13376
rect 12900 13330 12952 13336
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12728 11694 12756 13126
rect 12912 12986 12940 13330
rect 13004 13258 13032 13756
rect 12992 13252 13044 13258
rect 12992 13194 13044 13200
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 13004 12442 13032 12718
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 13004 11830 13032 12378
rect 12992 11824 13044 11830
rect 12992 11766 13044 11772
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12728 11354 12756 11630
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12992 11280 13044 11286
rect 12992 11222 13044 11228
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 13004 10810 13032 11222
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 10244 9738 10272 10542
rect 11750 10364 12046 10384
rect 11806 10362 11830 10364
rect 11886 10362 11910 10364
rect 11966 10362 11990 10364
rect 11828 10310 11830 10362
rect 11892 10310 11904 10362
rect 11966 10310 11968 10362
rect 11806 10308 11830 10310
rect 11886 10308 11910 10310
rect 11966 10308 11990 10310
rect 11750 10288 12046 10308
rect 10244 9722 10548 9738
rect 10244 9716 10560 9722
rect 10244 9710 10508 9716
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 9968 7954 9996 9114
rect 10244 8430 10272 9710
rect 10508 9658 10560 9664
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10704 9518 10732 9590
rect 13188 9586 13216 17478
rect 13464 17134 13492 17614
rect 13912 17536 13964 17542
rect 13912 17478 13964 17484
rect 13924 17202 13952 17478
rect 14449 17436 14745 17456
rect 14505 17434 14529 17436
rect 14585 17434 14609 17436
rect 14665 17434 14689 17436
rect 14527 17382 14529 17434
rect 14591 17382 14603 17434
rect 14665 17382 14667 17434
rect 14505 17380 14529 17382
rect 14585 17380 14609 17382
rect 14665 17380 14689 17382
rect 14449 17360 14745 17380
rect 15396 17338 15424 17614
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 15580 17134 15608 19071
rect 15672 17270 15700 19804
rect 17052 17814 17080 19804
rect 16028 17808 16080 17814
rect 16028 17750 16080 17756
rect 17040 17808 17092 17814
rect 17040 17750 17092 17756
rect 16040 17338 16068 17750
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 15660 17264 15712 17270
rect 15660 17206 15712 17212
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13372 15570 13400 16594
rect 13464 16114 13492 17070
rect 14556 17060 14608 17066
rect 14556 17002 14608 17008
rect 14568 16794 14596 17002
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 14449 16348 14745 16368
rect 14505 16346 14529 16348
rect 14585 16346 14609 16348
rect 14665 16346 14689 16348
rect 14527 16294 14529 16346
rect 14591 16294 14603 16346
rect 14665 16294 14667 16346
rect 14505 16292 14529 16294
rect 14585 16292 14609 16294
rect 14665 16292 14689 16294
rect 14449 16272 14745 16292
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13464 15706 13492 15914
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13360 15564 13412 15570
rect 13280 15524 13360 15552
rect 13280 13394 13308 15524
rect 13360 15506 13412 15512
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13832 15026 13860 15302
rect 14449 15260 14745 15280
rect 14505 15258 14529 15260
rect 14585 15258 14609 15260
rect 14665 15258 14689 15260
rect 14527 15206 14529 15258
rect 14591 15206 14603 15258
rect 14665 15206 14667 15258
rect 14505 15204 14529 15206
rect 14585 15204 14609 15206
rect 14665 15204 14689 15206
rect 14449 15184 14745 15204
rect 15304 15162 15332 15506
rect 14372 15156 14424 15162
rect 14372 15098 14424 15104
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 14384 14958 14412 15098
rect 14924 15088 14976 15094
rect 14924 15030 14976 15036
rect 14936 14958 14964 15030
rect 15028 15026 15056 15098
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 15304 14958 15332 15098
rect 14372 14952 14424 14958
rect 14924 14952 14976 14958
rect 14372 14894 14424 14900
rect 14844 14912 14924 14940
rect 14096 14544 14148 14550
rect 14096 14486 14148 14492
rect 13360 14340 13412 14346
rect 13360 14282 13412 14288
rect 13372 14074 13400 14282
rect 14108 14074 14136 14486
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 13360 13796 13412 13802
rect 13360 13738 13412 13744
rect 13372 13530 13400 13738
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13544 13456 13596 13462
rect 13544 13398 13596 13404
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13372 11898 13400 12242
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13464 11762 13492 12038
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13556 11694 13584 13398
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13648 12442 13676 13262
rect 14108 12782 14136 14010
rect 14292 13734 14320 14350
rect 14384 14074 14412 14894
rect 14449 14172 14745 14192
rect 14505 14170 14529 14172
rect 14585 14170 14609 14172
rect 14665 14170 14689 14172
rect 14527 14118 14529 14170
rect 14591 14118 14603 14170
rect 14665 14118 14667 14170
rect 14505 14116 14529 14118
rect 14585 14116 14609 14118
rect 14665 14116 14689 14118
rect 14449 14096 14745 14116
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 14292 12986 14320 13670
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14096 12776 14148 12782
rect 14016 12736 14096 12764
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13740 11694 13768 12038
rect 13924 11694 13952 12106
rect 14016 11762 14044 12736
rect 14096 12718 14148 12724
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 14108 11694 14136 12310
rect 14292 12238 14320 12922
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13372 11354 13400 11562
rect 13556 11354 13584 11630
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13740 11286 13768 11494
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 14016 10538 14044 11086
rect 14108 10674 14136 11494
rect 14384 11082 14412 13874
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14752 13394 14780 13670
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14449 13084 14745 13104
rect 14505 13082 14529 13084
rect 14585 13082 14609 13084
rect 14665 13082 14689 13084
rect 14527 13030 14529 13082
rect 14591 13030 14603 13082
rect 14665 13030 14667 13082
rect 14505 13028 14529 13030
rect 14585 13028 14609 13030
rect 14665 13028 14689 13030
rect 14449 13008 14745 13028
rect 14844 12986 14872 14912
rect 14924 14894 14976 14900
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15120 14822 15148 14894
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 14936 13410 14964 13806
rect 14936 13394 15056 13410
rect 14936 13388 15068 13394
rect 14936 13382 15016 13388
rect 15016 13330 15068 13336
rect 15120 12986 15148 14758
rect 15396 14482 15424 16390
rect 15384 14476 15436 14482
rect 15212 14436 15384 14464
rect 15212 13462 15240 14436
rect 15384 14418 15436 14424
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15304 13938 15332 14214
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15384 13796 15436 13802
rect 15384 13738 15436 13744
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 15396 13326 15424 13738
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15396 12782 15424 13262
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15212 12306 15240 12718
rect 15396 12374 15424 12718
rect 15488 12434 15516 16934
rect 15580 14958 15608 16934
rect 15764 16658 15792 17070
rect 16316 16658 16344 17478
rect 16762 17096 16818 17105
rect 16762 17031 16764 17040
rect 16816 17031 16818 17040
rect 16764 17002 16816 17008
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 16028 16652 16080 16658
rect 16304 16652 16356 16658
rect 16080 16612 16304 16640
rect 16028 16594 16080 16600
rect 16304 16594 16356 16600
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 15764 15570 15792 16594
rect 16040 16114 16068 16594
rect 16776 16250 16804 16594
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 16028 15972 16080 15978
rect 16028 15914 16080 15920
rect 16040 15706 16068 15914
rect 16028 15700 16080 15706
rect 16028 15642 16080 15648
rect 15752 15564 15804 15570
rect 15752 15506 15804 15512
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15568 14544 15620 14550
rect 15568 14486 15620 14492
rect 15580 13920 15608 14486
rect 15660 13932 15712 13938
rect 15580 13892 15660 13920
rect 15580 13394 15608 13892
rect 15660 13874 15712 13880
rect 16304 13796 16356 13802
rect 16304 13738 16356 13744
rect 16316 13530 16344 13738
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16500 13394 16528 15506
rect 16762 15056 16818 15065
rect 16762 14991 16818 15000
rect 16776 14958 16804 14991
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 15488 12406 15608 12434
rect 15384 12368 15436 12374
rect 15384 12310 15436 12316
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 14449 11996 14745 12016
rect 14505 11994 14529 11996
rect 14585 11994 14609 11996
rect 14665 11994 14689 11996
rect 14527 11942 14529 11994
rect 14591 11942 14603 11994
rect 14665 11942 14667 11994
rect 14505 11940 14529 11942
rect 14585 11940 14609 11942
rect 14665 11940 14689 11942
rect 14449 11920 14745 11940
rect 15212 11898 15240 12242
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15488 11762 15516 12242
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14844 11286 14872 11494
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 15384 11280 15436 11286
rect 15488 11268 15516 11698
rect 15436 11240 15516 11268
rect 15384 11222 15436 11228
rect 14372 11076 14424 11082
rect 14372 11018 14424 11024
rect 14449 10908 14745 10928
rect 14505 10906 14529 10908
rect 14585 10906 14609 10908
rect 14665 10906 14689 10908
rect 14527 10854 14529 10906
rect 14591 10854 14603 10906
rect 14665 10854 14667 10906
rect 14505 10852 14529 10854
rect 14585 10852 14609 10854
rect 14665 10852 14689 10854
rect 14449 10832 14745 10852
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14004 10532 14056 10538
rect 14004 10474 14056 10480
rect 14832 10532 14884 10538
rect 14832 10474 14884 10480
rect 14844 10266 14872 10474
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14449 9820 14745 9840
rect 14505 9818 14529 9820
rect 14585 9818 14609 9820
rect 14665 9818 14689 9820
rect 14527 9766 14529 9818
rect 14591 9766 14603 9818
rect 14665 9766 14667 9818
rect 14505 9764 14529 9766
rect 14585 9764 14609 9766
rect 14665 9764 14689 9766
rect 14449 9744 14745 9764
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11256 9382 11284 9454
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9968 7206 9996 7890
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9052 4380 9348 4400
rect 9108 4378 9132 4380
rect 9188 4378 9212 4380
rect 9268 4378 9292 4380
rect 9130 4326 9132 4378
rect 9194 4326 9206 4378
rect 9268 4326 9270 4378
rect 9108 4324 9132 4326
rect 9188 4324 9212 4326
rect 9268 4324 9292 4326
rect 9052 4304 9348 4324
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9052 3292 9348 3312
rect 9108 3290 9132 3292
rect 9188 3290 9212 3292
rect 9268 3290 9292 3292
rect 9130 3238 9132 3290
rect 9194 3238 9206 3290
rect 9268 3238 9270 3290
rect 9108 3236 9132 3238
rect 9188 3236 9212 3238
rect 9268 3236 9292 3238
rect 9052 3216 9348 3236
rect 9416 3194 9444 3470
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 9600 2990 9628 6598
rect 10232 5772 10284 5778
rect 10232 5714 10284 5720
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10152 4690 10180 5510
rect 10244 5234 10272 5714
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10244 5030 10272 5170
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9692 2650 9720 2858
rect 10152 2854 10180 3334
rect 10336 3194 10364 3674
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 10336 2774 10364 3130
rect 10520 2854 10548 8298
rect 10612 7546 10640 8978
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10980 8566 11008 8910
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 11256 8498 11284 9318
rect 11624 9178 11652 9318
rect 11750 9276 12046 9296
rect 11806 9274 11830 9276
rect 11886 9274 11910 9276
rect 11966 9274 11990 9276
rect 11828 9222 11830 9274
rect 11892 9222 11904 9274
rect 11966 9222 11968 9274
rect 11806 9220 11830 9222
rect 11886 9220 11910 9222
rect 11966 9220 11990 9222
rect 11750 9200 12046 9220
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 12176 9110 12204 9318
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12452 9042 12480 9522
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 11428 8968 11480 8974
rect 11348 8928 11428 8956
rect 11348 8838 11376 8928
rect 11428 8910 11480 8916
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10612 7410 10640 7482
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10704 5250 10732 8230
rect 11750 8188 12046 8208
rect 11806 8186 11830 8188
rect 11886 8186 11910 8188
rect 11966 8186 11990 8188
rect 11828 8134 11830 8186
rect 11892 8134 11904 8186
rect 11966 8134 11968 8186
rect 11806 8132 11830 8134
rect 11886 8132 11910 8134
rect 11966 8132 11990 8134
rect 11750 8112 12046 8132
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 11336 7472 11388 7478
rect 11336 7414 11388 7420
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10796 6254 10824 6938
rect 10980 6934 11008 7210
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 10876 6724 10928 6730
rect 10876 6666 10928 6672
rect 10888 6458 10916 6666
rect 11072 6458 11100 7278
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 11164 6186 11192 6802
rect 11348 6322 11376 7414
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 11750 7100 12046 7120
rect 11806 7098 11830 7100
rect 11886 7098 11910 7100
rect 11966 7098 11990 7100
rect 11828 7046 11830 7098
rect 11892 7046 11904 7098
rect 11966 7046 11968 7098
rect 11806 7044 11830 7046
rect 11886 7044 11910 7046
rect 11966 7044 11990 7046
rect 11750 7024 12046 7044
rect 12084 6866 12112 7278
rect 12544 6934 12572 8026
rect 12636 7342 12664 8978
rect 12820 8974 12848 9522
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 13004 9178 13032 9318
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13096 8498 13124 8910
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12820 7002 12848 7142
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 13096 6798 13124 8434
rect 13280 8430 13308 8978
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 11152 6180 11204 6186
rect 11152 6122 11204 6128
rect 11750 6012 12046 6032
rect 11806 6010 11830 6012
rect 11886 6010 11910 6012
rect 11966 6010 11990 6012
rect 11828 5958 11830 6010
rect 11892 5958 11904 6010
rect 11966 5958 11968 6010
rect 11806 5956 11830 5958
rect 11886 5956 11910 5958
rect 11966 5956 11990 5958
rect 11750 5936 12046 5956
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 10612 5222 10824 5250
rect 10612 5166 10640 5222
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10692 5160 10744 5166
rect 10796 5148 10824 5222
rect 11716 5166 11744 5646
rect 12084 5234 12112 5850
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12452 5370 12480 5714
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 10744 5120 10824 5148
rect 11704 5160 11756 5166
rect 10692 5102 10744 5108
rect 11704 5102 11756 5108
rect 12084 5030 12112 5170
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 11750 4924 12046 4944
rect 11806 4922 11830 4924
rect 11886 4922 11910 4924
rect 11966 4922 11990 4924
rect 11828 4870 11830 4922
rect 11892 4870 11904 4922
rect 11966 4870 11968 4922
rect 11806 4868 11830 4870
rect 11886 4868 11910 4870
rect 11966 4868 11990 4870
rect 11750 4848 12046 4868
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 11072 3738 11100 4626
rect 12452 4554 12480 5034
rect 12544 4622 12572 6734
rect 13280 6730 13308 7346
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13372 5234 13400 9318
rect 15488 9042 15516 9318
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 13912 8900 13964 8906
rect 13912 8842 13964 8848
rect 13924 8430 13952 8842
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 14016 7342 14044 8978
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 14108 7478 14136 8298
rect 14096 7472 14148 7478
rect 14096 7414 14148 7420
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13556 6254 13584 7142
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 14384 4826 14412 8774
rect 14449 8732 14745 8752
rect 14505 8730 14529 8732
rect 14585 8730 14609 8732
rect 14665 8730 14689 8732
rect 14527 8678 14529 8730
rect 14591 8678 14603 8730
rect 14665 8678 14667 8730
rect 14505 8676 14529 8678
rect 14585 8676 14609 8678
rect 14665 8676 14689 8678
rect 14449 8656 14745 8676
rect 14936 7818 14964 8978
rect 15580 8566 15608 12406
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15672 11626 15700 12242
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 15660 11620 15712 11626
rect 15660 11562 15712 11568
rect 16040 10674 16068 11630
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 16224 10606 16252 13330
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 16408 10985 16436 11630
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16394 10976 16450 10985
rect 16394 10911 16450 10920
rect 16500 10810 16528 11222
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16224 10130 16252 10542
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16684 9586 16712 14758
rect 16762 13016 16818 13025
rect 16762 12951 16818 12960
rect 16776 12782 16804 12951
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 15568 8560 15620 8566
rect 15568 8502 15620 8508
rect 15856 7954 15884 8978
rect 16132 8430 16160 9114
rect 16592 8498 16620 9318
rect 16776 8945 16804 9454
rect 16762 8936 16818 8945
rect 16762 8871 16818 8880
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 15948 7954 15976 8298
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 14924 7812 14976 7818
rect 14924 7754 14976 7760
rect 14449 7644 14745 7664
rect 14505 7642 14529 7644
rect 14585 7642 14609 7644
rect 14665 7642 14689 7644
rect 14527 7590 14529 7642
rect 14591 7590 14603 7642
rect 14665 7590 14667 7642
rect 14505 7588 14529 7590
rect 14585 7588 14609 7590
rect 14665 7588 14689 7590
rect 14449 7568 14745 7588
rect 14936 7342 14964 7754
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 15856 7002 15884 7890
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 14449 6556 14745 6576
rect 14505 6554 14529 6556
rect 14585 6554 14609 6556
rect 14665 6554 14689 6556
rect 14527 6502 14529 6554
rect 14591 6502 14603 6554
rect 14665 6502 14667 6554
rect 14505 6500 14529 6502
rect 14585 6500 14609 6502
rect 14665 6500 14689 6502
rect 14449 6480 14745 6500
rect 15856 6458 15884 6802
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 14449 5468 14745 5488
rect 14505 5466 14529 5468
rect 14585 5466 14609 5468
rect 14665 5466 14689 5468
rect 14527 5414 14529 5466
rect 14591 5414 14603 5466
rect 14665 5414 14667 5466
rect 14505 5412 14529 5414
rect 14585 5412 14609 5414
rect 14665 5412 14689 5414
rect 14449 5392 14745 5412
rect 15304 5234 15332 6190
rect 15856 5914 15884 6190
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15396 4826 15424 5102
rect 15856 5030 15884 5714
rect 15844 5024 15896 5030
rect 15844 4966 15896 4972
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10612 2990 10640 3538
rect 10980 3194 11008 3538
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10336 2746 10456 2774
rect 10428 2650 10456 2746
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 9052 2204 9348 2224
rect 9108 2202 9132 2204
rect 9188 2202 9212 2204
rect 9268 2202 9292 2204
rect 9130 2150 9132 2202
rect 9194 2150 9206 2202
rect 9268 2150 9270 2202
rect 9108 2148 9132 2150
rect 9188 2148 9212 2150
rect 9268 2148 9292 2150
rect 9052 2128 9348 2148
rect 9692 800 9720 2450
rect 10980 2378 11008 2858
rect 11072 2650 11100 3470
rect 11348 2990 11376 3878
rect 11750 3836 12046 3856
rect 11806 3834 11830 3836
rect 11886 3834 11910 3836
rect 11966 3834 11990 3836
rect 11828 3782 11830 3834
rect 11892 3782 11904 3834
rect 11966 3782 11968 3834
rect 11806 3780 11830 3782
rect 11886 3780 11910 3782
rect 11966 3780 11990 3782
rect 11750 3760 12046 3780
rect 12452 3194 12480 3878
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12544 3058 12572 4558
rect 14449 4380 14745 4400
rect 14505 4378 14529 4380
rect 14585 4378 14609 4380
rect 14665 4378 14689 4380
rect 14527 4326 14529 4378
rect 14591 4326 14603 4378
rect 14665 4326 14667 4378
rect 14505 4324 14529 4326
rect 14585 4324 14609 4326
rect 14665 4324 14689 4326
rect 14449 4304 14745 4324
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 12728 3670 12756 4082
rect 13268 4004 13320 4010
rect 13268 3946 13320 3952
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11750 2748 12046 2768
rect 11806 2746 11830 2748
rect 11886 2746 11910 2748
rect 11966 2746 11990 2748
rect 11828 2694 11830 2746
rect 11892 2694 11904 2746
rect 11966 2694 11968 2746
rect 11806 2692 11830 2694
rect 11886 2692 11910 2694
rect 11966 2692 11990 2694
rect 11750 2672 12046 2692
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 11072 800 11100 2450
rect 12452 800 12480 2450
rect 12544 2428 12572 2994
rect 13004 2582 13032 3470
rect 13188 3058 13216 3878
rect 13280 3602 13308 3946
rect 13648 3738 13676 4082
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13832 3670 13860 4014
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 13728 3460 13780 3466
rect 13728 3402 13780 3408
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 13648 2650 13676 2994
rect 13740 2990 13768 3402
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 12992 2576 13044 2582
rect 12992 2518 13044 2524
rect 13832 2514 13860 3606
rect 14200 3194 14228 4014
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14200 2650 14228 3130
rect 14292 2990 14320 3946
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14384 3058 14412 3878
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 14449 3292 14745 3312
rect 14505 3290 14529 3292
rect 14585 3290 14609 3292
rect 14665 3290 14689 3292
rect 14527 3238 14529 3290
rect 14591 3238 14603 3290
rect 14665 3238 14667 3290
rect 14505 3236 14529 3238
rect 14585 3236 14609 3238
rect 14665 3236 14689 3238
rect 14449 3216 14745 3236
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 15028 2990 15056 3470
rect 15396 3194 15424 4558
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 15488 3398 15516 3606
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14936 2650 14964 2790
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 12624 2440 12676 2446
rect 12544 2400 12624 2428
rect 12624 2382 12676 2388
rect 13924 1306 13952 2450
rect 14449 2204 14745 2224
rect 14505 2202 14529 2204
rect 14585 2202 14609 2204
rect 14665 2202 14689 2204
rect 14527 2150 14529 2202
rect 14591 2150 14603 2202
rect 14665 2150 14667 2202
rect 14505 2148 14529 2150
rect 14585 2148 14609 2150
rect 14665 2148 14689 2150
rect 14449 2128 14745 2148
rect 13832 1278 13952 1306
rect 13832 800 13860 1278
rect 15212 800 15240 2926
rect 15488 2530 15516 3334
rect 16592 3194 16620 6598
rect 16868 4010 16896 17478
rect 17040 17128 17092 17134
rect 17040 17070 17092 17076
rect 16946 6896 17002 6905
rect 16946 6831 16948 6840
rect 17000 6831 17002 6840
rect 16948 6802 17000 6808
rect 16946 4856 17002 4865
rect 16946 4791 17002 4800
rect 16960 4690 16988 4791
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 16856 4004 16908 4010
rect 16856 3946 16908 3952
rect 17052 3602 17080 17070
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16488 2984 16540 2990
rect 16488 2926 16540 2932
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16500 2825 16528 2926
rect 16486 2816 16542 2825
rect 16486 2751 16542 2760
rect 15488 2514 15608 2530
rect 15488 2508 15620 2514
rect 15488 2502 15568 2508
rect 15568 2450 15620 2456
rect 16580 2440 16632 2446
rect 16580 2382 16632 2388
rect 16592 800 16620 2382
rect 478 0 534 800
rect 1398 0 1454 800
rect 2778 0 2834 800
rect 4158 0 4214 800
rect 5538 0 5594 800
rect 6918 0 6974 800
rect 8298 0 8354 800
rect 9678 0 9734 800
rect 11058 0 11114 800
rect 12438 0 12494 800
rect 13818 0 13874 800
rect 15198 0 15254 800
rect 16578 0 16634 800
rect 16776 785 16804 2926
rect 17052 2514 17080 3538
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 16762 776 16818 785
rect 16762 711 16818 720
<< via2 >>
rect 1490 18400 1546 18456
rect 6353 17978 6409 17980
rect 6433 17978 6489 17980
rect 6513 17978 6569 17980
rect 6593 17978 6649 17980
rect 6353 17926 6379 17978
rect 6379 17926 6409 17978
rect 6433 17926 6443 17978
rect 6443 17926 6489 17978
rect 6513 17926 6559 17978
rect 6559 17926 6569 17978
rect 6593 17926 6623 17978
rect 6623 17926 6649 17978
rect 6353 17924 6409 17926
rect 6433 17924 6489 17926
rect 6513 17924 6569 17926
rect 6593 17924 6649 17926
rect 11750 17978 11806 17980
rect 11830 17978 11886 17980
rect 11910 17978 11966 17980
rect 11990 17978 12046 17980
rect 11750 17926 11776 17978
rect 11776 17926 11806 17978
rect 11830 17926 11840 17978
rect 11840 17926 11886 17978
rect 11910 17926 11956 17978
rect 11956 17926 11966 17978
rect 11990 17926 12020 17978
rect 12020 17926 12046 17978
rect 11750 17924 11806 17926
rect 11830 17924 11886 17926
rect 11910 17924 11966 17926
rect 11990 17924 12046 17926
rect 15566 19080 15622 19136
rect 1398 16360 1454 16416
rect 1398 14320 1454 14376
rect 1398 12300 1454 12336
rect 1398 12280 1400 12300
rect 1400 12280 1452 12300
rect 1452 12280 1454 12300
rect 1490 10260 1546 10296
rect 1490 10240 1492 10260
rect 1492 10240 1544 10260
rect 1544 10240 1546 10260
rect 1398 8200 1454 8256
rect 2870 15000 2926 15056
rect 3146 14864 3202 14920
rect 1398 6160 1454 6216
rect 1398 4140 1454 4176
rect 1398 4120 1400 4140
rect 1400 4120 1452 4140
rect 1452 4120 1454 4140
rect 3654 17434 3710 17436
rect 3734 17434 3790 17436
rect 3814 17434 3870 17436
rect 3894 17434 3950 17436
rect 3654 17382 3680 17434
rect 3680 17382 3710 17434
rect 3734 17382 3744 17434
rect 3744 17382 3790 17434
rect 3814 17382 3860 17434
rect 3860 17382 3870 17434
rect 3894 17382 3924 17434
rect 3924 17382 3950 17434
rect 3654 17380 3710 17382
rect 3734 17380 3790 17382
rect 3814 17380 3870 17382
rect 3894 17380 3950 17382
rect 3654 16346 3710 16348
rect 3734 16346 3790 16348
rect 3814 16346 3870 16348
rect 3894 16346 3950 16348
rect 3654 16294 3680 16346
rect 3680 16294 3710 16346
rect 3734 16294 3744 16346
rect 3744 16294 3790 16346
rect 3814 16294 3860 16346
rect 3860 16294 3870 16346
rect 3894 16294 3924 16346
rect 3924 16294 3950 16346
rect 3654 16292 3710 16294
rect 3734 16292 3790 16294
rect 3814 16292 3870 16294
rect 3894 16292 3950 16294
rect 3654 15258 3710 15260
rect 3734 15258 3790 15260
rect 3814 15258 3870 15260
rect 3894 15258 3950 15260
rect 3654 15206 3680 15258
rect 3680 15206 3710 15258
rect 3734 15206 3744 15258
rect 3744 15206 3790 15258
rect 3814 15206 3860 15258
rect 3860 15206 3870 15258
rect 3894 15206 3924 15258
rect 3924 15206 3950 15258
rect 3654 15204 3710 15206
rect 3734 15204 3790 15206
rect 3814 15204 3870 15206
rect 3894 15204 3950 15206
rect 3882 15000 3938 15056
rect 3698 14900 3700 14920
rect 3700 14900 3752 14920
rect 3752 14900 3754 14920
rect 3698 14864 3754 14900
rect 3654 14170 3710 14172
rect 3734 14170 3790 14172
rect 3814 14170 3870 14172
rect 3894 14170 3950 14172
rect 3654 14118 3680 14170
rect 3680 14118 3710 14170
rect 3734 14118 3744 14170
rect 3744 14118 3790 14170
rect 3814 14118 3860 14170
rect 3860 14118 3870 14170
rect 3894 14118 3924 14170
rect 3924 14118 3950 14170
rect 3654 14116 3710 14118
rect 3734 14116 3790 14118
rect 3814 14116 3870 14118
rect 3894 14116 3950 14118
rect 4066 13232 4122 13288
rect 3654 13082 3710 13084
rect 3734 13082 3790 13084
rect 3814 13082 3870 13084
rect 3894 13082 3950 13084
rect 3654 13030 3680 13082
rect 3680 13030 3710 13082
rect 3734 13030 3744 13082
rect 3744 13030 3790 13082
rect 3814 13030 3860 13082
rect 3860 13030 3870 13082
rect 3894 13030 3924 13082
rect 3924 13030 3950 13082
rect 3654 13028 3710 13030
rect 3734 13028 3790 13030
rect 3814 13028 3870 13030
rect 3894 13028 3950 13030
rect 3882 12824 3938 12880
rect 3654 11994 3710 11996
rect 3734 11994 3790 11996
rect 3814 11994 3870 11996
rect 3894 11994 3950 11996
rect 3654 11942 3680 11994
rect 3680 11942 3710 11994
rect 3734 11942 3744 11994
rect 3744 11942 3790 11994
rect 3814 11942 3860 11994
rect 3860 11942 3870 11994
rect 3894 11942 3924 11994
rect 3924 11942 3950 11994
rect 3654 11940 3710 11942
rect 3734 11940 3790 11942
rect 3814 11940 3870 11942
rect 3894 11940 3950 11942
rect 3654 10906 3710 10908
rect 3734 10906 3790 10908
rect 3814 10906 3870 10908
rect 3894 10906 3950 10908
rect 3654 10854 3680 10906
rect 3680 10854 3710 10906
rect 3734 10854 3744 10906
rect 3744 10854 3790 10906
rect 3814 10854 3860 10906
rect 3860 10854 3870 10906
rect 3894 10854 3924 10906
rect 3924 10854 3950 10906
rect 3654 10852 3710 10854
rect 3734 10852 3790 10854
rect 3814 10852 3870 10854
rect 3894 10852 3950 10854
rect 3654 9818 3710 9820
rect 3734 9818 3790 9820
rect 3814 9818 3870 9820
rect 3894 9818 3950 9820
rect 3654 9766 3680 9818
rect 3680 9766 3710 9818
rect 3734 9766 3744 9818
rect 3744 9766 3790 9818
rect 3814 9766 3860 9818
rect 3860 9766 3870 9818
rect 3894 9766 3924 9818
rect 3924 9766 3950 9818
rect 3654 9764 3710 9766
rect 3734 9764 3790 9766
rect 3814 9764 3870 9766
rect 3894 9764 3950 9766
rect 3654 8730 3710 8732
rect 3734 8730 3790 8732
rect 3814 8730 3870 8732
rect 3894 8730 3950 8732
rect 3654 8678 3680 8730
rect 3680 8678 3710 8730
rect 3734 8678 3744 8730
rect 3744 8678 3790 8730
rect 3814 8678 3860 8730
rect 3860 8678 3870 8730
rect 3894 8678 3924 8730
rect 3924 8678 3950 8730
rect 3654 8676 3710 8678
rect 3734 8676 3790 8678
rect 3814 8676 3870 8678
rect 3894 8676 3950 8678
rect 3654 7642 3710 7644
rect 3734 7642 3790 7644
rect 3814 7642 3870 7644
rect 3894 7642 3950 7644
rect 3654 7590 3680 7642
rect 3680 7590 3710 7642
rect 3734 7590 3744 7642
rect 3744 7590 3790 7642
rect 3814 7590 3860 7642
rect 3860 7590 3870 7642
rect 3894 7590 3924 7642
rect 3924 7590 3950 7642
rect 3654 7588 3710 7590
rect 3734 7588 3790 7590
rect 3814 7588 3870 7590
rect 3894 7588 3950 7590
rect 3654 6554 3710 6556
rect 3734 6554 3790 6556
rect 3814 6554 3870 6556
rect 3894 6554 3950 6556
rect 3654 6502 3680 6554
rect 3680 6502 3710 6554
rect 3734 6502 3744 6554
rect 3744 6502 3790 6554
rect 3814 6502 3860 6554
rect 3860 6502 3870 6554
rect 3894 6502 3924 6554
rect 3924 6502 3950 6554
rect 3654 6500 3710 6502
rect 3734 6500 3790 6502
rect 3814 6500 3870 6502
rect 3894 6500 3950 6502
rect 4710 15000 4766 15056
rect 3654 5466 3710 5468
rect 3734 5466 3790 5468
rect 3814 5466 3870 5468
rect 3894 5466 3950 5468
rect 3654 5414 3680 5466
rect 3680 5414 3710 5466
rect 3734 5414 3744 5466
rect 3744 5414 3790 5466
rect 3814 5414 3860 5466
rect 3860 5414 3870 5466
rect 3894 5414 3924 5466
rect 3924 5414 3950 5466
rect 3654 5412 3710 5414
rect 3734 5412 3790 5414
rect 3814 5412 3870 5414
rect 3894 5412 3950 5414
rect 3654 4378 3710 4380
rect 3734 4378 3790 4380
rect 3814 4378 3870 4380
rect 3894 4378 3950 4380
rect 3654 4326 3680 4378
rect 3680 4326 3710 4378
rect 3734 4326 3744 4378
rect 3744 4326 3790 4378
rect 3814 4326 3860 4378
rect 3860 4326 3870 4378
rect 3894 4326 3924 4378
rect 3924 4326 3950 4378
rect 3654 4324 3710 4326
rect 3734 4324 3790 4326
rect 3814 4324 3870 4326
rect 3894 4324 3950 4326
rect 6353 16890 6409 16892
rect 6433 16890 6489 16892
rect 6513 16890 6569 16892
rect 6593 16890 6649 16892
rect 6353 16838 6379 16890
rect 6379 16838 6409 16890
rect 6433 16838 6443 16890
rect 6443 16838 6489 16890
rect 6513 16838 6559 16890
rect 6559 16838 6569 16890
rect 6593 16838 6623 16890
rect 6623 16838 6649 16890
rect 6353 16836 6409 16838
rect 6433 16836 6489 16838
rect 6513 16836 6569 16838
rect 6593 16836 6649 16838
rect 6353 15802 6409 15804
rect 6433 15802 6489 15804
rect 6513 15802 6569 15804
rect 6593 15802 6649 15804
rect 6353 15750 6379 15802
rect 6379 15750 6409 15802
rect 6433 15750 6443 15802
rect 6443 15750 6489 15802
rect 6513 15750 6559 15802
rect 6559 15750 6569 15802
rect 6593 15750 6623 15802
rect 6623 15750 6649 15802
rect 6353 15748 6409 15750
rect 6433 15748 6489 15750
rect 6513 15748 6569 15750
rect 6593 15748 6649 15750
rect 6353 14714 6409 14716
rect 6433 14714 6489 14716
rect 6513 14714 6569 14716
rect 6593 14714 6649 14716
rect 6353 14662 6379 14714
rect 6379 14662 6409 14714
rect 6433 14662 6443 14714
rect 6443 14662 6489 14714
rect 6513 14662 6559 14714
rect 6559 14662 6569 14714
rect 6593 14662 6623 14714
rect 6623 14662 6649 14714
rect 6353 14660 6409 14662
rect 6433 14660 6489 14662
rect 6513 14660 6569 14662
rect 6593 14660 6649 14662
rect 6353 13626 6409 13628
rect 6433 13626 6489 13628
rect 6513 13626 6569 13628
rect 6593 13626 6649 13628
rect 6353 13574 6379 13626
rect 6379 13574 6409 13626
rect 6433 13574 6443 13626
rect 6443 13574 6489 13626
rect 6513 13574 6559 13626
rect 6559 13574 6569 13626
rect 6593 13574 6623 13626
rect 6623 13574 6649 13626
rect 6353 13572 6409 13574
rect 6433 13572 6489 13574
rect 6513 13572 6569 13574
rect 6593 13572 6649 13574
rect 5906 12824 5962 12880
rect 6353 12538 6409 12540
rect 6433 12538 6489 12540
rect 6513 12538 6569 12540
rect 6593 12538 6649 12540
rect 6353 12486 6379 12538
rect 6379 12486 6409 12538
rect 6433 12486 6443 12538
rect 6443 12486 6489 12538
rect 6513 12486 6559 12538
rect 6559 12486 6569 12538
rect 6593 12486 6623 12538
rect 6623 12486 6649 12538
rect 6353 12484 6409 12486
rect 6433 12484 6489 12486
rect 6513 12484 6569 12486
rect 6593 12484 6649 12486
rect 6353 11450 6409 11452
rect 6433 11450 6489 11452
rect 6513 11450 6569 11452
rect 6593 11450 6649 11452
rect 6353 11398 6379 11450
rect 6379 11398 6409 11450
rect 6433 11398 6443 11450
rect 6443 11398 6489 11450
rect 6513 11398 6559 11450
rect 6559 11398 6569 11450
rect 6593 11398 6623 11450
rect 6623 11398 6649 11450
rect 6353 11396 6409 11398
rect 6433 11396 6489 11398
rect 6513 11396 6569 11398
rect 6593 11396 6649 11398
rect 6353 10362 6409 10364
rect 6433 10362 6489 10364
rect 6513 10362 6569 10364
rect 6593 10362 6649 10364
rect 6353 10310 6379 10362
rect 6379 10310 6409 10362
rect 6433 10310 6443 10362
rect 6443 10310 6489 10362
rect 6513 10310 6559 10362
rect 6559 10310 6569 10362
rect 6593 10310 6623 10362
rect 6623 10310 6649 10362
rect 6353 10308 6409 10310
rect 6433 10308 6489 10310
rect 6513 10308 6569 10310
rect 6593 10308 6649 10310
rect 5998 8372 6000 8392
rect 6000 8372 6052 8392
rect 6052 8372 6054 8392
rect 3654 3290 3710 3292
rect 3734 3290 3790 3292
rect 3814 3290 3870 3292
rect 3894 3290 3950 3292
rect 3654 3238 3680 3290
rect 3680 3238 3710 3290
rect 3734 3238 3744 3290
rect 3744 3238 3790 3290
rect 3814 3238 3860 3290
rect 3860 3238 3870 3290
rect 3894 3238 3924 3290
rect 3924 3238 3950 3290
rect 3654 3236 3710 3238
rect 3734 3236 3790 3238
rect 3814 3236 3870 3238
rect 3894 3236 3950 3238
rect 2042 2080 2098 2136
rect 3654 2202 3710 2204
rect 3734 2202 3790 2204
rect 3814 2202 3870 2204
rect 3894 2202 3950 2204
rect 3654 2150 3680 2202
rect 3680 2150 3710 2202
rect 3734 2150 3744 2202
rect 3744 2150 3790 2202
rect 3814 2150 3860 2202
rect 3860 2150 3870 2202
rect 3894 2150 3924 2202
rect 3924 2150 3950 2202
rect 3654 2148 3710 2150
rect 3734 2148 3790 2150
rect 3814 2148 3870 2150
rect 3894 2148 3950 2150
rect 5998 8336 6054 8372
rect 6353 9274 6409 9276
rect 6433 9274 6489 9276
rect 6513 9274 6569 9276
rect 6593 9274 6649 9276
rect 6353 9222 6379 9274
rect 6379 9222 6409 9274
rect 6433 9222 6443 9274
rect 6443 9222 6489 9274
rect 6513 9222 6559 9274
rect 6559 9222 6569 9274
rect 6593 9222 6623 9274
rect 6623 9222 6649 9274
rect 6353 9220 6409 9222
rect 6433 9220 6489 9222
rect 6513 9220 6569 9222
rect 6593 9220 6649 9222
rect 6353 8186 6409 8188
rect 6433 8186 6489 8188
rect 6513 8186 6569 8188
rect 6593 8186 6649 8188
rect 6353 8134 6379 8186
rect 6379 8134 6409 8186
rect 6433 8134 6443 8186
rect 6443 8134 6489 8186
rect 6513 8134 6559 8186
rect 6559 8134 6569 8186
rect 6593 8134 6623 8186
rect 6623 8134 6649 8186
rect 6353 8132 6409 8134
rect 6433 8132 6489 8134
rect 6513 8132 6569 8134
rect 6593 8132 6649 8134
rect 6353 7098 6409 7100
rect 6433 7098 6489 7100
rect 6513 7098 6569 7100
rect 6593 7098 6649 7100
rect 6353 7046 6379 7098
rect 6379 7046 6409 7098
rect 6433 7046 6443 7098
rect 6443 7046 6489 7098
rect 6513 7046 6559 7098
rect 6559 7046 6569 7098
rect 6593 7046 6623 7098
rect 6623 7046 6649 7098
rect 6353 7044 6409 7046
rect 6433 7044 6489 7046
rect 6513 7044 6569 7046
rect 6593 7044 6649 7046
rect 7194 12824 7250 12880
rect 9052 17434 9108 17436
rect 9132 17434 9188 17436
rect 9212 17434 9268 17436
rect 9292 17434 9348 17436
rect 9052 17382 9078 17434
rect 9078 17382 9108 17434
rect 9132 17382 9142 17434
rect 9142 17382 9188 17434
rect 9212 17382 9258 17434
rect 9258 17382 9268 17434
rect 9292 17382 9322 17434
rect 9322 17382 9348 17434
rect 9052 17380 9108 17382
rect 9132 17380 9188 17382
rect 9212 17380 9268 17382
rect 9292 17380 9348 17382
rect 9052 16346 9108 16348
rect 9132 16346 9188 16348
rect 9212 16346 9268 16348
rect 9292 16346 9348 16348
rect 9052 16294 9078 16346
rect 9078 16294 9108 16346
rect 9132 16294 9142 16346
rect 9142 16294 9188 16346
rect 9212 16294 9258 16346
rect 9258 16294 9268 16346
rect 9292 16294 9322 16346
rect 9322 16294 9348 16346
rect 9052 16292 9108 16294
rect 9132 16292 9188 16294
rect 9212 16292 9268 16294
rect 9292 16292 9348 16294
rect 9052 15258 9108 15260
rect 9132 15258 9188 15260
rect 9212 15258 9268 15260
rect 9292 15258 9348 15260
rect 9052 15206 9078 15258
rect 9078 15206 9108 15258
rect 9132 15206 9142 15258
rect 9142 15206 9188 15258
rect 9212 15206 9258 15258
rect 9258 15206 9268 15258
rect 9292 15206 9322 15258
rect 9322 15206 9348 15258
rect 9052 15204 9108 15206
rect 9132 15204 9188 15206
rect 9212 15204 9268 15206
rect 9292 15204 9348 15206
rect 9052 14170 9108 14172
rect 9132 14170 9188 14172
rect 9212 14170 9268 14172
rect 9292 14170 9348 14172
rect 9052 14118 9078 14170
rect 9078 14118 9108 14170
rect 9132 14118 9142 14170
rect 9142 14118 9188 14170
rect 9212 14118 9258 14170
rect 9258 14118 9268 14170
rect 9292 14118 9322 14170
rect 9322 14118 9348 14170
rect 9052 14116 9108 14118
rect 9132 14116 9188 14118
rect 9212 14116 9268 14118
rect 9292 14116 9348 14118
rect 9052 13082 9108 13084
rect 9132 13082 9188 13084
rect 9212 13082 9268 13084
rect 9292 13082 9348 13084
rect 9052 13030 9078 13082
rect 9078 13030 9108 13082
rect 9132 13030 9142 13082
rect 9142 13030 9188 13082
rect 9212 13030 9258 13082
rect 9258 13030 9268 13082
rect 9292 13030 9322 13082
rect 9322 13030 9348 13082
rect 9052 13028 9108 13030
rect 9132 13028 9188 13030
rect 9212 13028 9268 13030
rect 9292 13028 9348 13030
rect 9052 11994 9108 11996
rect 9132 11994 9188 11996
rect 9212 11994 9268 11996
rect 9292 11994 9348 11996
rect 9052 11942 9078 11994
rect 9078 11942 9108 11994
rect 9132 11942 9142 11994
rect 9142 11942 9188 11994
rect 9212 11942 9258 11994
rect 9258 11942 9268 11994
rect 9292 11942 9322 11994
rect 9322 11942 9348 11994
rect 9052 11940 9108 11942
rect 9132 11940 9188 11942
rect 9212 11940 9268 11942
rect 9292 11940 9348 11942
rect 9052 10906 9108 10908
rect 9132 10906 9188 10908
rect 9212 10906 9268 10908
rect 9292 10906 9348 10908
rect 9052 10854 9078 10906
rect 9078 10854 9108 10906
rect 9132 10854 9142 10906
rect 9142 10854 9188 10906
rect 9212 10854 9258 10906
rect 9258 10854 9268 10906
rect 9292 10854 9322 10906
rect 9322 10854 9348 10906
rect 9052 10852 9108 10854
rect 9132 10852 9188 10854
rect 9212 10852 9268 10854
rect 9292 10852 9348 10854
rect 7562 9460 7564 9480
rect 7564 9460 7616 9480
rect 7616 9460 7618 9480
rect 7562 9424 7618 9460
rect 7746 9424 7802 9480
rect 8298 9424 8354 9480
rect 7654 8372 7656 8392
rect 7656 8372 7708 8392
rect 7708 8372 7710 8392
rect 7654 8336 7710 8372
rect 6353 6010 6409 6012
rect 6433 6010 6489 6012
rect 6513 6010 6569 6012
rect 6593 6010 6649 6012
rect 6353 5958 6379 6010
rect 6379 5958 6409 6010
rect 6433 5958 6443 6010
rect 6443 5958 6489 6010
rect 6513 5958 6559 6010
rect 6559 5958 6569 6010
rect 6593 5958 6623 6010
rect 6623 5958 6649 6010
rect 6353 5956 6409 5958
rect 6433 5956 6489 5958
rect 6513 5956 6569 5958
rect 6593 5956 6649 5958
rect 6353 4922 6409 4924
rect 6433 4922 6489 4924
rect 6513 4922 6569 4924
rect 6593 4922 6649 4924
rect 6353 4870 6379 4922
rect 6379 4870 6409 4922
rect 6433 4870 6443 4922
rect 6443 4870 6489 4922
rect 6513 4870 6559 4922
rect 6559 4870 6569 4922
rect 6593 4870 6623 4922
rect 6623 4870 6649 4922
rect 6353 4868 6409 4870
rect 6433 4868 6489 4870
rect 6513 4868 6569 4870
rect 6593 4868 6649 4870
rect 9052 9818 9108 9820
rect 9132 9818 9188 9820
rect 9212 9818 9268 9820
rect 9292 9818 9348 9820
rect 9052 9766 9078 9818
rect 9078 9766 9108 9818
rect 9132 9766 9142 9818
rect 9142 9766 9188 9818
rect 9212 9766 9258 9818
rect 9258 9766 9268 9818
rect 9292 9766 9322 9818
rect 9322 9766 9348 9818
rect 9052 9764 9108 9766
rect 9132 9764 9188 9766
rect 9212 9764 9268 9766
rect 9292 9764 9348 9766
rect 9052 8730 9108 8732
rect 9132 8730 9188 8732
rect 9212 8730 9268 8732
rect 9292 8730 9348 8732
rect 9052 8678 9078 8730
rect 9078 8678 9108 8730
rect 9132 8678 9142 8730
rect 9142 8678 9188 8730
rect 9212 8678 9258 8730
rect 9258 8678 9268 8730
rect 9292 8678 9322 8730
rect 9322 8678 9348 8730
rect 9052 8676 9108 8678
rect 9132 8676 9188 8678
rect 9212 8676 9268 8678
rect 9292 8676 9348 8678
rect 9052 7642 9108 7644
rect 9132 7642 9188 7644
rect 9212 7642 9268 7644
rect 9292 7642 9348 7644
rect 9052 7590 9078 7642
rect 9078 7590 9108 7642
rect 9132 7590 9142 7642
rect 9142 7590 9188 7642
rect 9212 7590 9258 7642
rect 9258 7590 9268 7642
rect 9292 7590 9322 7642
rect 9322 7590 9348 7642
rect 9052 7588 9108 7590
rect 9132 7588 9188 7590
rect 9212 7588 9268 7590
rect 9292 7588 9348 7590
rect 6353 3834 6409 3836
rect 6433 3834 6489 3836
rect 6513 3834 6569 3836
rect 6593 3834 6649 3836
rect 6353 3782 6379 3834
rect 6379 3782 6409 3834
rect 6433 3782 6443 3834
rect 6443 3782 6489 3834
rect 6513 3782 6559 3834
rect 6559 3782 6569 3834
rect 6593 3782 6623 3834
rect 6623 3782 6649 3834
rect 6353 3780 6409 3782
rect 6433 3780 6489 3782
rect 6513 3780 6569 3782
rect 6593 3780 6649 3782
rect 6353 2746 6409 2748
rect 6433 2746 6489 2748
rect 6513 2746 6569 2748
rect 6593 2746 6649 2748
rect 6353 2694 6379 2746
rect 6379 2694 6409 2746
rect 6433 2694 6443 2746
rect 6443 2694 6489 2746
rect 6513 2694 6559 2746
rect 6559 2694 6569 2746
rect 6593 2694 6623 2746
rect 6623 2694 6649 2746
rect 6353 2692 6409 2694
rect 6433 2692 6489 2694
rect 6513 2692 6569 2694
rect 6593 2692 6649 2694
rect 9052 6554 9108 6556
rect 9132 6554 9188 6556
rect 9212 6554 9268 6556
rect 9292 6554 9348 6556
rect 9052 6502 9078 6554
rect 9078 6502 9108 6554
rect 9132 6502 9142 6554
rect 9142 6502 9188 6554
rect 9212 6502 9258 6554
rect 9258 6502 9268 6554
rect 9292 6502 9322 6554
rect 9322 6502 9348 6554
rect 9052 6500 9108 6502
rect 9132 6500 9188 6502
rect 9212 6500 9268 6502
rect 9292 6500 9348 6502
rect 9052 5466 9108 5468
rect 9132 5466 9188 5468
rect 9212 5466 9268 5468
rect 9292 5466 9348 5468
rect 9052 5414 9078 5466
rect 9078 5414 9108 5466
rect 9132 5414 9142 5466
rect 9142 5414 9188 5466
rect 9212 5414 9258 5466
rect 9258 5414 9268 5466
rect 9292 5414 9322 5466
rect 9322 5414 9348 5466
rect 9052 5412 9108 5414
rect 9132 5412 9188 5414
rect 9212 5412 9268 5414
rect 9292 5412 9348 5414
rect 11750 16890 11806 16892
rect 11830 16890 11886 16892
rect 11910 16890 11966 16892
rect 11990 16890 12046 16892
rect 11750 16838 11776 16890
rect 11776 16838 11806 16890
rect 11830 16838 11840 16890
rect 11840 16838 11886 16890
rect 11910 16838 11956 16890
rect 11956 16838 11966 16890
rect 11990 16838 12020 16890
rect 12020 16838 12046 16890
rect 11750 16836 11806 16838
rect 11830 16836 11886 16838
rect 11910 16836 11966 16838
rect 11990 16836 12046 16838
rect 11750 15802 11806 15804
rect 11830 15802 11886 15804
rect 11910 15802 11966 15804
rect 11990 15802 12046 15804
rect 11750 15750 11776 15802
rect 11776 15750 11806 15802
rect 11830 15750 11840 15802
rect 11840 15750 11886 15802
rect 11910 15750 11956 15802
rect 11956 15750 11966 15802
rect 11990 15750 12020 15802
rect 12020 15750 12046 15802
rect 11750 15748 11806 15750
rect 11830 15748 11886 15750
rect 11910 15748 11966 15750
rect 11990 15748 12046 15750
rect 11750 14714 11806 14716
rect 11830 14714 11886 14716
rect 11910 14714 11966 14716
rect 11990 14714 12046 14716
rect 11750 14662 11776 14714
rect 11776 14662 11806 14714
rect 11830 14662 11840 14714
rect 11840 14662 11886 14714
rect 11910 14662 11956 14714
rect 11956 14662 11966 14714
rect 11990 14662 12020 14714
rect 12020 14662 12046 14714
rect 11750 14660 11806 14662
rect 11830 14660 11886 14662
rect 11910 14660 11966 14662
rect 11990 14660 12046 14662
rect 11750 13626 11806 13628
rect 11830 13626 11886 13628
rect 11910 13626 11966 13628
rect 11990 13626 12046 13628
rect 11750 13574 11776 13626
rect 11776 13574 11806 13626
rect 11830 13574 11840 13626
rect 11840 13574 11886 13626
rect 11910 13574 11956 13626
rect 11956 13574 11966 13626
rect 11990 13574 12020 13626
rect 12020 13574 12046 13626
rect 11750 13572 11806 13574
rect 11830 13572 11886 13574
rect 11910 13572 11966 13574
rect 11990 13572 12046 13574
rect 11750 12538 11806 12540
rect 11830 12538 11886 12540
rect 11910 12538 11966 12540
rect 11990 12538 12046 12540
rect 11750 12486 11776 12538
rect 11776 12486 11806 12538
rect 11830 12486 11840 12538
rect 11840 12486 11886 12538
rect 11910 12486 11956 12538
rect 11956 12486 11966 12538
rect 11990 12486 12020 12538
rect 12020 12486 12046 12538
rect 11750 12484 11806 12486
rect 11830 12484 11886 12486
rect 11910 12484 11966 12486
rect 11990 12484 12046 12486
rect 11750 11450 11806 11452
rect 11830 11450 11886 11452
rect 11910 11450 11966 11452
rect 11990 11450 12046 11452
rect 11750 11398 11776 11450
rect 11776 11398 11806 11450
rect 11830 11398 11840 11450
rect 11840 11398 11886 11450
rect 11910 11398 11956 11450
rect 11956 11398 11966 11450
rect 11990 11398 12020 11450
rect 12020 11398 12046 11450
rect 11750 11396 11806 11398
rect 11830 11396 11886 11398
rect 11910 11396 11966 11398
rect 11990 11396 12046 11398
rect 11750 10362 11806 10364
rect 11830 10362 11886 10364
rect 11910 10362 11966 10364
rect 11990 10362 12046 10364
rect 11750 10310 11776 10362
rect 11776 10310 11806 10362
rect 11830 10310 11840 10362
rect 11840 10310 11886 10362
rect 11910 10310 11956 10362
rect 11956 10310 11966 10362
rect 11990 10310 12020 10362
rect 12020 10310 12046 10362
rect 11750 10308 11806 10310
rect 11830 10308 11886 10310
rect 11910 10308 11966 10310
rect 11990 10308 12046 10310
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14609 17434 14665 17436
rect 14689 17434 14745 17436
rect 14449 17382 14475 17434
rect 14475 17382 14505 17434
rect 14529 17382 14539 17434
rect 14539 17382 14585 17434
rect 14609 17382 14655 17434
rect 14655 17382 14665 17434
rect 14689 17382 14719 17434
rect 14719 17382 14745 17434
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14609 17380 14665 17382
rect 14689 17380 14745 17382
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14609 16346 14665 16348
rect 14689 16346 14745 16348
rect 14449 16294 14475 16346
rect 14475 16294 14505 16346
rect 14529 16294 14539 16346
rect 14539 16294 14585 16346
rect 14609 16294 14655 16346
rect 14655 16294 14665 16346
rect 14689 16294 14719 16346
rect 14719 16294 14745 16346
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14609 16292 14665 16294
rect 14689 16292 14745 16294
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14609 15258 14665 15260
rect 14689 15258 14745 15260
rect 14449 15206 14475 15258
rect 14475 15206 14505 15258
rect 14529 15206 14539 15258
rect 14539 15206 14585 15258
rect 14609 15206 14655 15258
rect 14655 15206 14665 15258
rect 14689 15206 14719 15258
rect 14719 15206 14745 15258
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 14609 15204 14665 15206
rect 14689 15204 14745 15206
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14609 14170 14665 14172
rect 14689 14170 14745 14172
rect 14449 14118 14475 14170
rect 14475 14118 14505 14170
rect 14529 14118 14539 14170
rect 14539 14118 14585 14170
rect 14609 14118 14655 14170
rect 14655 14118 14665 14170
rect 14689 14118 14719 14170
rect 14719 14118 14745 14170
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14609 14116 14665 14118
rect 14689 14116 14745 14118
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14609 13082 14665 13084
rect 14689 13082 14745 13084
rect 14449 13030 14475 13082
rect 14475 13030 14505 13082
rect 14529 13030 14539 13082
rect 14539 13030 14585 13082
rect 14609 13030 14655 13082
rect 14655 13030 14665 13082
rect 14689 13030 14719 13082
rect 14719 13030 14745 13082
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14609 13028 14665 13030
rect 14689 13028 14745 13030
rect 16762 17060 16818 17096
rect 16762 17040 16764 17060
rect 16764 17040 16816 17060
rect 16816 17040 16818 17060
rect 16762 15000 16818 15056
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14609 11994 14665 11996
rect 14689 11994 14745 11996
rect 14449 11942 14475 11994
rect 14475 11942 14505 11994
rect 14529 11942 14539 11994
rect 14539 11942 14585 11994
rect 14609 11942 14655 11994
rect 14655 11942 14665 11994
rect 14689 11942 14719 11994
rect 14719 11942 14745 11994
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14609 11940 14665 11942
rect 14689 11940 14745 11942
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14609 10906 14665 10908
rect 14689 10906 14745 10908
rect 14449 10854 14475 10906
rect 14475 10854 14505 10906
rect 14529 10854 14539 10906
rect 14539 10854 14585 10906
rect 14609 10854 14655 10906
rect 14655 10854 14665 10906
rect 14689 10854 14719 10906
rect 14719 10854 14745 10906
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14609 10852 14665 10854
rect 14689 10852 14745 10854
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14609 9818 14665 9820
rect 14689 9818 14745 9820
rect 14449 9766 14475 9818
rect 14475 9766 14505 9818
rect 14529 9766 14539 9818
rect 14539 9766 14585 9818
rect 14609 9766 14655 9818
rect 14655 9766 14665 9818
rect 14689 9766 14719 9818
rect 14719 9766 14745 9818
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14609 9764 14665 9766
rect 14689 9764 14745 9766
rect 9052 4378 9108 4380
rect 9132 4378 9188 4380
rect 9212 4378 9268 4380
rect 9292 4378 9348 4380
rect 9052 4326 9078 4378
rect 9078 4326 9108 4378
rect 9132 4326 9142 4378
rect 9142 4326 9188 4378
rect 9212 4326 9258 4378
rect 9258 4326 9268 4378
rect 9292 4326 9322 4378
rect 9322 4326 9348 4378
rect 9052 4324 9108 4326
rect 9132 4324 9188 4326
rect 9212 4324 9268 4326
rect 9292 4324 9348 4326
rect 9052 3290 9108 3292
rect 9132 3290 9188 3292
rect 9212 3290 9268 3292
rect 9292 3290 9348 3292
rect 9052 3238 9078 3290
rect 9078 3238 9108 3290
rect 9132 3238 9142 3290
rect 9142 3238 9188 3290
rect 9212 3238 9258 3290
rect 9258 3238 9268 3290
rect 9292 3238 9322 3290
rect 9322 3238 9348 3290
rect 9052 3236 9108 3238
rect 9132 3236 9188 3238
rect 9212 3236 9268 3238
rect 9292 3236 9348 3238
rect 11750 9274 11806 9276
rect 11830 9274 11886 9276
rect 11910 9274 11966 9276
rect 11990 9274 12046 9276
rect 11750 9222 11776 9274
rect 11776 9222 11806 9274
rect 11830 9222 11840 9274
rect 11840 9222 11886 9274
rect 11910 9222 11956 9274
rect 11956 9222 11966 9274
rect 11990 9222 12020 9274
rect 12020 9222 12046 9274
rect 11750 9220 11806 9222
rect 11830 9220 11886 9222
rect 11910 9220 11966 9222
rect 11990 9220 12046 9222
rect 11750 8186 11806 8188
rect 11830 8186 11886 8188
rect 11910 8186 11966 8188
rect 11990 8186 12046 8188
rect 11750 8134 11776 8186
rect 11776 8134 11806 8186
rect 11830 8134 11840 8186
rect 11840 8134 11886 8186
rect 11910 8134 11956 8186
rect 11956 8134 11966 8186
rect 11990 8134 12020 8186
rect 12020 8134 12046 8186
rect 11750 8132 11806 8134
rect 11830 8132 11886 8134
rect 11910 8132 11966 8134
rect 11990 8132 12046 8134
rect 11750 7098 11806 7100
rect 11830 7098 11886 7100
rect 11910 7098 11966 7100
rect 11990 7098 12046 7100
rect 11750 7046 11776 7098
rect 11776 7046 11806 7098
rect 11830 7046 11840 7098
rect 11840 7046 11886 7098
rect 11910 7046 11956 7098
rect 11956 7046 11966 7098
rect 11990 7046 12020 7098
rect 12020 7046 12046 7098
rect 11750 7044 11806 7046
rect 11830 7044 11886 7046
rect 11910 7044 11966 7046
rect 11990 7044 12046 7046
rect 11750 6010 11806 6012
rect 11830 6010 11886 6012
rect 11910 6010 11966 6012
rect 11990 6010 12046 6012
rect 11750 5958 11776 6010
rect 11776 5958 11806 6010
rect 11830 5958 11840 6010
rect 11840 5958 11886 6010
rect 11910 5958 11956 6010
rect 11956 5958 11966 6010
rect 11990 5958 12020 6010
rect 12020 5958 12046 6010
rect 11750 5956 11806 5958
rect 11830 5956 11886 5958
rect 11910 5956 11966 5958
rect 11990 5956 12046 5958
rect 11750 4922 11806 4924
rect 11830 4922 11886 4924
rect 11910 4922 11966 4924
rect 11990 4922 12046 4924
rect 11750 4870 11776 4922
rect 11776 4870 11806 4922
rect 11830 4870 11840 4922
rect 11840 4870 11886 4922
rect 11910 4870 11956 4922
rect 11956 4870 11966 4922
rect 11990 4870 12020 4922
rect 12020 4870 12046 4922
rect 11750 4868 11806 4870
rect 11830 4868 11886 4870
rect 11910 4868 11966 4870
rect 11990 4868 12046 4870
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14609 8730 14665 8732
rect 14689 8730 14745 8732
rect 14449 8678 14475 8730
rect 14475 8678 14505 8730
rect 14529 8678 14539 8730
rect 14539 8678 14585 8730
rect 14609 8678 14655 8730
rect 14655 8678 14665 8730
rect 14689 8678 14719 8730
rect 14719 8678 14745 8730
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14609 8676 14665 8678
rect 14689 8676 14745 8678
rect 16394 10920 16450 10976
rect 16762 12960 16818 13016
rect 16762 8880 16818 8936
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14609 7642 14665 7644
rect 14689 7642 14745 7644
rect 14449 7590 14475 7642
rect 14475 7590 14505 7642
rect 14529 7590 14539 7642
rect 14539 7590 14585 7642
rect 14609 7590 14655 7642
rect 14655 7590 14665 7642
rect 14689 7590 14719 7642
rect 14719 7590 14745 7642
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14609 7588 14665 7590
rect 14689 7588 14745 7590
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14609 6554 14665 6556
rect 14689 6554 14745 6556
rect 14449 6502 14475 6554
rect 14475 6502 14505 6554
rect 14529 6502 14539 6554
rect 14539 6502 14585 6554
rect 14609 6502 14655 6554
rect 14655 6502 14665 6554
rect 14689 6502 14719 6554
rect 14719 6502 14745 6554
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14609 6500 14665 6502
rect 14689 6500 14745 6502
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14609 5466 14665 5468
rect 14689 5466 14745 5468
rect 14449 5414 14475 5466
rect 14475 5414 14505 5466
rect 14529 5414 14539 5466
rect 14539 5414 14585 5466
rect 14609 5414 14655 5466
rect 14655 5414 14665 5466
rect 14689 5414 14719 5466
rect 14719 5414 14745 5466
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 14609 5412 14665 5414
rect 14689 5412 14745 5414
rect 9052 2202 9108 2204
rect 9132 2202 9188 2204
rect 9212 2202 9268 2204
rect 9292 2202 9348 2204
rect 9052 2150 9078 2202
rect 9078 2150 9108 2202
rect 9132 2150 9142 2202
rect 9142 2150 9188 2202
rect 9212 2150 9258 2202
rect 9258 2150 9268 2202
rect 9292 2150 9322 2202
rect 9322 2150 9348 2202
rect 9052 2148 9108 2150
rect 9132 2148 9188 2150
rect 9212 2148 9268 2150
rect 9292 2148 9348 2150
rect 11750 3834 11806 3836
rect 11830 3834 11886 3836
rect 11910 3834 11966 3836
rect 11990 3834 12046 3836
rect 11750 3782 11776 3834
rect 11776 3782 11806 3834
rect 11830 3782 11840 3834
rect 11840 3782 11886 3834
rect 11910 3782 11956 3834
rect 11956 3782 11966 3834
rect 11990 3782 12020 3834
rect 12020 3782 12046 3834
rect 11750 3780 11806 3782
rect 11830 3780 11886 3782
rect 11910 3780 11966 3782
rect 11990 3780 12046 3782
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14609 4378 14665 4380
rect 14689 4378 14745 4380
rect 14449 4326 14475 4378
rect 14475 4326 14505 4378
rect 14529 4326 14539 4378
rect 14539 4326 14585 4378
rect 14609 4326 14655 4378
rect 14655 4326 14665 4378
rect 14689 4326 14719 4378
rect 14719 4326 14745 4378
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14609 4324 14665 4326
rect 14689 4324 14745 4326
rect 11750 2746 11806 2748
rect 11830 2746 11886 2748
rect 11910 2746 11966 2748
rect 11990 2746 12046 2748
rect 11750 2694 11776 2746
rect 11776 2694 11806 2746
rect 11830 2694 11840 2746
rect 11840 2694 11886 2746
rect 11910 2694 11956 2746
rect 11956 2694 11966 2746
rect 11990 2694 12020 2746
rect 12020 2694 12046 2746
rect 11750 2692 11806 2694
rect 11830 2692 11886 2694
rect 11910 2692 11966 2694
rect 11990 2692 12046 2694
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14609 3290 14665 3292
rect 14689 3290 14745 3292
rect 14449 3238 14475 3290
rect 14475 3238 14505 3290
rect 14529 3238 14539 3290
rect 14539 3238 14585 3290
rect 14609 3238 14655 3290
rect 14655 3238 14665 3290
rect 14689 3238 14719 3290
rect 14719 3238 14745 3290
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14609 3236 14665 3238
rect 14689 3236 14745 3238
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14609 2202 14665 2204
rect 14689 2202 14745 2204
rect 14449 2150 14475 2202
rect 14475 2150 14505 2202
rect 14529 2150 14539 2202
rect 14539 2150 14585 2202
rect 14609 2150 14655 2202
rect 14655 2150 14665 2202
rect 14689 2150 14719 2202
rect 14719 2150 14745 2202
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
rect 14609 2148 14665 2150
rect 14689 2148 14745 2150
rect 16946 6860 17002 6896
rect 16946 6840 16948 6860
rect 16948 6840 17000 6860
rect 17000 6840 17002 6860
rect 16946 4800 17002 4856
rect 16486 2760 16542 2816
rect 16762 720 16818 776
<< metal3 >>
rect 15561 19138 15627 19141
rect 17660 19138 18460 19168
rect 15561 19136 18460 19138
rect 15561 19080 15566 19136
rect 15622 19080 18460 19136
rect 15561 19078 18460 19080
rect 15561 19075 15627 19078
rect 17660 19048 18460 19078
rect 0 18458 800 18488
rect 1485 18458 1551 18461
rect 0 18456 1551 18458
rect 0 18400 1490 18456
rect 1546 18400 1551 18456
rect 0 18398 1551 18400
rect 0 18368 800 18398
rect 1485 18395 1551 18398
rect 6341 17984 6661 17985
rect 6341 17920 6349 17984
rect 6413 17920 6429 17984
rect 6493 17920 6509 17984
rect 6573 17920 6589 17984
rect 6653 17920 6661 17984
rect 6341 17919 6661 17920
rect 11738 17984 12058 17985
rect 11738 17920 11746 17984
rect 11810 17920 11826 17984
rect 11890 17920 11906 17984
rect 11970 17920 11986 17984
rect 12050 17920 12058 17984
rect 11738 17919 12058 17920
rect 3642 17440 3962 17441
rect 3642 17376 3650 17440
rect 3714 17376 3730 17440
rect 3794 17376 3810 17440
rect 3874 17376 3890 17440
rect 3954 17376 3962 17440
rect 3642 17375 3962 17376
rect 9040 17440 9360 17441
rect 9040 17376 9048 17440
rect 9112 17376 9128 17440
rect 9192 17376 9208 17440
rect 9272 17376 9288 17440
rect 9352 17376 9360 17440
rect 9040 17375 9360 17376
rect 14437 17440 14757 17441
rect 14437 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14605 17440
rect 14669 17376 14685 17440
rect 14749 17376 14757 17440
rect 14437 17375 14757 17376
rect 16757 17098 16823 17101
rect 17660 17098 18460 17128
rect 16757 17096 18460 17098
rect 16757 17040 16762 17096
rect 16818 17040 18460 17096
rect 16757 17038 18460 17040
rect 16757 17035 16823 17038
rect 17660 17008 18460 17038
rect 6341 16896 6661 16897
rect 6341 16832 6349 16896
rect 6413 16832 6429 16896
rect 6493 16832 6509 16896
rect 6573 16832 6589 16896
rect 6653 16832 6661 16896
rect 6341 16831 6661 16832
rect 11738 16896 12058 16897
rect 11738 16832 11746 16896
rect 11810 16832 11826 16896
rect 11890 16832 11906 16896
rect 11970 16832 11986 16896
rect 12050 16832 12058 16896
rect 11738 16831 12058 16832
rect 0 16418 800 16448
rect 1393 16418 1459 16421
rect 0 16416 1459 16418
rect 0 16360 1398 16416
rect 1454 16360 1459 16416
rect 0 16358 1459 16360
rect 0 16328 800 16358
rect 1393 16355 1459 16358
rect 3642 16352 3962 16353
rect 3642 16288 3650 16352
rect 3714 16288 3730 16352
rect 3794 16288 3810 16352
rect 3874 16288 3890 16352
rect 3954 16288 3962 16352
rect 3642 16287 3962 16288
rect 9040 16352 9360 16353
rect 9040 16288 9048 16352
rect 9112 16288 9128 16352
rect 9192 16288 9208 16352
rect 9272 16288 9288 16352
rect 9352 16288 9360 16352
rect 9040 16287 9360 16288
rect 14437 16352 14757 16353
rect 14437 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14605 16352
rect 14669 16288 14685 16352
rect 14749 16288 14757 16352
rect 14437 16287 14757 16288
rect 6341 15808 6661 15809
rect 6341 15744 6349 15808
rect 6413 15744 6429 15808
rect 6493 15744 6509 15808
rect 6573 15744 6589 15808
rect 6653 15744 6661 15808
rect 6341 15743 6661 15744
rect 11738 15808 12058 15809
rect 11738 15744 11746 15808
rect 11810 15744 11826 15808
rect 11890 15744 11906 15808
rect 11970 15744 11986 15808
rect 12050 15744 12058 15808
rect 11738 15743 12058 15744
rect 3642 15264 3962 15265
rect 3642 15200 3650 15264
rect 3714 15200 3730 15264
rect 3794 15200 3810 15264
rect 3874 15200 3890 15264
rect 3954 15200 3962 15264
rect 3642 15199 3962 15200
rect 9040 15264 9360 15265
rect 9040 15200 9048 15264
rect 9112 15200 9128 15264
rect 9192 15200 9208 15264
rect 9272 15200 9288 15264
rect 9352 15200 9360 15264
rect 9040 15199 9360 15200
rect 14437 15264 14757 15265
rect 14437 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14605 15264
rect 14669 15200 14685 15264
rect 14749 15200 14757 15264
rect 14437 15199 14757 15200
rect 2865 15058 2931 15061
rect 3877 15058 3943 15061
rect 4705 15058 4771 15061
rect 2865 15056 4771 15058
rect 2865 15000 2870 15056
rect 2926 15000 3882 15056
rect 3938 15000 4710 15056
rect 4766 15000 4771 15056
rect 2865 14998 4771 15000
rect 2865 14995 2931 14998
rect 3877 14995 3943 14998
rect 4705 14995 4771 14998
rect 16757 15058 16823 15061
rect 17660 15058 18460 15088
rect 16757 15056 18460 15058
rect 16757 15000 16762 15056
rect 16818 15000 18460 15056
rect 16757 14998 18460 15000
rect 16757 14995 16823 14998
rect 17660 14968 18460 14998
rect 3141 14922 3207 14925
rect 3693 14922 3759 14925
rect 3141 14920 3759 14922
rect 3141 14864 3146 14920
rect 3202 14864 3698 14920
rect 3754 14864 3759 14920
rect 3141 14862 3759 14864
rect 3141 14859 3207 14862
rect 3693 14859 3759 14862
rect 6341 14720 6661 14721
rect 6341 14656 6349 14720
rect 6413 14656 6429 14720
rect 6493 14656 6509 14720
rect 6573 14656 6589 14720
rect 6653 14656 6661 14720
rect 6341 14655 6661 14656
rect 11738 14720 12058 14721
rect 11738 14656 11746 14720
rect 11810 14656 11826 14720
rect 11890 14656 11906 14720
rect 11970 14656 11986 14720
rect 12050 14656 12058 14720
rect 11738 14655 12058 14656
rect 0 14378 800 14408
rect 1393 14378 1459 14381
rect 0 14376 1459 14378
rect 0 14320 1398 14376
rect 1454 14320 1459 14376
rect 0 14318 1459 14320
rect 0 14288 800 14318
rect 1393 14315 1459 14318
rect 3642 14176 3962 14177
rect 3642 14112 3650 14176
rect 3714 14112 3730 14176
rect 3794 14112 3810 14176
rect 3874 14112 3890 14176
rect 3954 14112 3962 14176
rect 3642 14111 3962 14112
rect 9040 14176 9360 14177
rect 9040 14112 9048 14176
rect 9112 14112 9128 14176
rect 9192 14112 9208 14176
rect 9272 14112 9288 14176
rect 9352 14112 9360 14176
rect 9040 14111 9360 14112
rect 14437 14176 14757 14177
rect 14437 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14605 14176
rect 14669 14112 14685 14176
rect 14749 14112 14757 14176
rect 14437 14111 14757 14112
rect 6341 13632 6661 13633
rect 6341 13568 6349 13632
rect 6413 13568 6429 13632
rect 6493 13568 6509 13632
rect 6573 13568 6589 13632
rect 6653 13568 6661 13632
rect 6341 13567 6661 13568
rect 11738 13632 12058 13633
rect 11738 13568 11746 13632
rect 11810 13568 11826 13632
rect 11890 13568 11906 13632
rect 11970 13568 11986 13632
rect 12050 13568 12058 13632
rect 11738 13567 12058 13568
rect 4061 13290 4127 13293
rect 4061 13288 4170 13290
rect 4061 13232 4066 13288
rect 4122 13232 4170 13288
rect 4061 13227 4170 13232
rect 3642 13088 3962 13089
rect 3642 13024 3650 13088
rect 3714 13024 3730 13088
rect 3794 13024 3810 13088
rect 3874 13024 3890 13088
rect 3954 13024 3962 13088
rect 3642 13023 3962 13024
rect 3877 12882 3943 12885
rect 4110 12882 4170 13227
rect 9040 13088 9360 13089
rect 9040 13024 9048 13088
rect 9112 13024 9128 13088
rect 9192 13024 9208 13088
rect 9272 13024 9288 13088
rect 9352 13024 9360 13088
rect 9040 13023 9360 13024
rect 14437 13088 14757 13089
rect 14437 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14605 13088
rect 14669 13024 14685 13088
rect 14749 13024 14757 13088
rect 14437 13023 14757 13024
rect 16757 13018 16823 13021
rect 17660 13018 18460 13048
rect 16757 13016 18460 13018
rect 16757 12960 16762 13016
rect 16818 12960 18460 13016
rect 16757 12958 18460 12960
rect 16757 12955 16823 12958
rect 17660 12928 18460 12958
rect 3877 12880 4170 12882
rect 3877 12824 3882 12880
rect 3938 12824 4170 12880
rect 3877 12822 4170 12824
rect 5901 12882 5967 12885
rect 7189 12882 7255 12885
rect 5901 12880 7255 12882
rect 5901 12824 5906 12880
rect 5962 12824 7194 12880
rect 7250 12824 7255 12880
rect 5901 12822 7255 12824
rect 3877 12819 3943 12822
rect 5901 12819 5967 12822
rect 7189 12819 7255 12822
rect 6341 12544 6661 12545
rect 6341 12480 6349 12544
rect 6413 12480 6429 12544
rect 6493 12480 6509 12544
rect 6573 12480 6589 12544
rect 6653 12480 6661 12544
rect 6341 12479 6661 12480
rect 11738 12544 12058 12545
rect 11738 12480 11746 12544
rect 11810 12480 11826 12544
rect 11890 12480 11906 12544
rect 11970 12480 11986 12544
rect 12050 12480 12058 12544
rect 11738 12479 12058 12480
rect 0 12338 800 12368
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 3642 12000 3962 12001
rect 3642 11936 3650 12000
rect 3714 11936 3730 12000
rect 3794 11936 3810 12000
rect 3874 11936 3890 12000
rect 3954 11936 3962 12000
rect 3642 11935 3962 11936
rect 9040 12000 9360 12001
rect 9040 11936 9048 12000
rect 9112 11936 9128 12000
rect 9192 11936 9208 12000
rect 9272 11936 9288 12000
rect 9352 11936 9360 12000
rect 9040 11935 9360 11936
rect 14437 12000 14757 12001
rect 14437 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14605 12000
rect 14669 11936 14685 12000
rect 14749 11936 14757 12000
rect 14437 11935 14757 11936
rect 6341 11456 6661 11457
rect 6341 11392 6349 11456
rect 6413 11392 6429 11456
rect 6493 11392 6509 11456
rect 6573 11392 6589 11456
rect 6653 11392 6661 11456
rect 6341 11391 6661 11392
rect 11738 11456 12058 11457
rect 11738 11392 11746 11456
rect 11810 11392 11826 11456
rect 11890 11392 11906 11456
rect 11970 11392 11986 11456
rect 12050 11392 12058 11456
rect 11738 11391 12058 11392
rect 16389 10978 16455 10981
rect 17660 10978 18460 11008
rect 16389 10976 18460 10978
rect 16389 10920 16394 10976
rect 16450 10920 18460 10976
rect 16389 10918 18460 10920
rect 16389 10915 16455 10918
rect 3642 10912 3962 10913
rect 3642 10848 3650 10912
rect 3714 10848 3730 10912
rect 3794 10848 3810 10912
rect 3874 10848 3890 10912
rect 3954 10848 3962 10912
rect 3642 10847 3962 10848
rect 9040 10912 9360 10913
rect 9040 10848 9048 10912
rect 9112 10848 9128 10912
rect 9192 10848 9208 10912
rect 9272 10848 9288 10912
rect 9352 10848 9360 10912
rect 9040 10847 9360 10848
rect 14437 10912 14757 10913
rect 14437 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14605 10912
rect 14669 10848 14685 10912
rect 14749 10848 14757 10912
rect 17660 10888 18460 10918
rect 14437 10847 14757 10848
rect 6341 10368 6661 10369
rect 0 10298 800 10328
rect 6341 10304 6349 10368
rect 6413 10304 6429 10368
rect 6493 10304 6509 10368
rect 6573 10304 6589 10368
rect 6653 10304 6661 10368
rect 6341 10303 6661 10304
rect 11738 10368 12058 10369
rect 11738 10304 11746 10368
rect 11810 10304 11826 10368
rect 11890 10304 11906 10368
rect 11970 10304 11986 10368
rect 12050 10304 12058 10368
rect 11738 10303 12058 10304
rect 1485 10298 1551 10301
rect 0 10296 1551 10298
rect 0 10240 1490 10296
rect 1546 10240 1551 10296
rect 0 10238 1551 10240
rect 0 10208 800 10238
rect 1485 10235 1551 10238
rect 3642 9824 3962 9825
rect 3642 9760 3650 9824
rect 3714 9760 3730 9824
rect 3794 9760 3810 9824
rect 3874 9760 3890 9824
rect 3954 9760 3962 9824
rect 3642 9759 3962 9760
rect 9040 9824 9360 9825
rect 9040 9760 9048 9824
rect 9112 9760 9128 9824
rect 9192 9760 9208 9824
rect 9272 9760 9288 9824
rect 9352 9760 9360 9824
rect 9040 9759 9360 9760
rect 14437 9824 14757 9825
rect 14437 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14605 9824
rect 14669 9760 14685 9824
rect 14749 9760 14757 9824
rect 14437 9759 14757 9760
rect 7557 9482 7623 9485
rect 7741 9482 7807 9485
rect 8293 9482 8359 9485
rect 7557 9480 8359 9482
rect 7557 9424 7562 9480
rect 7618 9424 7746 9480
rect 7802 9424 8298 9480
rect 8354 9424 8359 9480
rect 7557 9422 8359 9424
rect 7557 9419 7623 9422
rect 7741 9419 7807 9422
rect 8293 9419 8359 9422
rect 6341 9280 6661 9281
rect 6341 9216 6349 9280
rect 6413 9216 6429 9280
rect 6493 9216 6509 9280
rect 6573 9216 6589 9280
rect 6653 9216 6661 9280
rect 6341 9215 6661 9216
rect 11738 9280 12058 9281
rect 11738 9216 11746 9280
rect 11810 9216 11826 9280
rect 11890 9216 11906 9280
rect 11970 9216 11986 9280
rect 12050 9216 12058 9280
rect 11738 9215 12058 9216
rect 16757 8938 16823 8941
rect 17660 8938 18460 8968
rect 16757 8936 18460 8938
rect 16757 8880 16762 8936
rect 16818 8880 18460 8936
rect 16757 8878 18460 8880
rect 16757 8875 16823 8878
rect 17660 8848 18460 8878
rect 3642 8736 3962 8737
rect 3642 8672 3650 8736
rect 3714 8672 3730 8736
rect 3794 8672 3810 8736
rect 3874 8672 3890 8736
rect 3954 8672 3962 8736
rect 3642 8671 3962 8672
rect 9040 8736 9360 8737
rect 9040 8672 9048 8736
rect 9112 8672 9128 8736
rect 9192 8672 9208 8736
rect 9272 8672 9288 8736
rect 9352 8672 9360 8736
rect 9040 8671 9360 8672
rect 14437 8736 14757 8737
rect 14437 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14605 8736
rect 14669 8672 14685 8736
rect 14749 8672 14757 8736
rect 14437 8671 14757 8672
rect 5993 8394 6059 8397
rect 7649 8394 7715 8397
rect 5993 8392 7715 8394
rect 5993 8336 5998 8392
rect 6054 8336 7654 8392
rect 7710 8336 7715 8392
rect 5993 8334 7715 8336
rect 5993 8331 6059 8334
rect 7649 8331 7715 8334
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 6341 8192 6661 8193
rect 6341 8128 6349 8192
rect 6413 8128 6429 8192
rect 6493 8128 6509 8192
rect 6573 8128 6589 8192
rect 6653 8128 6661 8192
rect 6341 8127 6661 8128
rect 11738 8192 12058 8193
rect 11738 8128 11746 8192
rect 11810 8128 11826 8192
rect 11890 8128 11906 8192
rect 11970 8128 11986 8192
rect 12050 8128 12058 8192
rect 11738 8127 12058 8128
rect 3642 7648 3962 7649
rect 3642 7584 3650 7648
rect 3714 7584 3730 7648
rect 3794 7584 3810 7648
rect 3874 7584 3890 7648
rect 3954 7584 3962 7648
rect 3642 7583 3962 7584
rect 9040 7648 9360 7649
rect 9040 7584 9048 7648
rect 9112 7584 9128 7648
rect 9192 7584 9208 7648
rect 9272 7584 9288 7648
rect 9352 7584 9360 7648
rect 9040 7583 9360 7584
rect 14437 7648 14757 7649
rect 14437 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14605 7648
rect 14669 7584 14685 7648
rect 14749 7584 14757 7648
rect 14437 7583 14757 7584
rect 6341 7104 6661 7105
rect 6341 7040 6349 7104
rect 6413 7040 6429 7104
rect 6493 7040 6509 7104
rect 6573 7040 6589 7104
rect 6653 7040 6661 7104
rect 6341 7039 6661 7040
rect 11738 7104 12058 7105
rect 11738 7040 11746 7104
rect 11810 7040 11826 7104
rect 11890 7040 11906 7104
rect 11970 7040 11986 7104
rect 12050 7040 12058 7104
rect 11738 7039 12058 7040
rect 16941 6898 17007 6901
rect 17660 6898 18460 6928
rect 16941 6896 18460 6898
rect 16941 6840 16946 6896
rect 17002 6840 18460 6896
rect 16941 6838 18460 6840
rect 16941 6835 17007 6838
rect 17660 6808 18460 6838
rect 3642 6560 3962 6561
rect 3642 6496 3650 6560
rect 3714 6496 3730 6560
rect 3794 6496 3810 6560
rect 3874 6496 3890 6560
rect 3954 6496 3962 6560
rect 3642 6495 3962 6496
rect 9040 6560 9360 6561
rect 9040 6496 9048 6560
rect 9112 6496 9128 6560
rect 9192 6496 9208 6560
rect 9272 6496 9288 6560
rect 9352 6496 9360 6560
rect 9040 6495 9360 6496
rect 14437 6560 14757 6561
rect 14437 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14605 6560
rect 14669 6496 14685 6560
rect 14749 6496 14757 6560
rect 14437 6495 14757 6496
rect 0 6218 800 6248
rect 1393 6218 1459 6221
rect 0 6216 1459 6218
rect 0 6160 1398 6216
rect 1454 6160 1459 6216
rect 0 6158 1459 6160
rect 0 6128 800 6158
rect 1393 6155 1459 6158
rect 6341 6016 6661 6017
rect 6341 5952 6349 6016
rect 6413 5952 6429 6016
rect 6493 5952 6509 6016
rect 6573 5952 6589 6016
rect 6653 5952 6661 6016
rect 6341 5951 6661 5952
rect 11738 6016 12058 6017
rect 11738 5952 11746 6016
rect 11810 5952 11826 6016
rect 11890 5952 11906 6016
rect 11970 5952 11986 6016
rect 12050 5952 12058 6016
rect 11738 5951 12058 5952
rect 3642 5472 3962 5473
rect 3642 5408 3650 5472
rect 3714 5408 3730 5472
rect 3794 5408 3810 5472
rect 3874 5408 3890 5472
rect 3954 5408 3962 5472
rect 3642 5407 3962 5408
rect 9040 5472 9360 5473
rect 9040 5408 9048 5472
rect 9112 5408 9128 5472
rect 9192 5408 9208 5472
rect 9272 5408 9288 5472
rect 9352 5408 9360 5472
rect 9040 5407 9360 5408
rect 14437 5472 14757 5473
rect 14437 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14605 5472
rect 14669 5408 14685 5472
rect 14749 5408 14757 5472
rect 14437 5407 14757 5408
rect 6341 4928 6661 4929
rect 6341 4864 6349 4928
rect 6413 4864 6429 4928
rect 6493 4864 6509 4928
rect 6573 4864 6589 4928
rect 6653 4864 6661 4928
rect 6341 4863 6661 4864
rect 11738 4928 12058 4929
rect 11738 4864 11746 4928
rect 11810 4864 11826 4928
rect 11890 4864 11906 4928
rect 11970 4864 11986 4928
rect 12050 4864 12058 4928
rect 11738 4863 12058 4864
rect 16941 4858 17007 4861
rect 17660 4858 18460 4888
rect 16941 4856 18460 4858
rect 16941 4800 16946 4856
rect 17002 4800 18460 4856
rect 16941 4798 18460 4800
rect 16941 4795 17007 4798
rect 17660 4768 18460 4798
rect 3642 4384 3962 4385
rect 3642 4320 3650 4384
rect 3714 4320 3730 4384
rect 3794 4320 3810 4384
rect 3874 4320 3890 4384
rect 3954 4320 3962 4384
rect 3642 4319 3962 4320
rect 9040 4384 9360 4385
rect 9040 4320 9048 4384
rect 9112 4320 9128 4384
rect 9192 4320 9208 4384
rect 9272 4320 9288 4384
rect 9352 4320 9360 4384
rect 9040 4319 9360 4320
rect 14437 4384 14757 4385
rect 14437 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14605 4384
rect 14669 4320 14685 4384
rect 14749 4320 14757 4384
rect 14437 4319 14757 4320
rect 0 4178 800 4208
rect 1393 4178 1459 4181
rect 0 4176 1459 4178
rect 0 4120 1398 4176
rect 1454 4120 1459 4176
rect 0 4118 1459 4120
rect 0 4088 800 4118
rect 1393 4115 1459 4118
rect 6341 3840 6661 3841
rect 6341 3776 6349 3840
rect 6413 3776 6429 3840
rect 6493 3776 6509 3840
rect 6573 3776 6589 3840
rect 6653 3776 6661 3840
rect 6341 3775 6661 3776
rect 11738 3840 12058 3841
rect 11738 3776 11746 3840
rect 11810 3776 11826 3840
rect 11890 3776 11906 3840
rect 11970 3776 11986 3840
rect 12050 3776 12058 3840
rect 11738 3775 12058 3776
rect 3642 3296 3962 3297
rect 3642 3232 3650 3296
rect 3714 3232 3730 3296
rect 3794 3232 3810 3296
rect 3874 3232 3890 3296
rect 3954 3232 3962 3296
rect 3642 3231 3962 3232
rect 9040 3296 9360 3297
rect 9040 3232 9048 3296
rect 9112 3232 9128 3296
rect 9192 3232 9208 3296
rect 9272 3232 9288 3296
rect 9352 3232 9360 3296
rect 9040 3231 9360 3232
rect 14437 3296 14757 3297
rect 14437 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14605 3296
rect 14669 3232 14685 3296
rect 14749 3232 14757 3296
rect 14437 3231 14757 3232
rect 16481 2818 16547 2821
rect 17660 2818 18460 2848
rect 16481 2816 18460 2818
rect 16481 2760 16486 2816
rect 16542 2760 18460 2816
rect 16481 2758 18460 2760
rect 16481 2755 16547 2758
rect 6341 2752 6661 2753
rect 6341 2688 6349 2752
rect 6413 2688 6429 2752
rect 6493 2688 6509 2752
rect 6573 2688 6589 2752
rect 6653 2688 6661 2752
rect 6341 2687 6661 2688
rect 11738 2752 12058 2753
rect 11738 2688 11746 2752
rect 11810 2688 11826 2752
rect 11890 2688 11906 2752
rect 11970 2688 11986 2752
rect 12050 2688 12058 2752
rect 17660 2728 18460 2758
rect 11738 2687 12058 2688
rect 3642 2208 3962 2209
rect 0 2138 800 2168
rect 3642 2144 3650 2208
rect 3714 2144 3730 2208
rect 3794 2144 3810 2208
rect 3874 2144 3890 2208
rect 3954 2144 3962 2208
rect 3642 2143 3962 2144
rect 9040 2208 9360 2209
rect 9040 2144 9048 2208
rect 9112 2144 9128 2208
rect 9192 2144 9208 2208
rect 9272 2144 9288 2208
rect 9352 2144 9360 2208
rect 9040 2143 9360 2144
rect 14437 2208 14757 2209
rect 14437 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14605 2208
rect 14669 2144 14685 2208
rect 14749 2144 14757 2208
rect 14437 2143 14757 2144
rect 2037 2138 2103 2141
rect 0 2136 2103 2138
rect 0 2080 2042 2136
rect 2098 2080 2103 2136
rect 0 2078 2103 2080
rect 0 2048 800 2078
rect 2037 2075 2103 2078
rect 16757 778 16823 781
rect 17660 778 18460 808
rect 16757 776 18460 778
rect 16757 720 16762 776
rect 16818 720 18460 776
rect 16757 718 18460 720
rect 16757 715 16823 718
rect 17660 688 18460 718
<< via3 >>
rect 6349 17980 6413 17984
rect 6349 17924 6353 17980
rect 6353 17924 6409 17980
rect 6409 17924 6413 17980
rect 6349 17920 6413 17924
rect 6429 17980 6493 17984
rect 6429 17924 6433 17980
rect 6433 17924 6489 17980
rect 6489 17924 6493 17980
rect 6429 17920 6493 17924
rect 6509 17980 6573 17984
rect 6509 17924 6513 17980
rect 6513 17924 6569 17980
rect 6569 17924 6573 17980
rect 6509 17920 6573 17924
rect 6589 17980 6653 17984
rect 6589 17924 6593 17980
rect 6593 17924 6649 17980
rect 6649 17924 6653 17980
rect 6589 17920 6653 17924
rect 11746 17980 11810 17984
rect 11746 17924 11750 17980
rect 11750 17924 11806 17980
rect 11806 17924 11810 17980
rect 11746 17920 11810 17924
rect 11826 17980 11890 17984
rect 11826 17924 11830 17980
rect 11830 17924 11886 17980
rect 11886 17924 11890 17980
rect 11826 17920 11890 17924
rect 11906 17980 11970 17984
rect 11906 17924 11910 17980
rect 11910 17924 11966 17980
rect 11966 17924 11970 17980
rect 11906 17920 11970 17924
rect 11986 17980 12050 17984
rect 11986 17924 11990 17980
rect 11990 17924 12046 17980
rect 12046 17924 12050 17980
rect 11986 17920 12050 17924
rect 3650 17436 3714 17440
rect 3650 17380 3654 17436
rect 3654 17380 3710 17436
rect 3710 17380 3714 17436
rect 3650 17376 3714 17380
rect 3730 17436 3794 17440
rect 3730 17380 3734 17436
rect 3734 17380 3790 17436
rect 3790 17380 3794 17436
rect 3730 17376 3794 17380
rect 3810 17436 3874 17440
rect 3810 17380 3814 17436
rect 3814 17380 3870 17436
rect 3870 17380 3874 17436
rect 3810 17376 3874 17380
rect 3890 17436 3954 17440
rect 3890 17380 3894 17436
rect 3894 17380 3950 17436
rect 3950 17380 3954 17436
rect 3890 17376 3954 17380
rect 9048 17436 9112 17440
rect 9048 17380 9052 17436
rect 9052 17380 9108 17436
rect 9108 17380 9112 17436
rect 9048 17376 9112 17380
rect 9128 17436 9192 17440
rect 9128 17380 9132 17436
rect 9132 17380 9188 17436
rect 9188 17380 9192 17436
rect 9128 17376 9192 17380
rect 9208 17436 9272 17440
rect 9208 17380 9212 17436
rect 9212 17380 9268 17436
rect 9268 17380 9272 17436
rect 9208 17376 9272 17380
rect 9288 17436 9352 17440
rect 9288 17380 9292 17436
rect 9292 17380 9348 17436
rect 9348 17380 9352 17436
rect 9288 17376 9352 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 14605 17436 14669 17440
rect 14605 17380 14609 17436
rect 14609 17380 14665 17436
rect 14665 17380 14669 17436
rect 14605 17376 14669 17380
rect 14685 17436 14749 17440
rect 14685 17380 14689 17436
rect 14689 17380 14745 17436
rect 14745 17380 14749 17436
rect 14685 17376 14749 17380
rect 6349 16892 6413 16896
rect 6349 16836 6353 16892
rect 6353 16836 6409 16892
rect 6409 16836 6413 16892
rect 6349 16832 6413 16836
rect 6429 16892 6493 16896
rect 6429 16836 6433 16892
rect 6433 16836 6489 16892
rect 6489 16836 6493 16892
rect 6429 16832 6493 16836
rect 6509 16892 6573 16896
rect 6509 16836 6513 16892
rect 6513 16836 6569 16892
rect 6569 16836 6573 16892
rect 6509 16832 6573 16836
rect 6589 16892 6653 16896
rect 6589 16836 6593 16892
rect 6593 16836 6649 16892
rect 6649 16836 6653 16892
rect 6589 16832 6653 16836
rect 11746 16892 11810 16896
rect 11746 16836 11750 16892
rect 11750 16836 11806 16892
rect 11806 16836 11810 16892
rect 11746 16832 11810 16836
rect 11826 16892 11890 16896
rect 11826 16836 11830 16892
rect 11830 16836 11886 16892
rect 11886 16836 11890 16892
rect 11826 16832 11890 16836
rect 11906 16892 11970 16896
rect 11906 16836 11910 16892
rect 11910 16836 11966 16892
rect 11966 16836 11970 16892
rect 11906 16832 11970 16836
rect 11986 16892 12050 16896
rect 11986 16836 11990 16892
rect 11990 16836 12046 16892
rect 12046 16836 12050 16892
rect 11986 16832 12050 16836
rect 3650 16348 3714 16352
rect 3650 16292 3654 16348
rect 3654 16292 3710 16348
rect 3710 16292 3714 16348
rect 3650 16288 3714 16292
rect 3730 16348 3794 16352
rect 3730 16292 3734 16348
rect 3734 16292 3790 16348
rect 3790 16292 3794 16348
rect 3730 16288 3794 16292
rect 3810 16348 3874 16352
rect 3810 16292 3814 16348
rect 3814 16292 3870 16348
rect 3870 16292 3874 16348
rect 3810 16288 3874 16292
rect 3890 16348 3954 16352
rect 3890 16292 3894 16348
rect 3894 16292 3950 16348
rect 3950 16292 3954 16348
rect 3890 16288 3954 16292
rect 9048 16348 9112 16352
rect 9048 16292 9052 16348
rect 9052 16292 9108 16348
rect 9108 16292 9112 16348
rect 9048 16288 9112 16292
rect 9128 16348 9192 16352
rect 9128 16292 9132 16348
rect 9132 16292 9188 16348
rect 9188 16292 9192 16348
rect 9128 16288 9192 16292
rect 9208 16348 9272 16352
rect 9208 16292 9212 16348
rect 9212 16292 9268 16348
rect 9268 16292 9272 16348
rect 9208 16288 9272 16292
rect 9288 16348 9352 16352
rect 9288 16292 9292 16348
rect 9292 16292 9348 16348
rect 9348 16292 9352 16348
rect 9288 16288 9352 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 14605 16348 14669 16352
rect 14605 16292 14609 16348
rect 14609 16292 14665 16348
rect 14665 16292 14669 16348
rect 14605 16288 14669 16292
rect 14685 16348 14749 16352
rect 14685 16292 14689 16348
rect 14689 16292 14745 16348
rect 14745 16292 14749 16348
rect 14685 16288 14749 16292
rect 6349 15804 6413 15808
rect 6349 15748 6353 15804
rect 6353 15748 6409 15804
rect 6409 15748 6413 15804
rect 6349 15744 6413 15748
rect 6429 15804 6493 15808
rect 6429 15748 6433 15804
rect 6433 15748 6489 15804
rect 6489 15748 6493 15804
rect 6429 15744 6493 15748
rect 6509 15804 6573 15808
rect 6509 15748 6513 15804
rect 6513 15748 6569 15804
rect 6569 15748 6573 15804
rect 6509 15744 6573 15748
rect 6589 15804 6653 15808
rect 6589 15748 6593 15804
rect 6593 15748 6649 15804
rect 6649 15748 6653 15804
rect 6589 15744 6653 15748
rect 11746 15804 11810 15808
rect 11746 15748 11750 15804
rect 11750 15748 11806 15804
rect 11806 15748 11810 15804
rect 11746 15744 11810 15748
rect 11826 15804 11890 15808
rect 11826 15748 11830 15804
rect 11830 15748 11886 15804
rect 11886 15748 11890 15804
rect 11826 15744 11890 15748
rect 11906 15804 11970 15808
rect 11906 15748 11910 15804
rect 11910 15748 11966 15804
rect 11966 15748 11970 15804
rect 11906 15744 11970 15748
rect 11986 15804 12050 15808
rect 11986 15748 11990 15804
rect 11990 15748 12046 15804
rect 12046 15748 12050 15804
rect 11986 15744 12050 15748
rect 3650 15260 3714 15264
rect 3650 15204 3654 15260
rect 3654 15204 3710 15260
rect 3710 15204 3714 15260
rect 3650 15200 3714 15204
rect 3730 15260 3794 15264
rect 3730 15204 3734 15260
rect 3734 15204 3790 15260
rect 3790 15204 3794 15260
rect 3730 15200 3794 15204
rect 3810 15260 3874 15264
rect 3810 15204 3814 15260
rect 3814 15204 3870 15260
rect 3870 15204 3874 15260
rect 3810 15200 3874 15204
rect 3890 15260 3954 15264
rect 3890 15204 3894 15260
rect 3894 15204 3950 15260
rect 3950 15204 3954 15260
rect 3890 15200 3954 15204
rect 9048 15260 9112 15264
rect 9048 15204 9052 15260
rect 9052 15204 9108 15260
rect 9108 15204 9112 15260
rect 9048 15200 9112 15204
rect 9128 15260 9192 15264
rect 9128 15204 9132 15260
rect 9132 15204 9188 15260
rect 9188 15204 9192 15260
rect 9128 15200 9192 15204
rect 9208 15260 9272 15264
rect 9208 15204 9212 15260
rect 9212 15204 9268 15260
rect 9268 15204 9272 15260
rect 9208 15200 9272 15204
rect 9288 15260 9352 15264
rect 9288 15204 9292 15260
rect 9292 15204 9348 15260
rect 9348 15204 9352 15260
rect 9288 15200 9352 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 14605 15260 14669 15264
rect 14605 15204 14609 15260
rect 14609 15204 14665 15260
rect 14665 15204 14669 15260
rect 14605 15200 14669 15204
rect 14685 15260 14749 15264
rect 14685 15204 14689 15260
rect 14689 15204 14745 15260
rect 14745 15204 14749 15260
rect 14685 15200 14749 15204
rect 6349 14716 6413 14720
rect 6349 14660 6353 14716
rect 6353 14660 6409 14716
rect 6409 14660 6413 14716
rect 6349 14656 6413 14660
rect 6429 14716 6493 14720
rect 6429 14660 6433 14716
rect 6433 14660 6489 14716
rect 6489 14660 6493 14716
rect 6429 14656 6493 14660
rect 6509 14716 6573 14720
rect 6509 14660 6513 14716
rect 6513 14660 6569 14716
rect 6569 14660 6573 14716
rect 6509 14656 6573 14660
rect 6589 14716 6653 14720
rect 6589 14660 6593 14716
rect 6593 14660 6649 14716
rect 6649 14660 6653 14716
rect 6589 14656 6653 14660
rect 11746 14716 11810 14720
rect 11746 14660 11750 14716
rect 11750 14660 11806 14716
rect 11806 14660 11810 14716
rect 11746 14656 11810 14660
rect 11826 14716 11890 14720
rect 11826 14660 11830 14716
rect 11830 14660 11886 14716
rect 11886 14660 11890 14716
rect 11826 14656 11890 14660
rect 11906 14716 11970 14720
rect 11906 14660 11910 14716
rect 11910 14660 11966 14716
rect 11966 14660 11970 14716
rect 11906 14656 11970 14660
rect 11986 14716 12050 14720
rect 11986 14660 11990 14716
rect 11990 14660 12046 14716
rect 12046 14660 12050 14716
rect 11986 14656 12050 14660
rect 3650 14172 3714 14176
rect 3650 14116 3654 14172
rect 3654 14116 3710 14172
rect 3710 14116 3714 14172
rect 3650 14112 3714 14116
rect 3730 14172 3794 14176
rect 3730 14116 3734 14172
rect 3734 14116 3790 14172
rect 3790 14116 3794 14172
rect 3730 14112 3794 14116
rect 3810 14172 3874 14176
rect 3810 14116 3814 14172
rect 3814 14116 3870 14172
rect 3870 14116 3874 14172
rect 3810 14112 3874 14116
rect 3890 14172 3954 14176
rect 3890 14116 3894 14172
rect 3894 14116 3950 14172
rect 3950 14116 3954 14172
rect 3890 14112 3954 14116
rect 9048 14172 9112 14176
rect 9048 14116 9052 14172
rect 9052 14116 9108 14172
rect 9108 14116 9112 14172
rect 9048 14112 9112 14116
rect 9128 14172 9192 14176
rect 9128 14116 9132 14172
rect 9132 14116 9188 14172
rect 9188 14116 9192 14172
rect 9128 14112 9192 14116
rect 9208 14172 9272 14176
rect 9208 14116 9212 14172
rect 9212 14116 9268 14172
rect 9268 14116 9272 14172
rect 9208 14112 9272 14116
rect 9288 14172 9352 14176
rect 9288 14116 9292 14172
rect 9292 14116 9348 14172
rect 9348 14116 9352 14172
rect 9288 14112 9352 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 14605 14172 14669 14176
rect 14605 14116 14609 14172
rect 14609 14116 14665 14172
rect 14665 14116 14669 14172
rect 14605 14112 14669 14116
rect 14685 14172 14749 14176
rect 14685 14116 14689 14172
rect 14689 14116 14745 14172
rect 14745 14116 14749 14172
rect 14685 14112 14749 14116
rect 6349 13628 6413 13632
rect 6349 13572 6353 13628
rect 6353 13572 6409 13628
rect 6409 13572 6413 13628
rect 6349 13568 6413 13572
rect 6429 13628 6493 13632
rect 6429 13572 6433 13628
rect 6433 13572 6489 13628
rect 6489 13572 6493 13628
rect 6429 13568 6493 13572
rect 6509 13628 6573 13632
rect 6509 13572 6513 13628
rect 6513 13572 6569 13628
rect 6569 13572 6573 13628
rect 6509 13568 6573 13572
rect 6589 13628 6653 13632
rect 6589 13572 6593 13628
rect 6593 13572 6649 13628
rect 6649 13572 6653 13628
rect 6589 13568 6653 13572
rect 11746 13628 11810 13632
rect 11746 13572 11750 13628
rect 11750 13572 11806 13628
rect 11806 13572 11810 13628
rect 11746 13568 11810 13572
rect 11826 13628 11890 13632
rect 11826 13572 11830 13628
rect 11830 13572 11886 13628
rect 11886 13572 11890 13628
rect 11826 13568 11890 13572
rect 11906 13628 11970 13632
rect 11906 13572 11910 13628
rect 11910 13572 11966 13628
rect 11966 13572 11970 13628
rect 11906 13568 11970 13572
rect 11986 13628 12050 13632
rect 11986 13572 11990 13628
rect 11990 13572 12046 13628
rect 12046 13572 12050 13628
rect 11986 13568 12050 13572
rect 3650 13084 3714 13088
rect 3650 13028 3654 13084
rect 3654 13028 3710 13084
rect 3710 13028 3714 13084
rect 3650 13024 3714 13028
rect 3730 13084 3794 13088
rect 3730 13028 3734 13084
rect 3734 13028 3790 13084
rect 3790 13028 3794 13084
rect 3730 13024 3794 13028
rect 3810 13084 3874 13088
rect 3810 13028 3814 13084
rect 3814 13028 3870 13084
rect 3870 13028 3874 13084
rect 3810 13024 3874 13028
rect 3890 13084 3954 13088
rect 3890 13028 3894 13084
rect 3894 13028 3950 13084
rect 3950 13028 3954 13084
rect 3890 13024 3954 13028
rect 9048 13084 9112 13088
rect 9048 13028 9052 13084
rect 9052 13028 9108 13084
rect 9108 13028 9112 13084
rect 9048 13024 9112 13028
rect 9128 13084 9192 13088
rect 9128 13028 9132 13084
rect 9132 13028 9188 13084
rect 9188 13028 9192 13084
rect 9128 13024 9192 13028
rect 9208 13084 9272 13088
rect 9208 13028 9212 13084
rect 9212 13028 9268 13084
rect 9268 13028 9272 13084
rect 9208 13024 9272 13028
rect 9288 13084 9352 13088
rect 9288 13028 9292 13084
rect 9292 13028 9348 13084
rect 9348 13028 9352 13084
rect 9288 13024 9352 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 14605 13084 14669 13088
rect 14605 13028 14609 13084
rect 14609 13028 14665 13084
rect 14665 13028 14669 13084
rect 14605 13024 14669 13028
rect 14685 13084 14749 13088
rect 14685 13028 14689 13084
rect 14689 13028 14745 13084
rect 14745 13028 14749 13084
rect 14685 13024 14749 13028
rect 6349 12540 6413 12544
rect 6349 12484 6353 12540
rect 6353 12484 6409 12540
rect 6409 12484 6413 12540
rect 6349 12480 6413 12484
rect 6429 12540 6493 12544
rect 6429 12484 6433 12540
rect 6433 12484 6489 12540
rect 6489 12484 6493 12540
rect 6429 12480 6493 12484
rect 6509 12540 6573 12544
rect 6509 12484 6513 12540
rect 6513 12484 6569 12540
rect 6569 12484 6573 12540
rect 6509 12480 6573 12484
rect 6589 12540 6653 12544
rect 6589 12484 6593 12540
rect 6593 12484 6649 12540
rect 6649 12484 6653 12540
rect 6589 12480 6653 12484
rect 11746 12540 11810 12544
rect 11746 12484 11750 12540
rect 11750 12484 11806 12540
rect 11806 12484 11810 12540
rect 11746 12480 11810 12484
rect 11826 12540 11890 12544
rect 11826 12484 11830 12540
rect 11830 12484 11886 12540
rect 11886 12484 11890 12540
rect 11826 12480 11890 12484
rect 11906 12540 11970 12544
rect 11906 12484 11910 12540
rect 11910 12484 11966 12540
rect 11966 12484 11970 12540
rect 11906 12480 11970 12484
rect 11986 12540 12050 12544
rect 11986 12484 11990 12540
rect 11990 12484 12046 12540
rect 12046 12484 12050 12540
rect 11986 12480 12050 12484
rect 3650 11996 3714 12000
rect 3650 11940 3654 11996
rect 3654 11940 3710 11996
rect 3710 11940 3714 11996
rect 3650 11936 3714 11940
rect 3730 11996 3794 12000
rect 3730 11940 3734 11996
rect 3734 11940 3790 11996
rect 3790 11940 3794 11996
rect 3730 11936 3794 11940
rect 3810 11996 3874 12000
rect 3810 11940 3814 11996
rect 3814 11940 3870 11996
rect 3870 11940 3874 11996
rect 3810 11936 3874 11940
rect 3890 11996 3954 12000
rect 3890 11940 3894 11996
rect 3894 11940 3950 11996
rect 3950 11940 3954 11996
rect 3890 11936 3954 11940
rect 9048 11996 9112 12000
rect 9048 11940 9052 11996
rect 9052 11940 9108 11996
rect 9108 11940 9112 11996
rect 9048 11936 9112 11940
rect 9128 11996 9192 12000
rect 9128 11940 9132 11996
rect 9132 11940 9188 11996
rect 9188 11940 9192 11996
rect 9128 11936 9192 11940
rect 9208 11996 9272 12000
rect 9208 11940 9212 11996
rect 9212 11940 9268 11996
rect 9268 11940 9272 11996
rect 9208 11936 9272 11940
rect 9288 11996 9352 12000
rect 9288 11940 9292 11996
rect 9292 11940 9348 11996
rect 9348 11940 9352 11996
rect 9288 11936 9352 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 14605 11996 14669 12000
rect 14605 11940 14609 11996
rect 14609 11940 14665 11996
rect 14665 11940 14669 11996
rect 14605 11936 14669 11940
rect 14685 11996 14749 12000
rect 14685 11940 14689 11996
rect 14689 11940 14745 11996
rect 14745 11940 14749 11996
rect 14685 11936 14749 11940
rect 6349 11452 6413 11456
rect 6349 11396 6353 11452
rect 6353 11396 6409 11452
rect 6409 11396 6413 11452
rect 6349 11392 6413 11396
rect 6429 11452 6493 11456
rect 6429 11396 6433 11452
rect 6433 11396 6489 11452
rect 6489 11396 6493 11452
rect 6429 11392 6493 11396
rect 6509 11452 6573 11456
rect 6509 11396 6513 11452
rect 6513 11396 6569 11452
rect 6569 11396 6573 11452
rect 6509 11392 6573 11396
rect 6589 11452 6653 11456
rect 6589 11396 6593 11452
rect 6593 11396 6649 11452
rect 6649 11396 6653 11452
rect 6589 11392 6653 11396
rect 11746 11452 11810 11456
rect 11746 11396 11750 11452
rect 11750 11396 11806 11452
rect 11806 11396 11810 11452
rect 11746 11392 11810 11396
rect 11826 11452 11890 11456
rect 11826 11396 11830 11452
rect 11830 11396 11886 11452
rect 11886 11396 11890 11452
rect 11826 11392 11890 11396
rect 11906 11452 11970 11456
rect 11906 11396 11910 11452
rect 11910 11396 11966 11452
rect 11966 11396 11970 11452
rect 11906 11392 11970 11396
rect 11986 11452 12050 11456
rect 11986 11396 11990 11452
rect 11990 11396 12046 11452
rect 12046 11396 12050 11452
rect 11986 11392 12050 11396
rect 3650 10908 3714 10912
rect 3650 10852 3654 10908
rect 3654 10852 3710 10908
rect 3710 10852 3714 10908
rect 3650 10848 3714 10852
rect 3730 10908 3794 10912
rect 3730 10852 3734 10908
rect 3734 10852 3790 10908
rect 3790 10852 3794 10908
rect 3730 10848 3794 10852
rect 3810 10908 3874 10912
rect 3810 10852 3814 10908
rect 3814 10852 3870 10908
rect 3870 10852 3874 10908
rect 3810 10848 3874 10852
rect 3890 10908 3954 10912
rect 3890 10852 3894 10908
rect 3894 10852 3950 10908
rect 3950 10852 3954 10908
rect 3890 10848 3954 10852
rect 9048 10908 9112 10912
rect 9048 10852 9052 10908
rect 9052 10852 9108 10908
rect 9108 10852 9112 10908
rect 9048 10848 9112 10852
rect 9128 10908 9192 10912
rect 9128 10852 9132 10908
rect 9132 10852 9188 10908
rect 9188 10852 9192 10908
rect 9128 10848 9192 10852
rect 9208 10908 9272 10912
rect 9208 10852 9212 10908
rect 9212 10852 9268 10908
rect 9268 10852 9272 10908
rect 9208 10848 9272 10852
rect 9288 10908 9352 10912
rect 9288 10852 9292 10908
rect 9292 10852 9348 10908
rect 9348 10852 9352 10908
rect 9288 10848 9352 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 14605 10908 14669 10912
rect 14605 10852 14609 10908
rect 14609 10852 14665 10908
rect 14665 10852 14669 10908
rect 14605 10848 14669 10852
rect 14685 10908 14749 10912
rect 14685 10852 14689 10908
rect 14689 10852 14745 10908
rect 14745 10852 14749 10908
rect 14685 10848 14749 10852
rect 6349 10364 6413 10368
rect 6349 10308 6353 10364
rect 6353 10308 6409 10364
rect 6409 10308 6413 10364
rect 6349 10304 6413 10308
rect 6429 10364 6493 10368
rect 6429 10308 6433 10364
rect 6433 10308 6489 10364
rect 6489 10308 6493 10364
rect 6429 10304 6493 10308
rect 6509 10364 6573 10368
rect 6509 10308 6513 10364
rect 6513 10308 6569 10364
rect 6569 10308 6573 10364
rect 6509 10304 6573 10308
rect 6589 10364 6653 10368
rect 6589 10308 6593 10364
rect 6593 10308 6649 10364
rect 6649 10308 6653 10364
rect 6589 10304 6653 10308
rect 11746 10364 11810 10368
rect 11746 10308 11750 10364
rect 11750 10308 11806 10364
rect 11806 10308 11810 10364
rect 11746 10304 11810 10308
rect 11826 10364 11890 10368
rect 11826 10308 11830 10364
rect 11830 10308 11886 10364
rect 11886 10308 11890 10364
rect 11826 10304 11890 10308
rect 11906 10364 11970 10368
rect 11906 10308 11910 10364
rect 11910 10308 11966 10364
rect 11966 10308 11970 10364
rect 11906 10304 11970 10308
rect 11986 10364 12050 10368
rect 11986 10308 11990 10364
rect 11990 10308 12046 10364
rect 12046 10308 12050 10364
rect 11986 10304 12050 10308
rect 3650 9820 3714 9824
rect 3650 9764 3654 9820
rect 3654 9764 3710 9820
rect 3710 9764 3714 9820
rect 3650 9760 3714 9764
rect 3730 9820 3794 9824
rect 3730 9764 3734 9820
rect 3734 9764 3790 9820
rect 3790 9764 3794 9820
rect 3730 9760 3794 9764
rect 3810 9820 3874 9824
rect 3810 9764 3814 9820
rect 3814 9764 3870 9820
rect 3870 9764 3874 9820
rect 3810 9760 3874 9764
rect 3890 9820 3954 9824
rect 3890 9764 3894 9820
rect 3894 9764 3950 9820
rect 3950 9764 3954 9820
rect 3890 9760 3954 9764
rect 9048 9820 9112 9824
rect 9048 9764 9052 9820
rect 9052 9764 9108 9820
rect 9108 9764 9112 9820
rect 9048 9760 9112 9764
rect 9128 9820 9192 9824
rect 9128 9764 9132 9820
rect 9132 9764 9188 9820
rect 9188 9764 9192 9820
rect 9128 9760 9192 9764
rect 9208 9820 9272 9824
rect 9208 9764 9212 9820
rect 9212 9764 9268 9820
rect 9268 9764 9272 9820
rect 9208 9760 9272 9764
rect 9288 9820 9352 9824
rect 9288 9764 9292 9820
rect 9292 9764 9348 9820
rect 9348 9764 9352 9820
rect 9288 9760 9352 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 14605 9820 14669 9824
rect 14605 9764 14609 9820
rect 14609 9764 14665 9820
rect 14665 9764 14669 9820
rect 14605 9760 14669 9764
rect 14685 9820 14749 9824
rect 14685 9764 14689 9820
rect 14689 9764 14745 9820
rect 14745 9764 14749 9820
rect 14685 9760 14749 9764
rect 6349 9276 6413 9280
rect 6349 9220 6353 9276
rect 6353 9220 6409 9276
rect 6409 9220 6413 9276
rect 6349 9216 6413 9220
rect 6429 9276 6493 9280
rect 6429 9220 6433 9276
rect 6433 9220 6489 9276
rect 6489 9220 6493 9276
rect 6429 9216 6493 9220
rect 6509 9276 6573 9280
rect 6509 9220 6513 9276
rect 6513 9220 6569 9276
rect 6569 9220 6573 9276
rect 6509 9216 6573 9220
rect 6589 9276 6653 9280
rect 6589 9220 6593 9276
rect 6593 9220 6649 9276
rect 6649 9220 6653 9276
rect 6589 9216 6653 9220
rect 11746 9276 11810 9280
rect 11746 9220 11750 9276
rect 11750 9220 11806 9276
rect 11806 9220 11810 9276
rect 11746 9216 11810 9220
rect 11826 9276 11890 9280
rect 11826 9220 11830 9276
rect 11830 9220 11886 9276
rect 11886 9220 11890 9276
rect 11826 9216 11890 9220
rect 11906 9276 11970 9280
rect 11906 9220 11910 9276
rect 11910 9220 11966 9276
rect 11966 9220 11970 9276
rect 11906 9216 11970 9220
rect 11986 9276 12050 9280
rect 11986 9220 11990 9276
rect 11990 9220 12046 9276
rect 12046 9220 12050 9276
rect 11986 9216 12050 9220
rect 3650 8732 3714 8736
rect 3650 8676 3654 8732
rect 3654 8676 3710 8732
rect 3710 8676 3714 8732
rect 3650 8672 3714 8676
rect 3730 8732 3794 8736
rect 3730 8676 3734 8732
rect 3734 8676 3790 8732
rect 3790 8676 3794 8732
rect 3730 8672 3794 8676
rect 3810 8732 3874 8736
rect 3810 8676 3814 8732
rect 3814 8676 3870 8732
rect 3870 8676 3874 8732
rect 3810 8672 3874 8676
rect 3890 8732 3954 8736
rect 3890 8676 3894 8732
rect 3894 8676 3950 8732
rect 3950 8676 3954 8732
rect 3890 8672 3954 8676
rect 9048 8732 9112 8736
rect 9048 8676 9052 8732
rect 9052 8676 9108 8732
rect 9108 8676 9112 8732
rect 9048 8672 9112 8676
rect 9128 8732 9192 8736
rect 9128 8676 9132 8732
rect 9132 8676 9188 8732
rect 9188 8676 9192 8732
rect 9128 8672 9192 8676
rect 9208 8732 9272 8736
rect 9208 8676 9212 8732
rect 9212 8676 9268 8732
rect 9268 8676 9272 8732
rect 9208 8672 9272 8676
rect 9288 8732 9352 8736
rect 9288 8676 9292 8732
rect 9292 8676 9348 8732
rect 9348 8676 9352 8732
rect 9288 8672 9352 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 14605 8732 14669 8736
rect 14605 8676 14609 8732
rect 14609 8676 14665 8732
rect 14665 8676 14669 8732
rect 14605 8672 14669 8676
rect 14685 8732 14749 8736
rect 14685 8676 14689 8732
rect 14689 8676 14745 8732
rect 14745 8676 14749 8732
rect 14685 8672 14749 8676
rect 6349 8188 6413 8192
rect 6349 8132 6353 8188
rect 6353 8132 6409 8188
rect 6409 8132 6413 8188
rect 6349 8128 6413 8132
rect 6429 8188 6493 8192
rect 6429 8132 6433 8188
rect 6433 8132 6489 8188
rect 6489 8132 6493 8188
rect 6429 8128 6493 8132
rect 6509 8188 6573 8192
rect 6509 8132 6513 8188
rect 6513 8132 6569 8188
rect 6569 8132 6573 8188
rect 6509 8128 6573 8132
rect 6589 8188 6653 8192
rect 6589 8132 6593 8188
rect 6593 8132 6649 8188
rect 6649 8132 6653 8188
rect 6589 8128 6653 8132
rect 11746 8188 11810 8192
rect 11746 8132 11750 8188
rect 11750 8132 11806 8188
rect 11806 8132 11810 8188
rect 11746 8128 11810 8132
rect 11826 8188 11890 8192
rect 11826 8132 11830 8188
rect 11830 8132 11886 8188
rect 11886 8132 11890 8188
rect 11826 8128 11890 8132
rect 11906 8188 11970 8192
rect 11906 8132 11910 8188
rect 11910 8132 11966 8188
rect 11966 8132 11970 8188
rect 11906 8128 11970 8132
rect 11986 8188 12050 8192
rect 11986 8132 11990 8188
rect 11990 8132 12046 8188
rect 12046 8132 12050 8188
rect 11986 8128 12050 8132
rect 3650 7644 3714 7648
rect 3650 7588 3654 7644
rect 3654 7588 3710 7644
rect 3710 7588 3714 7644
rect 3650 7584 3714 7588
rect 3730 7644 3794 7648
rect 3730 7588 3734 7644
rect 3734 7588 3790 7644
rect 3790 7588 3794 7644
rect 3730 7584 3794 7588
rect 3810 7644 3874 7648
rect 3810 7588 3814 7644
rect 3814 7588 3870 7644
rect 3870 7588 3874 7644
rect 3810 7584 3874 7588
rect 3890 7644 3954 7648
rect 3890 7588 3894 7644
rect 3894 7588 3950 7644
rect 3950 7588 3954 7644
rect 3890 7584 3954 7588
rect 9048 7644 9112 7648
rect 9048 7588 9052 7644
rect 9052 7588 9108 7644
rect 9108 7588 9112 7644
rect 9048 7584 9112 7588
rect 9128 7644 9192 7648
rect 9128 7588 9132 7644
rect 9132 7588 9188 7644
rect 9188 7588 9192 7644
rect 9128 7584 9192 7588
rect 9208 7644 9272 7648
rect 9208 7588 9212 7644
rect 9212 7588 9268 7644
rect 9268 7588 9272 7644
rect 9208 7584 9272 7588
rect 9288 7644 9352 7648
rect 9288 7588 9292 7644
rect 9292 7588 9348 7644
rect 9348 7588 9352 7644
rect 9288 7584 9352 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 14605 7644 14669 7648
rect 14605 7588 14609 7644
rect 14609 7588 14665 7644
rect 14665 7588 14669 7644
rect 14605 7584 14669 7588
rect 14685 7644 14749 7648
rect 14685 7588 14689 7644
rect 14689 7588 14745 7644
rect 14745 7588 14749 7644
rect 14685 7584 14749 7588
rect 6349 7100 6413 7104
rect 6349 7044 6353 7100
rect 6353 7044 6409 7100
rect 6409 7044 6413 7100
rect 6349 7040 6413 7044
rect 6429 7100 6493 7104
rect 6429 7044 6433 7100
rect 6433 7044 6489 7100
rect 6489 7044 6493 7100
rect 6429 7040 6493 7044
rect 6509 7100 6573 7104
rect 6509 7044 6513 7100
rect 6513 7044 6569 7100
rect 6569 7044 6573 7100
rect 6509 7040 6573 7044
rect 6589 7100 6653 7104
rect 6589 7044 6593 7100
rect 6593 7044 6649 7100
rect 6649 7044 6653 7100
rect 6589 7040 6653 7044
rect 11746 7100 11810 7104
rect 11746 7044 11750 7100
rect 11750 7044 11806 7100
rect 11806 7044 11810 7100
rect 11746 7040 11810 7044
rect 11826 7100 11890 7104
rect 11826 7044 11830 7100
rect 11830 7044 11886 7100
rect 11886 7044 11890 7100
rect 11826 7040 11890 7044
rect 11906 7100 11970 7104
rect 11906 7044 11910 7100
rect 11910 7044 11966 7100
rect 11966 7044 11970 7100
rect 11906 7040 11970 7044
rect 11986 7100 12050 7104
rect 11986 7044 11990 7100
rect 11990 7044 12046 7100
rect 12046 7044 12050 7100
rect 11986 7040 12050 7044
rect 3650 6556 3714 6560
rect 3650 6500 3654 6556
rect 3654 6500 3710 6556
rect 3710 6500 3714 6556
rect 3650 6496 3714 6500
rect 3730 6556 3794 6560
rect 3730 6500 3734 6556
rect 3734 6500 3790 6556
rect 3790 6500 3794 6556
rect 3730 6496 3794 6500
rect 3810 6556 3874 6560
rect 3810 6500 3814 6556
rect 3814 6500 3870 6556
rect 3870 6500 3874 6556
rect 3810 6496 3874 6500
rect 3890 6556 3954 6560
rect 3890 6500 3894 6556
rect 3894 6500 3950 6556
rect 3950 6500 3954 6556
rect 3890 6496 3954 6500
rect 9048 6556 9112 6560
rect 9048 6500 9052 6556
rect 9052 6500 9108 6556
rect 9108 6500 9112 6556
rect 9048 6496 9112 6500
rect 9128 6556 9192 6560
rect 9128 6500 9132 6556
rect 9132 6500 9188 6556
rect 9188 6500 9192 6556
rect 9128 6496 9192 6500
rect 9208 6556 9272 6560
rect 9208 6500 9212 6556
rect 9212 6500 9268 6556
rect 9268 6500 9272 6556
rect 9208 6496 9272 6500
rect 9288 6556 9352 6560
rect 9288 6500 9292 6556
rect 9292 6500 9348 6556
rect 9348 6500 9352 6556
rect 9288 6496 9352 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 14605 6556 14669 6560
rect 14605 6500 14609 6556
rect 14609 6500 14665 6556
rect 14665 6500 14669 6556
rect 14605 6496 14669 6500
rect 14685 6556 14749 6560
rect 14685 6500 14689 6556
rect 14689 6500 14745 6556
rect 14745 6500 14749 6556
rect 14685 6496 14749 6500
rect 6349 6012 6413 6016
rect 6349 5956 6353 6012
rect 6353 5956 6409 6012
rect 6409 5956 6413 6012
rect 6349 5952 6413 5956
rect 6429 6012 6493 6016
rect 6429 5956 6433 6012
rect 6433 5956 6489 6012
rect 6489 5956 6493 6012
rect 6429 5952 6493 5956
rect 6509 6012 6573 6016
rect 6509 5956 6513 6012
rect 6513 5956 6569 6012
rect 6569 5956 6573 6012
rect 6509 5952 6573 5956
rect 6589 6012 6653 6016
rect 6589 5956 6593 6012
rect 6593 5956 6649 6012
rect 6649 5956 6653 6012
rect 6589 5952 6653 5956
rect 11746 6012 11810 6016
rect 11746 5956 11750 6012
rect 11750 5956 11806 6012
rect 11806 5956 11810 6012
rect 11746 5952 11810 5956
rect 11826 6012 11890 6016
rect 11826 5956 11830 6012
rect 11830 5956 11886 6012
rect 11886 5956 11890 6012
rect 11826 5952 11890 5956
rect 11906 6012 11970 6016
rect 11906 5956 11910 6012
rect 11910 5956 11966 6012
rect 11966 5956 11970 6012
rect 11906 5952 11970 5956
rect 11986 6012 12050 6016
rect 11986 5956 11990 6012
rect 11990 5956 12046 6012
rect 12046 5956 12050 6012
rect 11986 5952 12050 5956
rect 3650 5468 3714 5472
rect 3650 5412 3654 5468
rect 3654 5412 3710 5468
rect 3710 5412 3714 5468
rect 3650 5408 3714 5412
rect 3730 5468 3794 5472
rect 3730 5412 3734 5468
rect 3734 5412 3790 5468
rect 3790 5412 3794 5468
rect 3730 5408 3794 5412
rect 3810 5468 3874 5472
rect 3810 5412 3814 5468
rect 3814 5412 3870 5468
rect 3870 5412 3874 5468
rect 3810 5408 3874 5412
rect 3890 5468 3954 5472
rect 3890 5412 3894 5468
rect 3894 5412 3950 5468
rect 3950 5412 3954 5468
rect 3890 5408 3954 5412
rect 9048 5468 9112 5472
rect 9048 5412 9052 5468
rect 9052 5412 9108 5468
rect 9108 5412 9112 5468
rect 9048 5408 9112 5412
rect 9128 5468 9192 5472
rect 9128 5412 9132 5468
rect 9132 5412 9188 5468
rect 9188 5412 9192 5468
rect 9128 5408 9192 5412
rect 9208 5468 9272 5472
rect 9208 5412 9212 5468
rect 9212 5412 9268 5468
rect 9268 5412 9272 5468
rect 9208 5408 9272 5412
rect 9288 5468 9352 5472
rect 9288 5412 9292 5468
rect 9292 5412 9348 5468
rect 9348 5412 9352 5468
rect 9288 5408 9352 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 14605 5468 14669 5472
rect 14605 5412 14609 5468
rect 14609 5412 14665 5468
rect 14665 5412 14669 5468
rect 14605 5408 14669 5412
rect 14685 5468 14749 5472
rect 14685 5412 14689 5468
rect 14689 5412 14745 5468
rect 14745 5412 14749 5468
rect 14685 5408 14749 5412
rect 6349 4924 6413 4928
rect 6349 4868 6353 4924
rect 6353 4868 6409 4924
rect 6409 4868 6413 4924
rect 6349 4864 6413 4868
rect 6429 4924 6493 4928
rect 6429 4868 6433 4924
rect 6433 4868 6489 4924
rect 6489 4868 6493 4924
rect 6429 4864 6493 4868
rect 6509 4924 6573 4928
rect 6509 4868 6513 4924
rect 6513 4868 6569 4924
rect 6569 4868 6573 4924
rect 6509 4864 6573 4868
rect 6589 4924 6653 4928
rect 6589 4868 6593 4924
rect 6593 4868 6649 4924
rect 6649 4868 6653 4924
rect 6589 4864 6653 4868
rect 11746 4924 11810 4928
rect 11746 4868 11750 4924
rect 11750 4868 11806 4924
rect 11806 4868 11810 4924
rect 11746 4864 11810 4868
rect 11826 4924 11890 4928
rect 11826 4868 11830 4924
rect 11830 4868 11886 4924
rect 11886 4868 11890 4924
rect 11826 4864 11890 4868
rect 11906 4924 11970 4928
rect 11906 4868 11910 4924
rect 11910 4868 11966 4924
rect 11966 4868 11970 4924
rect 11906 4864 11970 4868
rect 11986 4924 12050 4928
rect 11986 4868 11990 4924
rect 11990 4868 12046 4924
rect 12046 4868 12050 4924
rect 11986 4864 12050 4868
rect 3650 4380 3714 4384
rect 3650 4324 3654 4380
rect 3654 4324 3710 4380
rect 3710 4324 3714 4380
rect 3650 4320 3714 4324
rect 3730 4380 3794 4384
rect 3730 4324 3734 4380
rect 3734 4324 3790 4380
rect 3790 4324 3794 4380
rect 3730 4320 3794 4324
rect 3810 4380 3874 4384
rect 3810 4324 3814 4380
rect 3814 4324 3870 4380
rect 3870 4324 3874 4380
rect 3810 4320 3874 4324
rect 3890 4380 3954 4384
rect 3890 4324 3894 4380
rect 3894 4324 3950 4380
rect 3950 4324 3954 4380
rect 3890 4320 3954 4324
rect 9048 4380 9112 4384
rect 9048 4324 9052 4380
rect 9052 4324 9108 4380
rect 9108 4324 9112 4380
rect 9048 4320 9112 4324
rect 9128 4380 9192 4384
rect 9128 4324 9132 4380
rect 9132 4324 9188 4380
rect 9188 4324 9192 4380
rect 9128 4320 9192 4324
rect 9208 4380 9272 4384
rect 9208 4324 9212 4380
rect 9212 4324 9268 4380
rect 9268 4324 9272 4380
rect 9208 4320 9272 4324
rect 9288 4380 9352 4384
rect 9288 4324 9292 4380
rect 9292 4324 9348 4380
rect 9348 4324 9352 4380
rect 9288 4320 9352 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 14605 4380 14669 4384
rect 14605 4324 14609 4380
rect 14609 4324 14665 4380
rect 14665 4324 14669 4380
rect 14605 4320 14669 4324
rect 14685 4380 14749 4384
rect 14685 4324 14689 4380
rect 14689 4324 14745 4380
rect 14745 4324 14749 4380
rect 14685 4320 14749 4324
rect 6349 3836 6413 3840
rect 6349 3780 6353 3836
rect 6353 3780 6409 3836
rect 6409 3780 6413 3836
rect 6349 3776 6413 3780
rect 6429 3836 6493 3840
rect 6429 3780 6433 3836
rect 6433 3780 6489 3836
rect 6489 3780 6493 3836
rect 6429 3776 6493 3780
rect 6509 3836 6573 3840
rect 6509 3780 6513 3836
rect 6513 3780 6569 3836
rect 6569 3780 6573 3836
rect 6509 3776 6573 3780
rect 6589 3836 6653 3840
rect 6589 3780 6593 3836
rect 6593 3780 6649 3836
rect 6649 3780 6653 3836
rect 6589 3776 6653 3780
rect 11746 3836 11810 3840
rect 11746 3780 11750 3836
rect 11750 3780 11806 3836
rect 11806 3780 11810 3836
rect 11746 3776 11810 3780
rect 11826 3836 11890 3840
rect 11826 3780 11830 3836
rect 11830 3780 11886 3836
rect 11886 3780 11890 3836
rect 11826 3776 11890 3780
rect 11906 3836 11970 3840
rect 11906 3780 11910 3836
rect 11910 3780 11966 3836
rect 11966 3780 11970 3836
rect 11906 3776 11970 3780
rect 11986 3836 12050 3840
rect 11986 3780 11990 3836
rect 11990 3780 12046 3836
rect 12046 3780 12050 3836
rect 11986 3776 12050 3780
rect 3650 3292 3714 3296
rect 3650 3236 3654 3292
rect 3654 3236 3710 3292
rect 3710 3236 3714 3292
rect 3650 3232 3714 3236
rect 3730 3292 3794 3296
rect 3730 3236 3734 3292
rect 3734 3236 3790 3292
rect 3790 3236 3794 3292
rect 3730 3232 3794 3236
rect 3810 3292 3874 3296
rect 3810 3236 3814 3292
rect 3814 3236 3870 3292
rect 3870 3236 3874 3292
rect 3810 3232 3874 3236
rect 3890 3292 3954 3296
rect 3890 3236 3894 3292
rect 3894 3236 3950 3292
rect 3950 3236 3954 3292
rect 3890 3232 3954 3236
rect 9048 3292 9112 3296
rect 9048 3236 9052 3292
rect 9052 3236 9108 3292
rect 9108 3236 9112 3292
rect 9048 3232 9112 3236
rect 9128 3292 9192 3296
rect 9128 3236 9132 3292
rect 9132 3236 9188 3292
rect 9188 3236 9192 3292
rect 9128 3232 9192 3236
rect 9208 3292 9272 3296
rect 9208 3236 9212 3292
rect 9212 3236 9268 3292
rect 9268 3236 9272 3292
rect 9208 3232 9272 3236
rect 9288 3292 9352 3296
rect 9288 3236 9292 3292
rect 9292 3236 9348 3292
rect 9348 3236 9352 3292
rect 9288 3232 9352 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 14605 3292 14669 3296
rect 14605 3236 14609 3292
rect 14609 3236 14665 3292
rect 14665 3236 14669 3292
rect 14605 3232 14669 3236
rect 14685 3292 14749 3296
rect 14685 3236 14689 3292
rect 14689 3236 14745 3292
rect 14745 3236 14749 3292
rect 14685 3232 14749 3236
rect 6349 2748 6413 2752
rect 6349 2692 6353 2748
rect 6353 2692 6409 2748
rect 6409 2692 6413 2748
rect 6349 2688 6413 2692
rect 6429 2748 6493 2752
rect 6429 2692 6433 2748
rect 6433 2692 6489 2748
rect 6489 2692 6493 2748
rect 6429 2688 6493 2692
rect 6509 2748 6573 2752
rect 6509 2692 6513 2748
rect 6513 2692 6569 2748
rect 6569 2692 6573 2748
rect 6509 2688 6573 2692
rect 6589 2748 6653 2752
rect 6589 2692 6593 2748
rect 6593 2692 6649 2748
rect 6649 2692 6653 2748
rect 6589 2688 6653 2692
rect 11746 2748 11810 2752
rect 11746 2692 11750 2748
rect 11750 2692 11806 2748
rect 11806 2692 11810 2748
rect 11746 2688 11810 2692
rect 11826 2748 11890 2752
rect 11826 2692 11830 2748
rect 11830 2692 11886 2748
rect 11886 2692 11890 2748
rect 11826 2688 11890 2692
rect 11906 2748 11970 2752
rect 11906 2692 11910 2748
rect 11910 2692 11966 2748
rect 11966 2692 11970 2748
rect 11906 2688 11970 2692
rect 11986 2748 12050 2752
rect 11986 2692 11990 2748
rect 11990 2692 12046 2748
rect 12046 2692 12050 2748
rect 11986 2688 12050 2692
rect 3650 2204 3714 2208
rect 3650 2148 3654 2204
rect 3654 2148 3710 2204
rect 3710 2148 3714 2204
rect 3650 2144 3714 2148
rect 3730 2204 3794 2208
rect 3730 2148 3734 2204
rect 3734 2148 3790 2204
rect 3790 2148 3794 2204
rect 3730 2144 3794 2148
rect 3810 2204 3874 2208
rect 3810 2148 3814 2204
rect 3814 2148 3870 2204
rect 3870 2148 3874 2204
rect 3810 2144 3874 2148
rect 3890 2204 3954 2208
rect 3890 2148 3894 2204
rect 3894 2148 3950 2204
rect 3950 2148 3954 2204
rect 3890 2144 3954 2148
rect 9048 2204 9112 2208
rect 9048 2148 9052 2204
rect 9052 2148 9108 2204
rect 9108 2148 9112 2204
rect 9048 2144 9112 2148
rect 9128 2204 9192 2208
rect 9128 2148 9132 2204
rect 9132 2148 9188 2204
rect 9188 2148 9192 2204
rect 9128 2144 9192 2148
rect 9208 2204 9272 2208
rect 9208 2148 9212 2204
rect 9212 2148 9268 2204
rect 9268 2148 9272 2204
rect 9208 2144 9272 2148
rect 9288 2204 9352 2208
rect 9288 2148 9292 2204
rect 9292 2148 9348 2204
rect 9348 2148 9352 2204
rect 9288 2144 9352 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
rect 14605 2204 14669 2208
rect 14605 2148 14609 2204
rect 14609 2148 14665 2204
rect 14665 2148 14669 2204
rect 14605 2144 14669 2148
rect 14685 2204 14749 2208
rect 14685 2148 14689 2204
rect 14689 2148 14745 2204
rect 14745 2148 14749 2204
rect 14685 2144 14749 2148
<< metal4 >>
rect 3642 17440 3963 18000
rect 3642 17376 3650 17440
rect 3714 17376 3730 17440
rect 3794 17376 3810 17440
rect 3874 17376 3890 17440
rect 3954 17376 3963 17440
rect 3642 16352 3963 17376
rect 3642 16288 3650 16352
rect 3714 16288 3730 16352
rect 3794 16288 3810 16352
rect 3874 16288 3890 16352
rect 3954 16288 3963 16352
rect 3642 15392 3963 16288
rect 3642 15264 3684 15392
rect 3920 15264 3963 15392
rect 3642 15200 3650 15264
rect 3954 15200 3963 15264
rect 3642 15156 3684 15200
rect 3920 15156 3963 15200
rect 3642 14176 3963 15156
rect 3642 14112 3650 14176
rect 3714 14112 3730 14176
rect 3794 14112 3810 14176
rect 3874 14112 3890 14176
rect 3954 14112 3963 14176
rect 3642 13088 3963 14112
rect 3642 13024 3650 13088
rect 3714 13024 3730 13088
rect 3794 13024 3810 13088
rect 3874 13024 3890 13088
rect 3954 13024 3963 13088
rect 3642 12000 3963 13024
rect 3642 11936 3650 12000
rect 3714 11936 3730 12000
rect 3794 11936 3810 12000
rect 3874 11936 3890 12000
rect 3954 11936 3963 12000
rect 3642 10912 3963 11936
rect 3642 10848 3650 10912
rect 3714 10848 3730 10912
rect 3794 10848 3810 10912
rect 3874 10848 3890 10912
rect 3954 10848 3963 10912
rect 3642 10134 3963 10848
rect 3642 9898 3684 10134
rect 3920 9898 3963 10134
rect 3642 9824 3963 9898
rect 3642 9760 3650 9824
rect 3714 9760 3730 9824
rect 3794 9760 3810 9824
rect 3874 9760 3890 9824
rect 3954 9760 3963 9824
rect 3642 8736 3963 9760
rect 3642 8672 3650 8736
rect 3714 8672 3730 8736
rect 3794 8672 3810 8736
rect 3874 8672 3890 8736
rect 3954 8672 3963 8736
rect 3642 7648 3963 8672
rect 3642 7584 3650 7648
rect 3714 7584 3730 7648
rect 3794 7584 3810 7648
rect 3874 7584 3890 7648
rect 3954 7584 3963 7648
rect 3642 6560 3963 7584
rect 3642 6496 3650 6560
rect 3714 6496 3730 6560
rect 3794 6496 3810 6560
rect 3874 6496 3890 6560
rect 3954 6496 3963 6560
rect 3642 5472 3963 6496
rect 3642 5408 3650 5472
rect 3714 5408 3730 5472
rect 3794 5408 3810 5472
rect 3874 5408 3890 5472
rect 3954 5408 3963 5472
rect 3642 4875 3963 5408
rect 3642 4639 3684 4875
rect 3920 4639 3963 4875
rect 3642 4384 3963 4639
rect 3642 4320 3650 4384
rect 3714 4320 3730 4384
rect 3794 4320 3810 4384
rect 3874 4320 3890 4384
rect 3954 4320 3963 4384
rect 3642 3296 3963 4320
rect 3642 3232 3650 3296
rect 3714 3232 3730 3296
rect 3794 3232 3810 3296
rect 3874 3232 3890 3296
rect 3954 3232 3963 3296
rect 3642 2208 3963 3232
rect 3642 2144 3650 2208
rect 3714 2144 3730 2208
rect 3794 2144 3810 2208
rect 3874 2144 3890 2208
rect 3954 2144 3963 2208
rect 3642 2128 3963 2144
rect 6341 17984 6661 18000
rect 6341 17920 6349 17984
rect 6413 17920 6429 17984
rect 6493 17920 6509 17984
rect 6573 17920 6589 17984
rect 6653 17920 6661 17984
rect 6341 16896 6661 17920
rect 6341 16832 6349 16896
rect 6413 16832 6429 16896
rect 6493 16832 6509 16896
rect 6573 16832 6589 16896
rect 6653 16832 6661 16896
rect 6341 15808 6661 16832
rect 6341 15744 6349 15808
rect 6413 15744 6429 15808
rect 6493 15744 6509 15808
rect 6573 15744 6589 15808
rect 6653 15744 6661 15808
rect 6341 14720 6661 15744
rect 6341 14656 6349 14720
rect 6413 14656 6429 14720
rect 6493 14656 6509 14720
rect 6573 14656 6589 14720
rect 6653 14656 6661 14720
rect 6341 13632 6661 14656
rect 6341 13568 6349 13632
rect 6413 13568 6429 13632
rect 6493 13568 6509 13632
rect 6573 13568 6589 13632
rect 6653 13568 6661 13632
rect 6341 12763 6661 13568
rect 6341 12544 6383 12763
rect 6619 12544 6661 12763
rect 6341 12480 6349 12544
rect 6413 12480 6429 12527
rect 6493 12480 6509 12527
rect 6573 12480 6589 12527
rect 6653 12480 6661 12544
rect 6341 11456 6661 12480
rect 6341 11392 6349 11456
rect 6413 11392 6429 11456
rect 6493 11392 6509 11456
rect 6573 11392 6589 11456
rect 6653 11392 6661 11456
rect 6341 10368 6661 11392
rect 6341 10304 6349 10368
rect 6413 10304 6429 10368
rect 6493 10304 6509 10368
rect 6573 10304 6589 10368
rect 6653 10304 6661 10368
rect 6341 9280 6661 10304
rect 6341 9216 6349 9280
rect 6413 9216 6429 9280
rect 6493 9216 6509 9280
rect 6573 9216 6589 9280
rect 6653 9216 6661 9280
rect 6341 8192 6661 9216
rect 6341 8128 6349 8192
rect 6413 8128 6429 8192
rect 6493 8128 6509 8192
rect 6573 8128 6589 8192
rect 6653 8128 6661 8192
rect 6341 7504 6661 8128
rect 6341 7268 6383 7504
rect 6619 7268 6661 7504
rect 6341 7104 6661 7268
rect 6341 7040 6349 7104
rect 6413 7040 6429 7104
rect 6493 7040 6509 7104
rect 6573 7040 6589 7104
rect 6653 7040 6661 7104
rect 6341 6016 6661 7040
rect 6341 5952 6349 6016
rect 6413 5952 6429 6016
rect 6493 5952 6509 6016
rect 6573 5952 6589 6016
rect 6653 5952 6661 6016
rect 6341 4928 6661 5952
rect 6341 4864 6349 4928
rect 6413 4864 6429 4928
rect 6493 4864 6509 4928
rect 6573 4864 6589 4928
rect 6653 4864 6661 4928
rect 6341 3840 6661 4864
rect 6341 3776 6349 3840
rect 6413 3776 6429 3840
rect 6493 3776 6509 3840
rect 6573 3776 6589 3840
rect 6653 3776 6661 3840
rect 6341 2752 6661 3776
rect 6341 2688 6349 2752
rect 6413 2688 6429 2752
rect 6493 2688 6509 2752
rect 6573 2688 6589 2752
rect 6653 2688 6661 2752
rect 6341 2128 6661 2688
rect 9040 17440 9360 18000
rect 9040 17376 9048 17440
rect 9112 17376 9128 17440
rect 9192 17376 9208 17440
rect 9272 17376 9288 17440
rect 9352 17376 9360 17440
rect 9040 16352 9360 17376
rect 9040 16288 9048 16352
rect 9112 16288 9128 16352
rect 9192 16288 9208 16352
rect 9272 16288 9288 16352
rect 9352 16288 9360 16352
rect 9040 15392 9360 16288
rect 9040 15264 9082 15392
rect 9318 15264 9360 15392
rect 9040 15200 9048 15264
rect 9352 15200 9360 15264
rect 9040 15156 9082 15200
rect 9318 15156 9360 15200
rect 9040 14176 9360 15156
rect 9040 14112 9048 14176
rect 9112 14112 9128 14176
rect 9192 14112 9208 14176
rect 9272 14112 9288 14176
rect 9352 14112 9360 14176
rect 9040 13088 9360 14112
rect 9040 13024 9048 13088
rect 9112 13024 9128 13088
rect 9192 13024 9208 13088
rect 9272 13024 9288 13088
rect 9352 13024 9360 13088
rect 9040 12000 9360 13024
rect 9040 11936 9048 12000
rect 9112 11936 9128 12000
rect 9192 11936 9208 12000
rect 9272 11936 9288 12000
rect 9352 11936 9360 12000
rect 9040 10912 9360 11936
rect 9040 10848 9048 10912
rect 9112 10848 9128 10912
rect 9192 10848 9208 10912
rect 9272 10848 9288 10912
rect 9352 10848 9360 10912
rect 9040 10134 9360 10848
rect 9040 9898 9082 10134
rect 9318 9898 9360 10134
rect 9040 9824 9360 9898
rect 9040 9760 9048 9824
rect 9112 9760 9128 9824
rect 9192 9760 9208 9824
rect 9272 9760 9288 9824
rect 9352 9760 9360 9824
rect 9040 8736 9360 9760
rect 9040 8672 9048 8736
rect 9112 8672 9128 8736
rect 9192 8672 9208 8736
rect 9272 8672 9288 8736
rect 9352 8672 9360 8736
rect 9040 7648 9360 8672
rect 9040 7584 9048 7648
rect 9112 7584 9128 7648
rect 9192 7584 9208 7648
rect 9272 7584 9288 7648
rect 9352 7584 9360 7648
rect 9040 6560 9360 7584
rect 9040 6496 9048 6560
rect 9112 6496 9128 6560
rect 9192 6496 9208 6560
rect 9272 6496 9288 6560
rect 9352 6496 9360 6560
rect 9040 5472 9360 6496
rect 9040 5408 9048 5472
rect 9112 5408 9128 5472
rect 9192 5408 9208 5472
rect 9272 5408 9288 5472
rect 9352 5408 9360 5472
rect 9040 4875 9360 5408
rect 9040 4639 9082 4875
rect 9318 4639 9360 4875
rect 9040 4384 9360 4639
rect 9040 4320 9048 4384
rect 9112 4320 9128 4384
rect 9192 4320 9208 4384
rect 9272 4320 9288 4384
rect 9352 4320 9360 4384
rect 9040 3296 9360 4320
rect 9040 3232 9048 3296
rect 9112 3232 9128 3296
rect 9192 3232 9208 3296
rect 9272 3232 9288 3296
rect 9352 3232 9360 3296
rect 9040 2208 9360 3232
rect 9040 2144 9048 2208
rect 9112 2144 9128 2208
rect 9192 2144 9208 2208
rect 9272 2144 9288 2208
rect 9352 2144 9360 2208
rect 9040 2128 9360 2144
rect 11738 17984 12059 18000
rect 11738 17920 11746 17984
rect 11810 17920 11826 17984
rect 11890 17920 11906 17984
rect 11970 17920 11986 17984
rect 12050 17920 12059 17984
rect 11738 16896 12059 17920
rect 11738 16832 11746 16896
rect 11810 16832 11826 16896
rect 11890 16832 11906 16896
rect 11970 16832 11986 16896
rect 12050 16832 12059 16896
rect 11738 15808 12059 16832
rect 11738 15744 11746 15808
rect 11810 15744 11826 15808
rect 11890 15744 11906 15808
rect 11970 15744 11986 15808
rect 12050 15744 12059 15808
rect 11738 14720 12059 15744
rect 11738 14656 11746 14720
rect 11810 14656 11826 14720
rect 11890 14656 11906 14720
rect 11970 14656 11986 14720
rect 12050 14656 12059 14720
rect 11738 13632 12059 14656
rect 11738 13568 11746 13632
rect 11810 13568 11826 13632
rect 11890 13568 11906 13632
rect 11970 13568 11986 13632
rect 12050 13568 12059 13632
rect 11738 12763 12059 13568
rect 11738 12544 11780 12763
rect 12016 12544 12059 12763
rect 11738 12480 11746 12544
rect 11810 12480 11826 12527
rect 11890 12480 11906 12527
rect 11970 12480 11986 12527
rect 12050 12480 12059 12544
rect 11738 11456 12059 12480
rect 11738 11392 11746 11456
rect 11810 11392 11826 11456
rect 11890 11392 11906 11456
rect 11970 11392 11986 11456
rect 12050 11392 12059 11456
rect 11738 10368 12059 11392
rect 11738 10304 11746 10368
rect 11810 10304 11826 10368
rect 11890 10304 11906 10368
rect 11970 10304 11986 10368
rect 12050 10304 12059 10368
rect 11738 9280 12059 10304
rect 11738 9216 11746 9280
rect 11810 9216 11826 9280
rect 11890 9216 11906 9280
rect 11970 9216 11986 9280
rect 12050 9216 12059 9280
rect 11738 8192 12059 9216
rect 11738 8128 11746 8192
rect 11810 8128 11826 8192
rect 11890 8128 11906 8192
rect 11970 8128 11986 8192
rect 12050 8128 12059 8192
rect 11738 7504 12059 8128
rect 11738 7268 11780 7504
rect 12016 7268 12059 7504
rect 11738 7104 12059 7268
rect 11738 7040 11746 7104
rect 11810 7040 11826 7104
rect 11890 7040 11906 7104
rect 11970 7040 11986 7104
rect 12050 7040 12059 7104
rect 11738 6016 12059 7040
rect 11738 5952 11746 6016
rect 11810 5952 11826 6016
rect 11890 5952 11906 6016
rect 11970 5952 11986 6016
rect 12050 5952 12059 6016
rect 11738 4928 12059 5952
rect 11738 4864 11746 4928
rect 11810 4864 11826 4928
rect 11890 4864 11906 4928
rect 11970 4864 11986 4928
rect 12050 4864 12059 4928
rect 11738 3840 12059 4864
rect 11738 3776 11746 3840
rect 11810 3776 11826 3840
rect 11890 3776 11906 3840
rect 11970 3776 11986 3840
rect 12050 3776 12059 3840
rect 11738 2752 12059 3776
rect 11738 2688 11746 2752
rect 11810 2688 11826 2752
rect 11890 2688 11906 2752
rect 11970 2688 11986 2752
rect 12050 2688 12059 2752
rect 11738 2128 12059 2688
rect 14437 17440 14757 18000
rect 14437 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14605 17440
rect 14669 17376 14685 17440
rect 14749 17376 14757 17440
rect 14437 16352 14757 17376
rect 14437 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14605 16352
rect 14669 16288 14685 16352
rect 14749 16288 14757 16352
rect 14437 15392 14757 16288
rect 14437 15264 14479 15392
rect 14715 15264 14757 15392
rect 14437 15200 14445 15264
rect 14749 15200 14757 15264
rect 14437 15156 14479 15200
rect 14715 15156 14757 15200
rect 14437 14176 14757 15156
rect 14437 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14605 14176
rect 14669 14112 14685 14176
rect 14749 14112 14757 14176
rect 14437 13088 14757 14112
rect 14437 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14605 13088
rect 14669 13024 14685 13088
rect 14749 13024 14757 13088
rect 14437 12000 14757 13024
rect 14437 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14605 12000
rect 14669 11936 14685 12000
rect 14749 11936 14757 12000
rect 14437 10912 14757 11936
rect 14437 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14605 10912
rect 14669 10848 14685 10912
rect 14749 10848 14757 10912
rect 14437 10134 14757 10848
rect 14437 9898 14479 10134
rect 14715 9898 14757 10134
rect 14437 9824 14757 9898
rect 14437 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14605 9824
rect 14669 9760 14685 9824
rect 14749 9760 14757 9824
rect 14437 8736 14757 9760
rect 14437 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14605 8736
rect 14669 8672 14685 8736
rect 14749 8672 14757 8736
rect 14437 7648 14757 8672
rect 14437 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14605 7648
rect 14669 7584 14685 7648
rect 14749 7584 14757 7648
rect 14437 6560 14757 7584
rect 14437 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14605 6560
rect 14669 6496 14685 6560
rect 14749 6496 14757 6560
rect 14437 5472 14757 6496
rect 14437 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14605 5472
rect 14669 5408 14685 5472
rect 14749 5408 14757 5472
rect 14437 4875 14757 5408
rect 14437 4639 14479 4875
rect 14715 4639 14757 4875
rect 14437 4384 14757 4639
rect 14437 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14605 4384
rect 14669 4320 14685 4384
rect 14749 4320 14757 4384
rect 14437 3296 14757 4320
rect 14437 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14605 3296
rect 14669 3232 14685 3296
rect 14749 3232 14757 3296
rect 14437 2208 14757 3232
rect 14437 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14605 2208
rect 14669 2144 14685 2208
rect 14749 2144 14757 2208
rect 14437 2128 14757 2144
<< via4 >>
rect 3684 15264 3920 15392
rect 3684 15200 3714 15264
rect 3714 15200 3730 15264
rect 3730 15200 3794 15264
rect 3794 15200 3810 15264
rect 3810 15200 3874 15264
rect 3874 15200 3890 15264
rect 3890 15200 3920 15264
rect 3684 15156 3920 15200
rect 3684 9898 3920 10134
rect 3684 4639 3920 4875
rect 6383 12544 6619 12763
rect 6383 12527 6413 12544
rect 6413 12527 6429 12544
rect 6429 12527 6493 12544
rect 6493 12527 6509 12544
rect 6509 12527 6573 12544
rect 6573 12527 6589 12544
rect 6589 12527 6619 12544
rect 6383 7268 6619 7504
rect 9082 15264 9318 15392
rect 9082 15200 9112 15264
rect 9112 15200 9128 15264
rect 9128 15200 9192 15264
rect 9192 15200 9208 15264
rect 9208 15200 9272 15264
rect 9272 15200 9288 15264
rect 9288 15200 9318 15264
rect 9082 15156 9318 15200
rect 9082 9898 9318 10134
rect 9082 4639 9318 4875
rect 11780 12544 12016 12763
rect 11780 12527 11810 12544
rect 11810 12527 11826 12544
rect 11826 12527 11890 12544
rect 11890 12527 11906 12544
rect 11906 12527 11970 12544
rect 11970 12527 11986 12544
rect 11986 12527 12016 12544
rect 11780 7268 12016 7504
rect 14479 15264 14715 15392
rect 14479 15200 14509 15264
rect 14509 15200 14525 15264
rect 14525 15200 14589 15264
rect 14589 15200 14605 15264
rect 14605 15200 14669 15264
rect 14669 15200 14685 15264
rect 14685 15200 14715 15264
rect 14479 15156 14715 15200
rect 14479 9898 14715 10134
rect 14479 4639 14715 4875
<< metal5 >>
rect 1104 15392 17296 15435
rect 1104 15156 3684 15392
rect 3920 15156 9082 15392
rect 9318 15156 14479 15392
rect 14715 15156 17296 15392
rect 1104 15114 17296 15156
rect 1104 12763 17296 12805
rect 1104 12527 6383 12763
rect 6619 12527 11780 12763
rect 12016 12527 17296 12763
rect 1104 12485 17296 12527
rect 1104 10134 17296 10176
rect 1104 9898 3684 10134
rect 3920 9898 9082 10134
rect 9318 9898 14479 10134
rect 14715 9898 17296 10134
rect 1104 9856 17296 9898
rect 1104 7504 17296 7547
rect 1104 7268 6383 7504
rect 6619 7268 11780 7504
rect 12016 7268 17296 7504
rect 1104 7226 17296 7268
rect 1104 4875 17296 4917
rect 1104 4639 3684 4875
rect 3920 4639 9082 4875
rect 9318 4639 14479 4875
rect 14715 4639 17296 4875
rect 1104 4597 17296 4639
use sky130_fd_sc_hd__decap_3  FILLER_1_9
timestamp 1619617919
transform 1 0 1932 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output45
timestamp 1619617919
transform -1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1619617919
transform 1 0 2024 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1619617919
transform -1 0 1656 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1619617919
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1619617919
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ringosc.ibufp11
timestamp 1619617919
transform -1 0 1932 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  ringosc.ibufp10
timestamp 1619617919
transform -1 0 2484 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1619617919
transform 1 0 1748 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21
timestamp 1619617919
transform 1 0 3036 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17
timestamp 1619617919
transform 1 0 2668 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1619617919
transform 1 0 2300 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1619617919
transform -1 0 3036 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfrbp_2  idiv2
timestamp 1619617919
transform 1 0 2484 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_4  irb
timestamp 1619617919
transform -1 0 5244 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1619617919
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1619617919
transform -1 0 4416 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1619617919
transform -1 0 5796 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30
timestamp 1619617919
transform 1 0 3864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36
timestamp 1619617919
transform 1 0 4416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45
timestamp 1619617919
transform 1 0 5244 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1619617919
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_51
timestamp 1619617919
transform 1 0 5796 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1619617919
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1619617919
transform 1 0 6348 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51
timestamp 1619617919
transform 1 0 5796 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1619617919
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1619617919
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_4  ringosc.dstage\[11\].id.delayen0
timestamp 1619617919
transform 1 0 6440 0 1 2720
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69
timestamp 1619617919
transform 1 0 7452 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1619617919
transform -1 0 7176 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1619617919
transform -1 0 7452 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[11\].id.delayenb1
timestamp 1619617919
transform -1 0 8096 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_0_82
timestamp 1619617919
transform 1 0 8648 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77
timestamp 1619617919
transform 1 0 8188 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1619617919
transform 1 0 8280 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1619617919
transform 1 0 8096 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1619617919
transform 1 0 8372 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1619617919
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1619617919
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86
timestamp 1619617919
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1619617919
transform 1 0 9660 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1619617919
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp 1619617919
transform -1 0 10028 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96
timestamp 1619617919
transform 1 0 9936 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb1
timestamp 1619617919
transform 1 0 10028 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_1_104
timestamp 1619617919
transform 1 0 10672 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_106
timestamp 1619617919
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102
timestamp 1619617919
transform 1 0 10488 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1619617919
transform 1 0 11040 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1619617919
transform 1 0 10580 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1619617919
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_1_115
timestamp 1619617919
transform 1 0 11684 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117
timestamp 1619617919
transform 1 0 11868 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115
timestamp 1619617919
transform 1 0 11684 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111
timestamp 1619617919
transform 1 0 11316 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1619617919
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1619617919
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  input1
timestamp 1619617919
transform 1 0 12420 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1619617919
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1619617919
transform -1 0 14352 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _324_
timestamp 1619617919
transform -1 0 13984 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1619617919
transform 1 0 14536 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1619617919
transform 1 0 13248 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1619617919
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1619617919
transform -1 0 14352 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output43
timestamp 1619617919
transform 1 0 14536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144
timestamp 1619617919
transform 1 0 14352 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1619617919
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_158
timestamp 1619617919
transform 1 0 15640 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1619617919
transform 1 0 15364 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_172
timestamp 1619617919
transform 1 0 16928 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_164
timestamp 1619617919
transform 1 0 16192 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1619617919
transform 1 0 16284 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1619617919
transform 1 0 16560 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1619617919
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1619617919
transform -1 0 17296 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1619617919
transform -1 0 17296 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfrbp_1  idiv16
timestamp 1619617919
transform -1 0 17020 0 -1 2720
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1619617919
transform 1 0 3220 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1619617919
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1619617919
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_15
timestamp 1619617919
transform 1 0 2484 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfrbp_2  idiv4
timestamp 1619617919
transform -1 0 6072 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1619617919
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1619617919
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[11\].id.delayen1
timestamp 1619617919
transform -1 0 7820 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb0
timestamp 1619617919
transform 1 0 6072 0 -1 3808
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  FILLER_2_65
timestamp 1619617919
transform 1 0 7084 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_73
timestamp 1619617919
transform 1 0 7820 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1619617919
transform -1 0 8740 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1619617919
transform 1 0 9936 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen1
timestamp 1619617919
transform 1 0 9384 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1619617919
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_83
timestamp 1619617919
transform 1 0 8740 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_87
timestamp 1619617919
transform 1 0 9108 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_95
timestamp 1619617919
transform 1 0 9844 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_99
timestamp 1619617919
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen0
timestamp 1619617919
transform -1 0 11500 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb0
timestamp 1619617919
transform -1 0 11040 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_2_113
timestamp 1619617919
transform 1 0 11500 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1619617919
transform 1 0 13616 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _322_
timestamp 1619617919
transform -1 0 13616 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfrbp_2  idiv8
timestamp 1619617919
transform 1 0 14720 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1619617919
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_125
timestamp 1619617919
transform 1 0 12604 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_139
timestamp 1619617919
transform 1 0 13892 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_144
timestamp 1619617919
transform 1 0 14352 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1619617919
transform -1 0 17296 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_172
timestamp 1619617919
transform 1 0 16928 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1619617919
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output41
timestamp 1619617919
transform -1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_7
timestamp 1619617919
transform 1 0 1748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_19
timestamp 1619617919
transform 1 0 2852 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01
timestamp 1619617919
transform 1 0 3680 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_3_27
timestamp 1619617919
transform 1 0 3588 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_41
timestamp 1619617919
transform 1 0 4876 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1619617919
transform 1 0 7084 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.delayen1
timestamp 1619617919
transform 1 0 6624 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1619617919
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_53
timestamp 1619617919
transform 1 0 5980 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_58
timestamp 1619617919
transform 1 0 6440 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_68
timestamp 1619617919
transform 1 0 7360 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_80
timestamp 1619617919
transform 1 0 8464 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_92
timestamp 1619617919
transform 1 0 9568 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1619617919
transform 1 0 12052 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1619617919
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1619617919
transform 1 0 10672 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_112
timestamp 1619617919
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1619617919
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _323_
timestamp 1619617919
transform -1 0 13800 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _325_
timestamp 1619617919
transform 1 0 13800 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_128
timestamp 1619617919
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_146
timestamp 1619617919
transform 1 0 14536 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1619617919
transform -1 0 17296 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1619617919
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_158
timestamp 1619617919
transform 1 0 15640 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_170
timestamp 1619617919
transform 1 0 16744 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_172
timestamp 1619617919
transform 1 0 16928 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen0
timestamp 1619617919
transform 1 0 2392 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb0
timestamp 1619617919
transform 1 0 1748 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1619617919
transform 1 0 2852 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1619617919
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1619617919
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_22
timestamp 1619617919
transform 1 0 3128 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00
timestamp 1619617919
transform -1 0 4416 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0
timestamp 1619617919
transform -1 0 4876 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb0
timestamp 1619617919
transform 1 0 4876 0 -1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1619617919
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_28
timestamp 1619617919
transform 1 0 3680 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_30
timestamp 1619617919
transform 1 0 3864 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.delayen0
timestamp 1619617919
transform 1 0 5980 0 -1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_2  ringosc.iss.delayenb1
timestamp 1619617919
transform 1 0 6992 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1619617919
transform 1 0 7636 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_52
timestamp 1619617919
transform 1 0 5888 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_74
timestamp 1619617919
transform 1 0 7912 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen0
timestamp 1619617919
transform 1 0 9108 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb0
timestamp 1619617919
transform 1 0 8188 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1619617919
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1619617919
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_92
timestamp 1619617919
transform 1 0 9568 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1619617919
transform -1 0 11224 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_104
timestamp 1619617919
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_110
timestamp 1619617919
transform 1 0 11224 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_122
timestamp 1619617919
transform 1 0 12328 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp 1619617919
transform -1 0 15364 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1619617919
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_134
timestamp 1619617919
transform 1 0 13432 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_142
timestamp 1619617919
transform 1 0 14168 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_144
timestamp 1619617919
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1619617919
transform -1 0 17296 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1619617919
transform -1 0 17020 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_155
timestamp 1619617919
transform 1 0 15364 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_167
timestamp 1619617919
transform 1 0 16468 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1619617919
transform 1 0 2852 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen1
timestamp 1619617919
transform 1 0 2392 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb1
timestamp 1619617919
transform 1 0 1748 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1619617919
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1619617919
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_22
timestamp 1619617919
transform 1 0 3128 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1
timestamp 1619617919
transform 1 0 5428 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.reseten0
timestamp 1619617919
transform 1 0 4416 0 1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_5_34
timestamp 1619617919
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _356_
timestamp 1619617919
transform -1 0 8648 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1619617919
transform 1 0 6440 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1619617919
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp 1619617919
transform 1 0 5704 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_56
timestamp 1619617919
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_67
timestamp 1619617919
transform 1 0 7268 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _377_
timestamp 1619617919
transform -1 0 9844 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb1
timestamp 1619617919
transform -1 0 10672 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_5_82
timestamp 1619617919
transform 1 0 8648 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_95
timestamp 1619617919
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0
timestamp 1619617919
transform 1 0 12328 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb1
timestamp 1619617919
transform 1 0 11684 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1619617919
transform 1 0 11132 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen1
timestamp 1619617919
transform 1 0 10672 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1619617919
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_112
timestamp 1619617919
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen0
timestamp 1619617919
transform 1 0 13340 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb0
timestamp 1619617919
transform -1 0 13340 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 1619617919
transform 1 0 13800 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1619617919
transform 1 0 14444 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb1
timestamp 1619617919
transform -1 0 15456 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_5_141
timestamp 1619617919
transform 1 0 14076 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1619617919
transform 1 0 15916 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen1
timestamp 1619617919
transform 1 0 15456 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1619617919
transform -1 0 17296 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1619617919
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_164
timestamp 1619617919
transform 1 0 16192 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_170
timestamp 1619617919
transform 1 0 16744 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_172
timestamp 1619617919
transform 1 0 16928 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _360_
timestamp 1619617919
transform -1 0 2392 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb0
timestamp 1619617919
transform -1 0 3956 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1619617919
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1619617919
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1619617919
transform -1 0 1656 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_6
timestamp 1619617919
transform 1 0 1656 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_18
timestamp 1619617919
transform 1 0 2760 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1619617919
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_14
timestamp 1619617919
transform 1 0 2392 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _196_
timestamp 1619617919
transform -1 0 4876 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _303_
timestamp 1619617919
transform 1 0 5520 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1619617919
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_26
timestamp 1619617919
transform 1 0 3496 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_30
timestamp 1619617919
transform 1 0 3864 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1619617919
transform 1 0 4876 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_31
timestamp 1619617919
transform 1 0 3956 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_43
timestamp 1619617919
transform 1 0 5060 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_47
timestamp 1619617919
transform 1 0 5428 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _306_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 7912 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1619617919
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1619617919
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1619617919
transform 1 0 5980 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1619617919
transform 1 0 7084 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_54
timestamp 1619617919
transform 1 0 6072 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_58
timestamp 1619617919
transform 1 0 6440 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_71
timestamp 1619617919
transform 1 0 7636 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1619617919
transform -1 0 10304 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1619617919
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_77
timestamp 1619617919
transform 1 0 8188 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1619617919
transform 1 0 8924 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_87
timestamp 1619617919
transform 1 0 9108 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_95
timestamp 1619617919
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1619617919
transform 1 0 8464 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_92
timestamp 1619617919
transform 1 0 9568 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_110
timestamp 1619617919
transform 1 0 11224 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1619617919
transform 1 0 10948 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1619617919
transform -1 0 10948 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_120
timestamp 1619617919
transform 1 0 12144 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_112
timestamp 1619617919
transform 1 0 11408 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1619617919
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen1
timestamp 1619617919
transform 1 0 11684 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1619617919
transform 1 0 12236 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_115
timestamp 1619617919
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_124
timestamp 1619617919
transform 1 0 12512 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_100
timestamp 1619617919
transform 1 0 10304 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb0
timestamp 1619617919
transform 1 0 14812 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1619617919
transform -1 0 13708 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1619617919
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_136
timestamp 1619617919
transform 1 0 13616 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_142
timestamp 1619617919
transform 1 0 14168 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_144
timestamp 1619617919
transform 1 0 14352 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_127
timestamp 1619617919
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1619617919
transform 1 0 13708 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_156
timestamp 1619617919
transform 1 0 15456 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen0
timestamp 1619617919
transform 1 0 15456 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_7_161
timestamp 1619617919
transform 1 0 15916 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_162
timestamp 1619617919
transform 1 0 16008 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1619617919
transform 1 0 15732 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_172
timestamp 1619617919
transform 1 0 16928 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1619617919
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_170
timestamp 1619617919
transform 1 0 16744 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1619617919
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1619617919
transform -1 0 17296 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1619617919
transform -1 0 17296 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1619617919
transform -1 0 2392 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1619617919
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1619617919
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_14
timestamp 1619617919
transform 1 0 2392 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _314_
timestamp 1619617919
transform 1 0 5428 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1619617919
transform 1 0 5152 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1619617919
transform 1 0 3864 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[5\].id.delayenb1
timestamp 1619617919
transform 1 0 4508 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1619617919
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_26
timestamp 1619617919
transform 1 0 3496 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _321_
timestamp 1619617919
transform 1 0 7268 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _369_
timestamp 1619617919
transform -1 0 8740 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1619617919
transform 1 0 5980 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_65
timestamp 1619617919
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_73
timestamp 1619617919
transform 1 0 7820 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _312_
timestamp 1619617919
transform -1 0 9660 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb1
timestamp 1619617919
transform 1 0 9844 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1619617919
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_83
timestamp 1619617919
transform 1 0 8740 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1619617919
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_2  _368_
timestamp 1619617919
transform 1 0 12144 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen1
timestamp 1619617919
transform 1 0 10488 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[4\].id.delayenb0
timestamp 1619617919
transform -1 0 12144 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_8_107
timestamp 1619617919
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1619617919
transform 1 0 13248 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1619617919
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_129
timestamp 1619617919
transform 1 0 12972 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1619617919
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1619617919
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1619617919
transform 1 0 16192 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1619617919
transform -1 0 17296 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1619617919
transform 1 0 16744 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_156
timestamp 1619617919
transform 1 0 15456 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_168
timestamp 1619617919
transform 1 0 16560 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1619617919
transform -1 0 2760 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1619617919
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1619617919
transform 1 0 1380 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_11
timestamp 1619617919
transform 1 0 2116 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_18
timestamp 1619617919
transform 1 0 2760 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1619617919
transform -1 0 5336 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[5\].id.delayen1
timestamp 1619617919
transform 1 0 3864 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1619617919
transform 1 0 4324 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_38
timestamp 1619617919
transform 1 0 4600 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_46
timestamp 1619617919
transform 1 0 5336 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1619617919
transform -1 0 8096 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _354_
timestamp 1619617919
transform 1 0 6440 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1619617919
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_54
timestamp 1619617919
transform 1 0 6072 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_67
timestamp 1619617919
transform 1 0 7268 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _315_
timestamp 1619617919
transform 1 0 8740 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _319_
timestamp 1619617919
transform -1 0 8648 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _374_
timestamp 1619617919
transform -1 0 10488 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_82
timestamp 1619617919
transform 1 0 8648 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_88
timestamp 1619617919
transform 1 0 9200 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_92
timestamp 1619617919
transform 1 0 9568 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _291_
timestamp 1619617919
transform 1 0 12420 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1619617919
transform -1 0 11500 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1619617919
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_102
timestamp 1619617919
transform 1 0 10488 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1619617919
transform 1 0 11500 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_115
timestamp 1619617919
transform 1 0 11684 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen0
timestamp 1619617919
transform 1 0 13800 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb0
timestamp 1619617919
transform 1 0 13156 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_9_128
timestamp 1619617919
transform 1 0 12880 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_143
timestamp 1619617919
transform 1 0 14260 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1619617919
transform -1 0 17296 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1619617919
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_155
timestamp 1619617919
transform 1 0 15364 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_167
timestamp 1619617919
transform 1 0 16468 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_172
timestamp 1619617919
transform 1 0 16928 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb0
timestamp 1619617919
transform 1 0 1380 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1619617919
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_10
timestamp 1619617919
transform 1 0 2024 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_22
timestamp 1619617919
transform 1 0 3128 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _372_
timestamp 1619617919
transform -1 0 6440 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1619617919
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_28
timestamp 1619617919
transform 1 0 3680 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1619617919
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_42
timestamp 1619617919
transform 1 0 4968 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_48
timestamp 1619617919
transform 1 0 5520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1619617919
transform -1 0 8004 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _302_
timestamp 1619617919
transform 1 0 7268 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _307_
timestamp 1619617919
transform 1 0 6440 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_10_65
timestamp 1619617919
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_71
timestamp 1619617919
transform 1 0 7636 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1619617919
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  repeater46
timestamp 1619617919
transform -1 0 10212 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_75
timestamp 1619617919
transform 1 0 8004 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_83
timestamp 1619617919
transform 1 0 8740 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_99
timestamp 1619617919
transform 1 0 10212 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_111
timestamp 1619617919
transform 1 0 11316 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1619617919
transform 1 0 12420 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1619617919
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_135
timestamp 1619617919
transform 1 0 13524 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_144
timestamp 1619617919
transform 1 0 14352 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen0
timestamp 1619617919
transform -1 0 16376 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb0
timestamp 1619617919
transform 1 0 15272 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1619617919
transform -1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1619617919
transform -1 0 17296 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_166
timestamp 1619617919
transform 1 0 16376 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_172
timestamp 1619617919
transform 1 0 16928 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen0
timestamp 1619617919
transform 1 0 1840 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen1
timestamp 1619617919
transform 1 0 3220 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb1
timestamp 1619617919
transform -1 0 3220 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1619617919
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output39
timestamp 1619617919
transform -1 0 1748 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1619617919
transform 1 0 1748 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_13
timestamp 1619617919
transform 1 0 2300 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _304_
timestamp 1619617919
transform 1 0 5336 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1619617919
transform 1 0 4140 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1619617919
transform 1 0 3680 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_31
timestamp 1619617919
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_42
timestamp 1619617919
transform 1 0 4968 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _296_
timestamp 1619617919
transform -1 0 6900 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1619617919
transform 1 0 6900 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _298_
timestamp 1619617919
transform -1 0 8004 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _300_
timestamp 1619617919
transform 1 0 5980 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1619617919
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_66
timestamp 1619617919
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _301_
timestamp 1619617919
transform 1 0 8004 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _308_
timestamp 1619617919
transform 1 0 9200 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_11_79
timestamp 1619617919
transform 1 0 8372 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_87
timestamp 1619617919
transform 1 0 9108 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_95
timestamp 1619617919
transform 1 0 9844 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1619617919
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _365_
timestamp 1619617919
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1619617919
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_103
timestamp 1619617919
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_115
timestamp 1619617919
transform 1 0 11684 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _347_
timestamp 1619617919
transform 1 0 13248 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1619617919
transform 1 0 13892 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_135
timestamp 1619617919
transform 1 0 13524 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_142
timestamp 1619617919
transform 1 0 14168 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1619617919
transform -1 0 16192 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1619617919
transform -1 0 17296 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1619617919
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_154
timestamp 1619617919
transform 1 0 15272 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_160
timestamp 1619617919
transform 1 0 15824 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_164
timestamp 1619617919
transform 1 0 16192 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_170
timestamp 1619617919
transform 1 0 16744 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_172
timestamp 1619617919
transform 1 0 16928 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1619617919
transform -1 0 3036 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1619617919
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1619617919
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_15
timestamp 1619617919
transform 1 0 2484 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_21
timestamp 1619617919
transform 1 0 3036 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _294_
timestamp 1619617919
transform 1 0 5336 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _366_
timestamp 1619617919
transform 1 0 4508 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1619617919
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_30
timestamp 1619617919
transform 1 0 3864 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_36
timestamp 1619617919
transform 1 0 4416 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_51
timestamp 1619617919
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_63
timestamp 1619617919
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _254_
timestamp 1619617919
transform 1 0 9936 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _311_
timestamp 1619617919
transform 1 0 8096 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _316_
timestamp 1619617919
transform -1 0 9936 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1619617919
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_75
timestamp 1619617919
transform 1 0 8004 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1619617919
transform 1 0 8924 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _290_
timestamp 1619617919
transform 1 0 10580 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _292_
timestamp 1619617919
transform 1 0 12236 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _371_
timestamp 1619617919
transform -1 0 12052 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_108
timestamp 1619617919
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_119
timestamp 1619617919
transform 1 0 12052 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1619617919
transform 1 0 14812 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen1
timestamp 1619617919
transform 1 0 14352 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb1
timestamp 1619617919
transform 1 0 13340 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1619617919
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_126
timestamp 1619617919
transform 1 0 12696 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_132
timestamp 1619617919
transform 1 0 13248 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_140
timestamp 1619617919
transform 1 0 13984 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1619617919
transform 1 0 16560 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen1
timestamp 1619617919
transform 1 0 16100 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb1
timestamp 1619617919
transform 1 0 15456 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1619617919
transform -1 0 17296 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_152
timestamp 1619617919
transform 1 0 15088 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_171
timestamp 1619617919
transform 1 0 16836 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_7
timestamp 1619617919
transform 1 0 1748 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output40
timestamp 1619617919
transform -1 0 1748 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1619617919
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1619617919
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _364_
timestamp 1619617919
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_15
timestamp 1619617919
transform 1 0 2484 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_12
timestamp 1619617919
transform 1 0 2208 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb1
timestamp 1619617919
transform -1 0 3220 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1619617919
transform 1 0 2576 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_20
timestamp 1619617919
transform 1 0 2944 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen1
timestamp 1619617919
transform 1 0 3220 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_14_33
timestamp 1619617919
transform 1 0 4140 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_28
timestamp 1619617919
transform 1 0 3680 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_28
timestamp 1619617919
transform 1 0 3680 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1619617919
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1619617919
transform 1 0 3864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1619617919
transform 1 0 3956 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_46
timestamp 1619617919
transform 1 0 5336 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1619617919
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1619617919
transform -1 0 5336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_8  _197_
timestamp 1619617919
transform -1 0 5704 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_14_61
timestamp 1619617919
transform 1 0 6716 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_55
timestamp 1619617919
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1619617919
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _305_
timestamp 1619617919
transform 1 0 6072 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _293_
timestamp 1619617919
transform -1 0 6164 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _248_
timestamp 1619617919
transform 1 0 6440 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_13_74
timestamp 1619617919
transform 1 0 7912 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _310_
timestamp 1619617919
transform -1 0 7636 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1619617919
transform -1 0 7912 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1619617919
transform 1 0 6900 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1619617919
transform 1 0 7084 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1619617919
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_1  _309_
timestamp 1619617919
transform 1 0 8004 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _317_
timestamp 1619617919
transform -1 0 9660 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _320_
timestamp 1619617919
transform 1 0 9108 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1619617919
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_80
timestamp 1619617919
transform 1 0 8464 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_86
timestamp 1619617919
transform 1 0 9016 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_93
timestamp 1619617919
transform 1 0 9660 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_80
timestamp 1619617919
transform 1 0 8464 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_96
timestamp 1619617919
transform 1 0 9936 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_105
timestamp 1619617919
transform 1 0 10764 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_101
timestamp 1619617919
transform 1 0 10396 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _318_
timestamp 1619617919
transform 1 0 11040 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _313_
timestamp 1619617919
transform -1 0 10764 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_124
timestamp 1619617919
transform 1 0 12512 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1619617919
transform 1 0 11500 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1619617919
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1619617919
transform 1 0 11684 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_120
timestamp 1619617919
transform 1 0 12144 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_108
timestamp 1619617919
transform 1 0 11040 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1619617919
transform -1 0 14996 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1619617919
transform -1 0 13432 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1619617919
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_134
timestamp 1619617919
transform 1 0 13432 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_146
timestamp 1619617919
transform 1 0 14536 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_132
timestamp 1619617919
transform 1 0 13248 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_140
timestamp 1619617919
transform 1 0 13984 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_144
timestamp 1619617919
transform 1 0 14352 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_159
timestamp 1619617919
transform 1 0 15732 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _373_
timestamp 1619617919
transform -1 0 15732 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_171
timestamp 1619617919
transform 1 0 16836 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_163
timestamp 1619617919
transform 1 0 16100 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_172
timestamp 1619617919
transform 1 0 16928 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1619617919
transform 1 0 16468 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1619617919
transform 1 0 16560 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1619617919
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1619617919
transform -1 0 17296 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1619617919
transform -1 0 17296 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_151
timestamp 1619617919
transform 1 0 14996 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1619617919
transform -1 0 2208 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1619617919
transform -1 0 3220 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1619617919
transform 1 0 2576 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1619617919
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_12
timestamp 1619617919
transform 1 0 2208 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_23
timestamp 1619617919
transform 1 0 3220 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _392_
timestamp 1619617919
transform 1 0 4140 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_15_31
timestamp 1619617919
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1619617919
transform 1 0 6900 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1619617919
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_54
timestamp 1619617919
transform 1 0 6072 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_58
timestamp 1619617919
transform 1 0 6440 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_62
timestamp 1619617919
transform 1 0 6808 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_66
timestamp 1619617919
transform 1 0 7176 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_74
timestamp 1619617919
transform 1 0 7912 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1619617919
transform 1 0 10212 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1619617919
transform 1 0 8188 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1619617919
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_98
timestamp 1619617919
transform 1 0 10120 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1619617919
transform -1 0 11500 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1619617919
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_102
timestamp 1619617919
transform 1 0 10488 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1619617919
transform 1 0 11500 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_115
timestamp 1619617919
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _341_
timestamp 1619617919
transform 1 0 12880 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _385_
timestamp 1619617919
transform 1 0 13800 0 1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_15_127
timestamp 1619617919
transform 1 0 12788 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_131
timestamp 1619617919
transform 1 0 13156 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_137
timestamp 1619617919
transform 1 0 13708 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1619617919
transform -1 0 16468 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1619617919
transform -1 0 17296 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1619617919
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_161
timestamp 1619617919
transform 1 0 15916 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_167
timestamp 1619617919
transform 1 0 16468 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_172
timestamp 1619617919
transform 1 0 16928 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen0
timestamp 1619617919
transform 1 0 2116 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb0
timestamp 1619617919
transform 1 0 1472 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1619617919
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1619617919
transform 1 0 1380 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_16
timestamp 1619617919
transform 1 0 2576 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _246_
timestamp 1619617919
transform 1 0 5152 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _273_
timestamp 1619617919
transform 1 0 4232 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1619617919
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_28
timestamp 1619617919
transform 1 0 3680 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_30
timestamp 1619617919
transform 1 0 3864 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_38
timestamp 1619617919
transform 1 0 4600 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _258_
timestamp 1619617919
transform 1 0 6992 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1619617919
transform -1 0 6992 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _261_
timestamp 1619617919
transform -1 0 8096 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_51
timestamp 1619617919
transform 1 0 5796 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1619617919
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_71
timestamp 1619617919
transform 1 0 7636 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _395_
timestamp 1619617919
transform 1 0 9108 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1619617919
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_76
timestamp 1619617919
transform 1 0 8096 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_84
timestamp 1619617919
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _199_
timestamp 1619617919
transform -1 0 11684 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_4  _386_
timestamp 1619617919
transform -1 0 14076 0 -1 11424
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  FILLER_16_115
timestamp 1619617919
transform 1 0 11684 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _200_
timestamp 1619617919
transform 1 0 14536 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1619617919
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1619617919
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_144
timestamp 1619617919
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _400_
timestamp 1619617919
transform 1 0 15180 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1619617919
transform -1 0 17296 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1619617919
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1619617919
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1619617919
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1619617919
transform -1 0 5244 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _272_
timestamp 1619617919
transform -1 0 4968 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_27
timestamp 1619617919
transform 1 0 3588 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_33
timestamp 1619617919
transform 1 0 4140 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_45
timestamp 1619617919
transform 1 0 5244 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1619617919
transform 1 0 7452 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _260_
timestamp 1619617919
transform 1 0 6716 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1619617919
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_58
timestamp 1619617919
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_72
timestamp 1619617919
transform 1 0 7728 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1619617919
transform -1 0 9752 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_84
timestamp 1619617919
transform 1 0 8832 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_90
timestamp 1619617919
transform 1 0 9384 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_94
timestamp 1619617919
transform 1 0 9752 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1619617919
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_106
timestamp 1619617919
transform 1 0 10856 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_115
timestamp 1619617919
transform 1 0 11684 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1619617919
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1619617919
transform 1 0 13248 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _286_
timestamp 1619617919
transform -1 0 13248 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _287_
timestamp 1619617919
transform 1 0 13524 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _288_
timestamp 1619617919
transform 1 0 14352 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_17_149
timestamp 1619617919
transform 1 0 14812 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _209_
timestamp 1619617919
transform 1 0 15364 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1619617919
transform -1 0 17296 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1619617919
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1619617919
transform -1 0 16836 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_163
timestamp 1619617919
transform 1 0 16100 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1619617919
transform 1 0 16468 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_172
timestamp 1619617919
transform 1 0 16928 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1619617919
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1619617919
transform -1 0 1656 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_6
timestamp 1619617919
transform 1 0 1656 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_18
timestamp 1619617919
transform 1 0 2760 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _270_
timestamp 1619617919
transform -1 0 4232 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1619617919
transform 1 0 4232 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1619617919
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_26
timestamp 1619617919
transform 1 0 3496 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_37
timestamp 1619617919
transform 1 0 4508 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_49
timestamp 1619617919
transform 1 0 5612 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _252_
timestamp 1619617919
transform 1 0 7268 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _256_
timestamp 1619617919
transform -1 0 7084 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_65
timestamp 1619617919
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_74
timestamp 1619617919
transform 1 0 7912 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1619617919
transform 1 0 9384 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp 1619617919
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1619617919
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_87
timestamp 1619617919
transform 1 0 9108 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_96
timestamp 1619617919
transform 1 0 9936 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _401_
timestamp 1619617919
transform 1 0 10304 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_18_120
timestamp 1619617919
transform 1 0 12144 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1619617919
transform 1 0 13892 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _279_
timestamp 1619617919
transform -1 0 13432 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _285_
timestamp 1619617919
transform -1 0 13800 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1619617919
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_128
timestamp 1619617919
transform 1 0 12880 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_138
timestamp 1619617919
transform 1 0 13800 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_142
timestamp 1619617919
transform 1 0 14168 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_144
timestamp 1619617919
transform 1 0 14352 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _210_
timestamp 1619617919
transform 1 0 15180 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1619617919
transform -1 0 17296 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1619617919
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_160
timestamp 1619617919
transform 1 0 15824 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_172
timestamp 1619617919
transform 1 0 16928 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_9
timestamp 1619617919
transform 1 0 1932 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1619617919
transform 1 0 1380 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1619617919
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1619617919
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1619617919
transform 1 0 2024 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_21
timestamp 1619617919
transform 1 0 3036 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_13
timestamp 1619617919
transform 1 0 2300 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _275_
timestamp 1619617919
transform 1 0 3312 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _274_
timestamp 1619617919
transform -1 0 3772 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _391_
timestamp 1619617919
transform -1 0 3312 0 1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__o22a_1  _244_
timestamp 1619617919
transform 1 0 3864 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1619617919
transform 1 0 4048 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _250_
timestamp 1619617919
transform -1 0 5152 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _269_
timestamp 1619617919
transform -1 0 4968 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1619617919
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_35
timestamp 1619617919
transform 1 0 4324 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_44
timestamp 1619617919
transform 1 0 5152 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_42
timestamp 1619617919
transform 1 0 4968 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_62
timestamp 1619617919
transform 1 0 6808 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_50
timestamp 1619617919
transform 1 0 5704 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_56
timestamp 1619617919
transform 1 0 6256 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1619617919
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _263_
timestamp 1619617919
transform -1 0 6808 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _262_
timestamp 1619617919
transform 1 0 5980 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _251_
timestamp 1619617919
transform -1 0 7084 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_19_65
timestamp 1619617919
transform 1 0 7084 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _266_
timestamp 1619617919
transform -1 0 8280 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _265_
timestamp 1619617919
transform 1 0 7176 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1619617919
transform 1 0 7636 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1619617919
transform 1 0 7360 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_74
timestamp 1619617919
transform 1 0 7912 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _394_
timestamp 1619617919
transform 1 0 8280 0 1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1619617919
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_99
timestamp 1619617919
transform 1 0 10212 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_87
timestamp 1619617919
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_99
timestamp 1619617919
transform 1 0 10212 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_103
timestamp 1619617919
transform 1 0 10580 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_103
timestamp 1619617919
transform 1 0 10580 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _224_
timestamp 1619617919
transform 1 0 10672 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _212_
timestamp 1619617919
transform 1 0 10672 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_115
timestamp 1619617919
transform 1 0 11684 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1619617919
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1619617919
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_1  _223_
timestamp 1619617919
transform 1 0 11684 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1619617919
transform -1 0 11684 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_123
timestamp 1619617919
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_122
timestamp 1619617919
transform 1 0 12328 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _207_
timestamp 1619617919
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_135
timestamp 1619617919
transform 1 0 13524 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_126
timestamp 1619617919
transform 1 0 12696 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _343_
timestamp 1619617919
transform -1 0 13524 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _284_
timestamp 1619617919
transform 1 0 12604 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1619617919
transform -1 0 13064 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_144
timestamp 1619617919
transform 1 0 14352 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_147
timestamp 1619617919
transform 1 0 14628 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_142
timestamp 1619617919
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1619617919
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2ai_1  _228_
timestamp 1619617919
transform -1 0 15364 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1619617919
transform 1 0 14352 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_130
timestamp 1619617919
transform 1 0 13064 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_158
timestamp 1619617919
transform 1 0 15640 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _208_
timestamp 1619617919
transform 1 0 14904 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1619617919
transform -1 0 15640 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1619617919
transform 1 0 16284 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_164
timestamp 1619617919
transform 1 0 16192 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1619617919
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1619617919
transform -1 0 16836 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1619617919
transform 1 0 16468 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_168
timestamp 1619617919
transform 1 0 16560 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1619617919
transform -1 0 17296 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1619617919
transform -1 0 17296 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_172
timestamp 1619617919
transform 1 0 16928 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_172
timestamp 1619617919
transform 1 0 16928 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_155
timestamp 1619617919
transform 1 0 15364 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1619617919
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1619617919
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1619617919
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1619617919
transform 1 0 3956 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _268_
timestamp 1619617919
transform 1 0 5244 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1619617919
transform 1 0 3588 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_34
timestamp 1619617919
transform 1 0 4232 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_42
timestamp 1619617919
transform 1 0 4968 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _267_
timestamp 1619617919
transform -1 0 6256 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1619617919
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_56
timestamp 1619617919
transform 1 0 6256 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1619617919
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_70
timestamp 1619617919
transform 1 0 7544 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _219_
timestamp 1619617919
transform 1 0 10120 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _220_
timestamp 1619617919
transform 1 0 9384 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _221_
timestamp 1619617919
transform -1 0 9292 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _222_
timestamp 1619617919
transform -1 0 8832 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_89
timestamp 1619617919
transform 1 0 9292 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _206_
timestamp 1619617919
transform 1 0 10672 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _384_
timestamp 1619617919
transform 1 0 12328 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1619617919
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_107
timestamp 1619617919
transform 1 0 10948 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1619617919
transform 1 0 11500 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_115
timestamp 1619617919
transform 1 0 11684 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1619617919
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_1  _227_
timestamp 1619617919
transform 1 0 14444 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_142
timestamp 1619617919
transform 1 0 14168 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _399_
timestamp 1619617919
transform 1 0 14996 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1619617919
transform -1 0 17296 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1619617919
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_172
timestamp 1619617919
transform 1 0 16928 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _276_
timestamp 1619617919
transform 1 0 2944 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1619617919
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1619617919
transform -1 0 1656 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_6
timestamp 1619617919
transform 1 0 1656 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_18
timestamp 1619617919
transform 1 0 2760 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1619617919
transform 1 0 3956 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _242_
timestamp 1619617919
transform -1 0 3772 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _393_
timestamp 1619617919
transform 1 0 4508 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1619617919
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_30
timestamp 1619617919
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_34
timestamp 1619617919
transform 1 0 4232 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1619617919
transform -1 0 7912 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_58
timestamp 1619617919
transform 1 0 6440 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_70
timestamp 1619617919
transform 1 0 7544 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_74
timestamp 1619617919
transform 1 0 7912 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__o2bb2a_1  _213_
timestamp 1619617919
transform -1 0 10672 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1619617919
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_87
timestamp 1619617919
transform 1 0 9108 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_95
timestamp 1619617919
transform 1 0 9844 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a311o_1  _289_
timestamp 1619617919
transform 1 0 12512 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _402_
timestamp 1619617919
transform -1 0 12512 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1619617919
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_132
timestamp 1619617919
transform 1 0 13248 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_140
timestamp 1619617919
transform 1 0 13984 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_144
timestamp 1619617919
transform 1 0 14352 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _201_
timestamp 1619617919
transform 1 0 14904 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1619617919
transform -1 0 17296 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_157
timestamp 1619617919
transform 1 0 15548 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_169
timestamp 1619617919
transform 1 0 16652 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _277_
timestamp 1619617919
transform 1 0 3220 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _390_
timestamp 1619617919
transform -1 0 3220 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1619617919
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1619617919
transform 1 0 3956 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1619617919
transform -1 0 5704 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_34
timestamp 1619617919
transform 1 0 4232 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_46
timestamp 1619617919
transform 1 0 5336 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1619617919
transform -1 0 7452 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _194_
timestamp 1619617919
transform 1 0 6440 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _237_
timestamp 1619617919
transform 1 0 7452 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_4  _238_
timestamp 1619617919
transform 1 0 7912 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1619617919
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_50
timestamp 1619617919
transform 1 0 5704 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_56
timestamp 1619617919
transform 1 0 6256 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_65
timestamp 1619617919
transform 1 0 7084 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _236_
timestamp 1619617919
transform -1 0 9844 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_95
timestamp 1619617919
transform 1 0 9844 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _198_
timestamp 1619617919
transform 1 0 10580 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1619617919
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_110
timestamp 1619617919
transform 1 0 11224 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_115
timestamp 1619617919
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _231_
timestamp 1619617919
transform -1 0 15364 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _232_
timestamp 1619617919
transform 1 0 13984 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_127
timestamp 1619617919
transform 1 0 12788 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_139
timestamp 1619617919
transform 1 0 13892 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _229_
timestamp 1619617919
transform 1 0 15364 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1619617919
transform -1 0 17296 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1619617919
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1619617919
transform 1 0 16560 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_158
timestamp 1619617919
transform 1 0 15640 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1619617919
transform 1 0 16376 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_172
timestamp 1619617919
transform 1 0 16928 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _240_
timestamp 1619617919
transform 1 0 3036 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1619617919
transform 1 0 1932 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1619617919
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_3
timestamp 1619617919
transform 1 0 1380 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_12
timestamp 1619617919
transform 1 0 2208 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_20
timestamp 1619617919
transform 1 0 2944 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1619617919
transform 1 0 4784 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _241_
timestamp 1619617919
transform -1 0 4140 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1619617919
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_28
timestamp 1619617919
transform 1 0 3680 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_33
timestamp 1619617919
transform 1 0 4140 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_39
timestamp 1619617919
transform 1 0 4692 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_43
timestamp 1619617919
transform 1 0 5060 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a221oi_2  _226_
timestamp 1619617919
transform -1 0 8096 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_55
timestamp 1619617919
transform 1 0 6164 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_63
timestamp 1619617919
transform 1 0 6900 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _214_
timestamp 1619617919
transform -1 0 10488 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1619617919
transform -1 0 9384 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_2  _234_
timestamp 1619617919
transform 1 0 8096 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1619617919
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1619617919
transform 1 0 8924 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_90
timestamp 1619617919
transform 1 0 9384 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_96
timestamp 1619617919
transform 1 0 9936 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _283_
timestamp 1619617919
transform 1 0 11960 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_102
timestamp 1619617919
transform 1 0 10488 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_114
timestamp 1619617919
transform 1 0 11592 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1619617919
transform -1 0 14628 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1619617919
transform 1 0 12788 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp 1619617919
transform -1 0 13616 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1619617919
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_130
timestamp 1619617919
transform 1 0 13064 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_136
timestamp 1619617919
transform 1 0 13616 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_142
timestamp 1619617919
transform 1 0 14168 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_147
timestamp 1619617919
transform 1 0 14628 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp 1619617919
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1619617919
transform -1 0 17296 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1619617919
transform 1 0 15732 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_166
timestamp 1619617919
transform 1 0 16376 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_172
timestamp 1619617919
transform 1 0 16928 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1619617919
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1619617919
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_6
timestamp 1619617919
transform 1 0 1656 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_18
timestamp 1619617919
transform 1 0 2760 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _398_
timestamp 1619617919
transform 1 0 3864 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__a22o_1  _202_
timestamp 1619617919
transform -1 0 6348 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _233_
timestamp 1619617919
transform 1 0 6440 0 1 15776
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1619617919
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_68
timestamp 1619617919
transform 1 0 7360 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _216_
timestamp 1619617919
transform -1 0 10580 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _218_
timestamp 1619617919
transform -1 0 9752 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_80
timestamp 1619617919
transform 1 0 8464 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_88
timestamp 1619617919
transform 1 0 9200 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _215_
timestamp 1619617919
transform -1 0 11316 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _387_
timestamp 1619617919
transform 1 0 12420 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1619617919
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_111
timestamp 1619617919
transform 1 0 11316 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_115
timestamp 1619617919
transform 1 0 11684 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_144
timestamp 1619617919
transform 1 0 14352 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _383_
timestamp 1619617919
transform 1 0 14996 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1619617919
transform -1 0 17296 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1619617919
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_150
timestamp 1619617919
transform 1 0 14904 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_172
timestamp 1619617919
transform 1 0 16928 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_8
timestamp 1619617919
transform 1 0 1840 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1619617919
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1619617919
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1619617919
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _349_
timestamp 1619617919
transform 1 0 1564 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_24
timestamp 1619617919
transform 1 0 3312 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _338_
timestamp 1619617919
transform 1 0 3036 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _278_
timestamp 1619617919
transform 1 0 2392 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1619617919
transform -1 0 3496 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _389_
timestamp 1619617919
transform 1 0 1380 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__or2_1  _204_
timestamp 1619617919
transform -1 0 5704 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1619617919
transform -1 0 4876 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _396_
timestamp 1619617919
transform 1 0 3404 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1619617919
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_26
timestamp 1619617919
transform 1 0 3496 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_30
timestamp 1619617919
transform 1 0 3864 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1619617919
transform 1 0 4876 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _203_
timestamp 1619617919
transform -1 0 7084 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _397_
timestamp 1619617919
transform 1 0 6256 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1619617919
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_53
timestamp 1619617919
transform 1 0 5980 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_50
timestamp 1619617919
transform 1 0 5704 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_56
timestamp 1619617919
transform 1 0 6256 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_65
timestamp 1619617919
transform 1 0 7084 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_73
timestamp 1619617919
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1619617919
transform 1 0 8924 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_79
timestamp 1619617919
transform 1 0 8372 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1619617919
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1619617919
transform 1 0 8096 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_95
timestamp 1619617919
transform 1 0 9844 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_95
timestamp 1619617919
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_87
timestamp 1619617919
transform 1 0 9108 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _205_
timestamp 1619617919
transform 1 0 10028 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _195_
timestamp 1619617919
transform -1 0 10580 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _403_
timestamp 1619617919
transform 1 0 8004 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_27_111
timestamp 1619617919
transform 1 0 11316 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_103
timestamp 1619617919
transform 1 0 10580 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_111
timestamp 1619617919
transform 1 0 11316 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_107
timestamp 1619617919
transform 1 0 10948 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1619617919
transform 1 0 10672 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1619617919
transform 1 0 11040 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1619617919
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_1  _282_
timestamp 1619617919
transform 1 0 11408 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_116
timestamp 1619617919
transform 1 0 11776 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _388_
timestamp 1619617919
transform 1 0 11684 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp 1619617919
transform -1 0 14628 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _381_
timestamp 1619617919
transform 1 0 13616 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1619617919
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_128
timestamp 1619617919
transform 1 0 12880 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_140
timestamp 1619617919
transform 1 0 13984 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_147
timestamp 1619617919
transform 1 0 14628 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_155
timestamp 1619617919
transform 1 0 15364 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1619617919
transform -1 0 15732 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _345_
timestamp 1619617919
transform -1 0 16008 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_172
timestamp 1619617919
transform 1 0 16928 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_165
timestamp 1619617919
transform 1 0 16284 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output42
timestamp 1619617919
transform 1 0 16468 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1619617919
transform 1 0 16008 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1619617919
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1619617919
transform -1 0 17296 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1619617919
transform -1 0 17296 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _193_
timestamp 1619617919
transform -1 0 17020 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1619617919
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1619617919
transform 1 0 1840 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1619617919
transform 1 0 3220 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1619617919
transform 1 0 2116 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output44
timestamp 1619617919
transform -1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1619617919
transform 1 0 1748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_14
timestamp 1619617919
transform 1 0 2392 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_22
timestamp 1619617919
transform 1 0 3128 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 1619617919
transform -1 0 4508 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1619617919
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1619617919
transform 1 0 4600 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_26
timestamp 1619617919
transform 1 0 3496 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_30
timestamp 1619617919
transform 1 0 3864 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_37
timestamp 1619617919
transform 1 0 4508 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1619617919
transform 1 0 4876 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1619617919
transform 1 0 6440 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1619617919
transform 1 0 5980 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1619617919
transform -1 0 7636 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_56
timestamp 1619617919
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_59
timestamp 1619617919
transform 1 0 6532 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_67
timestamp 1619617919
transform 1 0 7268 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_71
timestamp 1619617919
transform 1 0 7636 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp 1619617919
transform -1 0 9016 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1619617919
transform 1 0 9108 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1619617919
transform -1 0 10396 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1619617919
transform 1 0 9200 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_86
timestamp 1619617919
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_91
timestamp 1619617919
transform 1 0 9476 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_97
timestamp 1619617919
transform 1 0 10028 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _339_
timestamp 1619617919
transform -1 0 12604 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1619617919
transform 1 0 11776 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1619617919
transform 1 0 11500 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_101
timestamp 1619617919
transform 1 0 10396 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_117
timestamp 1619617919
transform 1 0 11868 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_121
timestamp 1619617919
transform 1 0 12236 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _382_
timestamp 1619617919
transform 1 0 14720 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1619617919
transform 1 0 14444 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1619617919
transform -1 0 13156 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1619617919
transform 1 0 14168 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_125
timestamp 1619617919
transform 1 0 12604 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_131
timestamp 1619617919
transform 1 0 13156 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_139
timestamp 1619617919
transform 1 0 13892 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_146
timestamp 1619617919
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1619617919
transform -1 0 17296 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1619617919
transform -1 0 17020 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_168
timestamp 1619617919
transform 1 0 16560 0 -1 17952
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 8168 800 8288 6 clockc
port 0 nsew signal tristate
rlabel metal3 s 0 10208 800 10328 6 clockd[0]
port 1 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 clockd[1]
port 2 nsew signal tristate
rlabel metal3 s 17660 17008 18460 17128 6 clockd[2]
port 3 nsew signal tristate
rlabel metal2 s 16578 0 16634 800 6 clockd[3]
port 4 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 clockp[0]
port 5 nsew signal tristate
rlabel metal2 s 1398 0 1454 800 6 clockp[1]
port 6 nsew signal tristate
rlabel metal2 s 12438 0 12494 800 6 dco
port 7 nsew signal input
rlabel metal3 s 17660 12928 18460 13048 6 div[0]
port 8 nsew signal input
rlabel metal2 s 15658 19804 15714 20604 6 div[1]
port 9 nsew signal input
rlabel metal2 s 5998 19804 6054 20604 6 div[2]
port 10 nsew signal input
rlabel metal2 s 478 0 534 800 6 div[3]
port 11 nsew signal input
rlabel metal2 s 11518 19804 11574 20604 6 div[4]
port 12 nsew signal input
rlabel metal2 s 12898 19804 12954 20604 6 ext_trim[0]
port 13 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 ext_trim[10]
port 14 nsew signal input
rlabel metal2 s 1858 19804 1914 20604 6 ext_trim[11]
port 15 nsew signal input
rlabel metal3 s 17660 4768 18460 4888 6 ext_trim[12]
port 16 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 ext_trim[13]
port 17 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 ext_trim[14]
port 18 nsew signal input
rlabel metal3 s 17660 14968 18460 15088 6 ext_trim[15]
port 19 nsew signal input
rlabel metal2 s 3238 19804 3294 20604 6 ext_trim[16]
port 20 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 ext_trim[17]
port 21 nsew signal input
rlabel metal2 s 4618 19804 4674 20604 6 ext_trim[18]
port 22 nsew signal input
rlabel metal3 s 17660 8848 18460 8968 6 ext_trim[19]
port 23 nsew signal input
rlabel metal2 s 10138 19804 10194 20604 6 ext_trim[1]
port 24 nsew signal input
rlabel metal2 s 8758 19804 8814 20604 6 ext_trim[20]
port 25 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 ext_trim[21]
port 26 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 ext_trim[22]
port 27 nsew signal input
rlabel metal3 s 17660 19048 18460 19168 6 ext_trim[23]
port 28 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 ext_trim[24]
port 29 nsew signal input
rlabel metal2 s 7378 19804 7434 20604 6 ext_trim[25]
port 30 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 ext_trim[2]
port 31 nsew signal input
rlabel metal3 s 17660 6808 18460 6928 6 ext_trim[3]
port 32 nsew signal input
rlabel metal3 s 17660 688 18460 808 6 ext_trim[4]
port 33 nsew signal input
rlabel metal3 s 17660 10888 18460 11008 6 ext_trim[5]
port 34 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 ext_trim[6]
port 35 nsew signal input
rlabel metal2 s 478 19804 534 20604 6 ext_trim[7]
port 36 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 ext_trim[8]
port 37 nsew signal input
rlabel metal3 s 17660 2728 18460 2848 6 ext_trim[9]
port 38 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 extclk_sel
port 39 nsew signal input
rlabel metal2 s 14278 19804 14334 20604 6 osc
port 40 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 reset
port 41 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 sel[0]
port 42 nsew signal input
rlabel metal2 s 17038 19804 17094 20604 6 sel[1]
port 43 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 sel[2]
port 44 nsew signal input
rlabel metal4 s 14437 2128 14757 18000 6 VPWR
port 45 nsew power bidirectional
rlabel metal4 s 9040 2128 9360 18000 6 VPWR
port 46 nsew power bidirectional
rlabel metal4 s 3643 2128 3963 18000 6 VPWR
port 47 nsew power bidirectional
rlabel metal5 s 1104 15115 17296 15435 6 VPWR
port 48 nsew power bidirectional
rlabel metal5 s 1104 9856 17296 10176 6 VPWR
port 49 nsew power bidirectional
rlabel metal5 s 1104 4597 17296 4917 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 11739 2128 12059 18000 6 VGND
port 51 nsew ground bidirectional
rlabel metal4 s 6341 2128 6661 18000 6 VGND
port 52 nsew ground bidirectional
rlabel metal5 s 1104 12485 17296 12805 6 VGND
port 53 nsew ground bidirectional
rlabel metal5 s 1104 7227 17296 7547 6 VGND
port 54 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 18460 20604
<< end >>
