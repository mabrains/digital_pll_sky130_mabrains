magic
tech sky130A
magscale 1 2
timestamp 1619593287
<< locali >>
rect 13921 20247 13955 20485
rect 6285 18207 6319 18309
rect 11437 12087 11471 12257
<< viali >>
rect 1501 22729 1535 22763
rect 12265 22661 12299 22695
rect 2329 22525 2363 22559
rect 2789 22525 2823 22559
rect 4629 22525 4663 22559
rect 6009 22525 6043 22559
rect 7849 22525 7883 22559
rect 9873 22525 9907 22559
rect 10885 22525 10919 22559
rect 12449 22525 12483 22559
rect 12909 22525 12943 22559
rect 14933 22525 14967 22559
rect 16681 22525 16715 22559
rect 18153 22525 18187 22559
rect 20453 22525 20487 22559
rect 21097 22525 21131 22559
rect 1593 22457 1627 22491
rect 2145 22389 2179 22423
rect 2973 22389 3007 22423
rect 4813 22389 4847 22423
rect 5825 22389 5859 22423
rect 8033 22389 8067 22423
rect 9689 22389 9723 22423
rect 10701 22389 10735 22423
rect 13093 22389 13127 22423
rect 15117 22389 15151 22423
rect 16497 22389 16531 22423
rect 17969 22389 18003 22423
rect 20269 22389 20303 22423
rect 20913 22389 20947 22423
rect 19993 22185 20027 22219
rect 8401 22049 8435 22083
rect 9505 22049 9539 22083
rect 13093 22049 13127 22083
rect 14933 22049 14967 22083
rect 16681 22049 16715 22083
rect 20177 22049 20211 22083
rect 21097 22049 21131 22083
rect 5181 21981 5215 22015
rect 5457 21981 5491 22015
rect 10701 21981 10735 22015
rect 10977 21981 11011 22015
rect 17325 21981 17359 22015
rect 17601 21981 17635 22015
rect 20913 21913 20947 21947
rect 6929 21845 6963 21879
rect 8585 21845 8619 21879
rect 9689 21845 9723 21879
rect 12449 21845 12483 21879
rect 13277 21845 13311 21879
rect 14749 21845 14783 21879
rect 16865 21845 16899 21879
rect 19073 21845 19107 21879
rect 1777 21641 1811 21675
rect 6837 21641 6871 21675
rect 11069 21641 11103 21675
rect 12081 21641 12115 21675
rect 17325 21641 17359 21675
rect 2513 21573 2547 21607
rect 15209 21573 15243 21607
rect 7481 21505 7515 21539
rect 7757 21505 7791 21539
rect 9689 21505 9723 21539
rect 13277 21505 13311 21539
rect 14749 21505 14783 21539
rect 18797 21505 18831 21539
rect 21005 21505 21039 21539
rect 1961 21437 1995 21471
rect 2697 21437 2731 21471
rect 3433 21437 3467 21471
rect 5089 21437 5123 21471
rect 5733 21437 5767 21471
rect 7021 21437 7055 21471
rect 10057 21437 10091 21471
rect 10517 21437 10551 21471
rect 10885 21437 10919 21471
rect 12265 21437 12299 21471
rect 13001 21437 13035 21471
rect 15393 21437 15427 21471
rect 16037 21437 16071 21471
rect 19073 21437 19107 21471
rect 20177 21437 20211 21471
rect 20361 21437 20395 21471
rect 20913 21437 20947 21471
rect 9873 21369 9907 21403
rect 10701 21369 10735 21403
rect 10793 21369 10827 21403
rect 3617 21301 3651 21335
rect 5273 21301 5307 21335
rect 5917 21301 5951 21335
rect 9229 21301 9263 21335
rect 15853 21301 15887 21335
rect 19901 21301 19935 21335
rect 5825 21097 5859 21131
rect 17509 21097 17543 21131
rect 18153 21097 18187 21131
rect 6193 21029 6227 21063
rect 6331 21029 6365 21063
rect 6018 20961 6052 20995
rect 6112 20961 6146 20995
rect 8217 20961 8251 20995
rect 10609 20961 10643 20995
rect 10793 20961 10827 20995
rect 11069 20961 11103 20995
rect 11437 20961 11471 20995
rect 15209 20961 15243 20995
rect 17693 20961 17727 20995
rect 18337 20961 18371 20995
rect 20177 20961 20211 20995
rect 20913 20961 20947 20995
rect 6469 20893 6503 20927
rect 11253 20893 11287 20927
rect 15485 20893 15519 20927
rect 8401 20757 8435 20791
rect 16957 20757 16991 20791
rect 19993 20757 20027 20791
rect 21005 20757 21039 20791
rect 14013 20553 14047 20587
rect 21097 20553 21131 20587
rect 6929 20485 6963 20519
rect 10609 20485 10643 20519
rect 13921 20485 13955 20519
rect 3249 20417 3283 20451
rect 4997 20417 5031 20451
rect 6837 20417 6871 20451
rect 8401 20417 8435 20451
rect 8677 20417 8711 20451
rect 1409 20349 1443 20383
rect 5641 20349 5675 20383
rect 7021 20349 7055 20383
rect 7113 20349 7147 20383
rect 10793 20349 10827 20383
rect 10885 20349 10919 20383
rect 11161 20349 11195 20383
rect 3525 20281 3559 20315
rect 10977 20281 11011 20315
rect 19625 20417 19659 20451
rect 14197 20349 14231 20383
rect 14289 20349 14323 20383
rect 14565 20349 14599 20383
rect 15025 20349 15059 20383
rect 19349 20349 19383 20383
rect 14381 20281 14415 20315
rect 1593 20213 1627 20247
rect 5549 20213 5583 20247
rect 10149 20213 10183 20247
rect 13921 20213 13955 20247
rect 15117 20213 15151 20247
rect 4813 20009 4847 20043
rect 7573 20009 7607 20043
rect 9505 20009 9539 20043
rect 20637 20009 20671 20043
rect 6193 19941 6227 19975
rect 7205 19941 7239 19975
rect 15025 19941 15059 19975
rect 15117 19941 15151 19975
rect 15945 19941 15979 19975
rect 4997 19873 5031 19907
rect 5089 19873 5123 19907
rect 5365 19873 5399 19907
rect 6377 19873 6411 19907
rect 6469 19873 6503 19907
rect 6745 19873 6779 19907
rect 7389 19873 7423 19907
rect 8033 19873 8067 19907
rect 9689 19873 9723 19907
rect 11897 19873 11931 19907
rect 14933 19873 14967 19907
rect 15301 19873 15335 19907
rect 15761 19873 15795 19907
rect 16037 19873 16071 19907
rect 20821 19873 20855 19907
rect 13185 19805 13219 19839
rect 13553 19805 13587 19839
rect 13645 19805 13679 19839
rect 14749 19737 14783 19771
rect 15761 19737 15795 19771
rect 5273 19669 5307 19703
rect 6653 19669 6687 19703
rect 8125 19669 8159 19703
rect 11805 19669 11839 19703
rect 13829 19669 13863 19703
rect 4445 19465 4479 19499
rect 5825 19465 5859 19499
rect 6929 19465 6963 19499
rect 15117 19465 15151 19499
rect 16405 19465 16439 19499
rect 12633 19329 12667 19363
rect 14105 19329 14139 19363
rect 14197 19329 14231 19363
rect 15945 19329 15979 19363
rect 17693 19329 17727 19363
rect 2421 19261 2455 19295
rect 4629 19261 4663 19295
rect 5733 19261 5767 19295
rect 5917 19261 5951 19295
rect 6837 19261 6871 19295
rect 7757 19261 7791 19295
rect 12173 19261 12207 19295
rect 12357 19261 12391 19295
rect 12449 19261 12483 19295
rect 13829 19261 13863 19295
rect 14013 19261 14047 19295
rect 14381 19261 14415 19295
rect 15025 19261 15059 19295
rect 15669 19261 15703 19295
rect 15853 19261 15887 19295
rect 16037 19261 16071 19295
rect 16221 19261 16255 19295
rect 17877 19261 17911 19295
rect 17969 19261 18003 19295
rect 18521 19261 18555 19295
rect 19441 19261 19475 19295
rect 19625 19261 19659 19295
rect 7849 19193 7883 19227
rect 12725 19193 12759 19227
rect 12817 19193 12851 19227
rect 17693 19193 17727 19227
rect 2605 19125 2639 19159
rect 14565 19125 14599 19159
rect 18613 19125 18647 19159
rect 19533 19125 19567 19159
rect 13461 18921 13495 18955
rect 18889 18921 18923 18955
rect 5825 18853 5859 18887
rect 13645 18853 13679 18887
rect 16221 18853 16255 18887
rect 18981 18853 19015 18887
rect 6009 18785 6043 18819
rect 6469 18785 6503 18819
rect 7389 18785 7423 18819
rect 7849 18785 7883 18819
rect 11713 18785 11747 18819
rect 11805 18785 11839 18819
rect 11989 18785 12023 18819
rect 12265 18785 12299 18819
rect 12541 18785 12575 18819
rect 13829 18785 13863 18819
rect 18613 18785 18647 18819
rect 19073 18785 19107 18819
rect 11161 18717 11195 18751
rect 15945 18717 15979 18751
rect 5641 18581 5675 18615
rect 6561 18581 6595 18615
rect 7297 18581 7331 18615
rect 7941 18581 7975 18615
rect 17693 18581 17727 18615
rect 8309 18377 8343 18411
rect 12081 18377 12115 18411
rect 12449 18377 12483 18411
rect 13829 18377 13863 18411
rect 16313 18377 16347 18411
rect 17325 18377 17359 18411
rect 18245 18377 18279 18411
rect 18797 18377 18831 18411
rect 6285 18309 6319 18343
rect 13001 18309 13035 18343
rect 8861 18241 8895 18275
rect 9045 18241 9079 18275
rect 11069 18241 11103 18275
rect 12173 18241 12207 18275
rect 4537 18173 4571 18207
rect 5365 18173 5399 18207
rect 5457 18173 5491 18207
rect 5825 18173 5859 18207
rect 6285 18173 6319 18207
rect 7021 18173 7055 18207
rect 8033 18173 8067 18207
rect 8125 18173 8159 18207
rect 8401 18173 8435 18207
rect 9137 18173 9171 18207
rect 9873 18173 9907 18207
rect 10977 18173 11011 18207
rect 12081 18173 12115 18207
rect 13093 18173 13127 18207
rect 13737 18173 13771 18207
rect 13921 18173 13955 18207
rect 16221 18173 16255 18207
rect 16405 18173 16439 18207
rect 17509 18173 17543 18207
rect 18337 18173 18371 18207
rect 18981 18173 19015 18207
rect 19165 18173 19199 18207
rect 19257 18173 19291 18207
rect 19349 18173 19383 18207
rect 19533 18173 19567 18207
rect 21097 18173 21131 18207
rect 5181 18105 5215 18139
rect 5549 18105 5583 18139
rect 5687 18105 5721 18139
rect 6837 18105 6871 18139
rect 4721 18037 4755 18071
rect 7205 18037 7239 18071
rect 7849 18037 7883 18071
rect 8861 18037 8895 18071
rect 10057 18037 10091 18071
rect 20913 18037 20947 18071
rect 6561 17833 6595 17867
rect 8309 17833 8343 17867
rect 12725 17833 12759 17867
rect 15209 17833 15243 17867
rect 15393 17833 15427 17867
rect 4537 17765 4571 17799
rect 7941 17765 7975 17799
rect 8033 17765 8067 17799
rect 9781 17765 9815 17799
rect 1409 17697 1443 17731
rect 4261 17697 4295 17731
rect 6745 17697 6779 17731
rect 6837 17697 6871 17731
rect 7113 17697 7147 17731
rect 7665 17697 7699 17731
rect 7758 17697 7792 17731
rect 8130 17697 8164 17731
rect 9505 17697 9539 17731
rect 11989 17697 12023 17731
rect 12357 17697 12391 17731
rect 12817 17697 12851 17731
rect 15268 17697 15302 17731
rect 17601 17697 17635 17731
rect 19073 17697 19107 17731
rect 19993 17697 20027 17731
rect 20177 17697 20211 17731
rect 20269 17697 20303 17731
rect 20407 17697 20441 17731
rect 12081 17629 12115 17663
rect 12541 17629 12575 17663
rect 14749 17629 14783 17663
rect 1593 17493 1627 17527
rect 6009 17493 6043 17527
rect 7021 17493 7055 17527
rect 11253 17493 11287 17527
rect 14841 17493 14875 17527
rect 17417 17493 17451 17527
rect 18981 17493 19015 17527
rect 20545 17493 20579 17527
rect 8033 17289 8067 17323
rect 8125 17289 8159 17323
rect 12081 17289 12115 17323
rect 18889 17289 18923 17323
rect 21097 17289 21131 17323
rect 7113 17153 7147 17187
rect 7205 17153 7239 17187
rect 7941 17153 7975 17187
rect 19625 17153 19659 17187
rect 5917 17085 5951 17119
rect 7021 17085 7055 17119
rect 7297 17085 7331 17119
rect 7481 17085 7515 17119
rect 8217 17085 8251 17119
rect 8677 17085 8711 17119
rect 15485 17085 15519 17119
rect 17509 17085 17543 17119
rect 17601 17085 17635 17119
rect 17877 17085 17911 17119
rect 17969 17085 18003 17119
rect 18429 17085 18463 17119
rect 18705 17085 18739 17119
rect 19349 17085 19383 17119
rect 5825 17017 5859 17051
rect 12265 17017 12299 17051
rect 12449 17017 12483 17051
rect 15209 17017 15243 17051
rect 17693 17017 17727 17051
rect 6837 16949 6871 16983
rect 8769 16949 8803 16983
rect 13737 16949 13771 16983
rect 17325 16949 17359 16983
rect 18521 16949 18555 16983
rect 1869 16745 1903 16779
rect 2513 16745 2547 16779
rect 11437 16745 11471 16779
rect 12081 16745 12115 16779
rect 15301 16745 15335 16779
rect 18061 16745 18095 16779
rect 20085 16745 20119 16779
rect 20821 16745 20855 16779
rect 14933 16677 14967 16711
rect 16589 16677 16623 16711
rect 1685 16609 1719 16643
rect 2329 16609 2363 16643
rect 7297 16609 7331 16643
rect 7389 16609 7423 16643
rect 11805 16609 11839 16643
rect 11897 16609 11931 16643
rect 13645 16609 13679 16643
rect 13829 16609 13863 16643
rect 14749 16609 14783 16643
rect 15021 16609 15055 16643
rect 15163 16609 15197 16643
rect 16313 16609 16347 16643
rect 18889 16609 18923 16643
rect 19993 16609 20027 16643
rect 20177 16609 20211 16643
rect 21005 16609 21039 16643
rect 18981 16541 19015 16575
rect 13829 16473 13863 16507
rect 2697 16201 2731 16235
rect 12817 16201 12851 16235
rect 19165 16201 19199 16235
rect 20729 16201 20763 16235
rect 7021 16133 7055 16167
rect 17325 16133 17359 16167
rect 3341 16065 3375 16099
rect 6837 16065 6871 16099
rect 8769 16065 8803 16099
rect 8953 16065 8987 16099
rect 13369 16065 13403 16099
rect 13921 16065 13955 16099
rect 17877 16065 17911 16099
rect 2605 15997 2639 16031
rect 7113 15997 7147 16031
rect 9045 15997 9079 16031
rect 10517 15997 10551 16031
rect 12998 15997 13032 16031
rect 13461 15997 13495 16031
rect 14105 15997 14139 16031
rect 14381 15997 14415 16031
rect 17509 15997 17543 16031
rect 18981 15997 19015 16031
rect 19165 15997 19199 16031
rect 19533 15997 19567 16031
rect 20913 15997 20947 16031
rect 3617 15929 3651 15963
rect 17693 15929 17727 15963
rect 5089 15861 5123 15895
rect 6837 15861 6871 15895
rect 8769 15861 8803 15895
rect 10701 15861 10735 15895
rect 13001 15861 13035 15895
rect 14289 15861 14323 15895
rect 17601 15861 17635 15895
rect 19441 15861 19475 15895
rect 4445 15657 4479 15691
rect 5089 15657 5123 15691
rect 14749 15657 14783 15691
rect 16957 15657 16991 15691
rect 20913 15657 20947 15691
rect 5365 15589 5399 15623
rect 9781 15589 9815 15623
rect 1409 15521 1443 15555
rect 4629 15521 4663 15555
rect 5273 15521 5307 15555
rect 5457 15521 5491 15555
rect 5595 15521 5629 15555
rect 6377 15521 6411 15555
rect 6837 15521 6871 15555
rect 6930 15521 6964 15555
rect 7067 15521 7101 15555
rect 7205 15521 7239 15555
rect 7302 15521 7336 15555
rect 7941 15521 7975 15555
rect 8034 15521 8068 15555
rect 8217 15521 8251 15555
rect 8309 15521 8343 15555
rect 8447 15521 8481 15555
rect 9505 15521 9539 15555
rect 15025 15521 15059 15555
rect 17049 15521 17083 15555
rect 18337 15521 18371 15555
rect 21097 15521 21131 15555
rect 5733 15453 5767 15487
rect 6285 15453 6319 15487
rect 14933 15453 14967 15487
rect 15301 15453 15335 15487
rect 15393 15453 15427 15487
rect 1593 15317 1627 15351
rect 7481 15317 7515 15351
rect 8585 15317 8619 15351
rect 11253 15317 11287 15351
rect 18245 15317 18279 15351
rect 4997 15113 5031 15147
rect 5549 15113 5583 15147
rect 8401 15113 8435 15147
rect 8953 15113 8987 15147
rect 10149 15113 10183 15147
rect 14381 15113 14415 15147
rect 15485 15113 15519 15147
rect 17325 15113 17359 15147
rect 17509 15113 17543 15147
rect 7205 15045 7239 15079
rect 7941 15045 7975 15079
rect 9413 15045 9447 15079
rect 18337 15045 18371 15079
rect 7113 14977 7147 15011
rect 7481 14977 7515 15011
rect 9965 14977 9999 15011
rect 14933 14977 14967 15011
rect 16313 14977 16347 15011
rect 17601 14977 17635 15011
rect 1869 14909 1903 14943
rect 4905 14909 4939 14943
rect 5089 14909 5123 14943
rect 5733 14909 5767 14943
rect 6837 14909 6871 14943
rect 7021 14909 7055 14943
rect 7297 14909 7331 14943
rect 8125 14909 8159 14943
rect 8217 14909 8251 14943
rect 8493 14909 8527 14943
rect 9137 14909 9171 14943
rect 9229 14909 9263 14943
rect 9505 14909 9539 14943
rect 10241 14909 10275 14943
rect 12541 14909 12575 14943
rect 14562 14909 14596 14943
rect 15025 14909 15059 14943
rect 15485 14909 15519 14943
rect 15761 14909 15795 14943
rect 16405 14909 16439 14943
rect 17693 14909 17727 14943
rect 18521 14909 18555 14943
rect 18705 14909 18739 14943
rect 18889 14909 18923 14943
rect 19349 14909 19383 14943
rect 5917 14841 5951 14875
rect 18613 14841 18647 14875
rect 19625 14841 19659 14875
rect 2053 14773 2087 14807
rect 2697 14773 2731 14807
rect 2789 14773 2823 14807
rect 9965 14773 9999 14807
rect 12357 14773 12391 14807
rect 14565 14773 14599 14807
rect 15669 14773 15703 14807
rect 21097 14773 21131 14807
rect 6193 14569 6227 14603
rect 7297 14569 7331 14603
rect 8493 14569 8527 14603
rect 9965 14569 9999 14603
rect 10609 14569 10643 14603
rect 19993 14569 20027 14603
rect 20177 14569 20211 14603
rect 6469 14501 6503 14535
rect 6561 14501 6595 14535
rect 11437 14501 11471 14535
rect 15025 14501 15059 14535
rect 15117 14501 15151 14535
rect 2329 14433 2363 14467
rect 6377 14433 6411 14467
rect 6745 14433 6779 14467
rect 7389 14433 7423 14467
rect 8401 14433 8435 14467
rect 9873 14433 9907 14467
rect 10517 14433 10551 14467
rect 14933 14433 14967 14467
rect 15301 14433 15335 14467
rect 16221 14433 16255 14467
rect 16957 14433 16991 14467
rect 17141 14433 17175 14467
rect 18061 14433 18095 14467
rect 18337 14433 18371 14467
rect 18429 14433 18463 14467
rect 18613 14433 18647 14467
rect 20174 14433 20208 14467
rect 20545 14433 20579 14467
rect 1961 14365 1995 14399
rect 2789 14365 2823 14399
rect 3157 14365 3191 14399
rect 11161 14365 11195 14399
rect 17049 14365 17083 14399
rect 17233 14365 17267 14399
rect 18245 14365 18279 14399
rect 20637 14365 20671 14399
rect 16313 14297 16347 14331
rect 2329 14229 2363 14263
rect 2973 14229 3007 14263
rect 12909 14229 12943 14263
rect 14749 14229 14783 14263
rect 17417 14229 17451 14263
rect 17877 14229 17911 14263
rect 1961 14025 1995 14059
rect 8585 14025 8619 14059
rect 15761 14025 15795 14059
rect 17417 14025 17451 14059
rect 17509 14025 17543 14059
rect 19441 14025 19475 14059
rect 20729 14025 20763 14059
rect 3525 13957 3559 13991
rect 3985 13957 4019 13991
rect 9505 13957 9539 13991
rect 2421 13889 2455 13923
rect 2513 13889 2547 13923
rect 3157 13889 3191 13923
rect 10149 13889 10183 13923
rect 14289 13889 14323 13923
rect 17325 13889 17359 13923
rect 4169 13821 4203 13855
rect 8677 13821 8711 13855
rect 9965 13821 9999 13855
rect 14013 13821 14047 13855
rect 17601 13821 17635 13855
rect 18061 13821 18095 13855
rect 18245 13821 18279 13855
rect 19579 13821 19613 13855
rect 19717 13821 19751 13855
rect 19993 13821 20027 13855
rect 20913 13821 20947 13855
rect 2329 13753 2363 13787
rect 19809 13753 19843 13787
rect 3525 13685 3559 13719
rect 9873 13685 9907 13719
rect 18429 13685 18463 13719
rect 2421 13481 2455 13515
rect 3157 13481 3191 13515
rect 4629 13481 4663 13515
rect 6745 13481 6779 13515
rect 8309 13481 8343 13515
rect 9873 13481 9907 13515
rect 15025 13481 15059 13515
rect 15577 13481 15611 13515
rect 4721 13413 4755 13447
rect 16221 13413 16255 13447
rect 17969 13413 18003 13447
rect 2053 13345 2087 13379
rect 2421 13345 2455 13379
rect 3341 13345 3375 13379
rect 5825 13345 5859 13379
rect 6929 13345 6963 13379
rect 7113 13345 7147 13379
rect 7573 13345 7607 13379
rect 8401 13345 8435 13379
rect 10149 13345 10183 13379
rect 10609 13345 10643 13379
rect 12265 13345 12299 13379
rect 14933 13345 14967 13379
rect 15117 13345 15151 13379
rect 15761 13345 15795 13379
rect 4813 13277 4847 13311
rect 5641 13277 5675 13311
rect 5917 13277 5951 13311
rect 6009 13277 6043 13311
rect 6101 13277 6135 13311
rect 11989 13277 12023 13311
rect 12173 13277 12207 13311
rect 18245 13277 18279 13311
rect 7665 13209 7699 13243
rect 10241 13209 10275 13243
rect 10333 13209 10367 13243
rect 4261 13141 4295 13175
rect 6929 13141 6963 13175
rect 10425 13141 10459 13175
rect 12633 13141 12667 13175
rect 1501 12937 1535 12971
rect 3157 12937 3191 12971
rect 3985 12937 4019 12971
rect 9413 12937 9447 12971
rect 9781 12869 9815 12903
rect 2789 12801 2823 12835
rect 3617 12801 3651 12835
rect 9505 12801 9539 12835
rect 12265 12801 12299 12835
rect 12449 12801 12483 12835
rect 18245 12801 18279 12835
rect 18521 12801 18555 12835
rect 20269 12801 20303 12835
rect 3985 12733 4019 12767
rect 6837 12733 6871 12767
rect 7021 12733 7055 12767
rect 8217 12733 8251 12767
rect 8585 12733 8619 12767
rect 9413 12733 9447 12767
rect 10977 12733 11011 12767
rect 11161 12733 11195 12767
rect 13553 12733 13587 12767
rect 21097 12733 21131 12767
rect 1593 12665 1627 12699
rect 3157 12665 3191 12699
rect 8401 12665 8435 12699
rect 13369 12665 13403 12699
rect 7113 12597 7147 12631
rect 11069 12597 11103 12631
rect 12541 12597 12575 12631
rect 12909 12597 12943 12631
rect 13737 12597 13771 12631
rect 20913 12597 20947 12631
rect 4353 12393 4387 12427
rect 11897 12393 11931 12427
rect 12357 12393 12391 12427
rect 15117 12393 15151 12427
rect 15209 12393 15243 12427
rect 17325 12393 17359 12427
rect 19993 12393 20027 12427
rect 6101 12325 6135 12359
rect 6469 12325 6503 12359
rect 11713 12325 11747 12359
rect 4261 12257 4295 12291
rect 6285 12257 6319 12291
rect 7205 12257 7239 12291
rect 7941 12257 7975 12291
rect 8217 12257 8251 12291
rect 10057 12257 10091 12291
rect 10241 12257 10275 12291
rect 10425 12257 10459 12291
rect 10517 12257 10551 12291
rect 11437 12257 11471 12291
rect 11529 12257 11563 12291
rect 12541 12257 12575 12291
rect 12633 12257 12667 12291
rect 17509 12257 17543 12291
rect 20177 12257 20211 12291
rect 20913 12257 20947 12291
rect 7849 12189 7883 12223
rect 10333 12189 10367 12223
rect 10793 12121 10827 12155
rect 15301 12189 15335 12223
rect 7297 12053 7331 12087
rect 11437 12053 11471 12087
rect 14749 12053 14783 12087
rect 20729 12053 20763 12087
rect 5825 11849 5859 11883
rect 3709 11781 3743 11815
rect 13277 11781 13311 11815
rect 1961 11713 1995 11747
rect 2145 11713 2179 11747
rect 3525 11713 3559 11747
rect 6837 11713 6871 11747
rect 8861 11713 8895 11747
rect 10609 11713 10643 11747
rect 12909 11713 12943 11747
rect 15577 11713 15611 11747
rect 3893 11645 3927 11679
rect 4537 11645 4571 11679
rect 5641 11645 5675 11679
rect 5917 11645 5951 11679
rect 8585 11645 8619 11679
rect 8677 11645 8711 11679
rect 8769 11645 8803 11679
rect 10701 11645 10735 11679
rect 10885 11645 10919 11679
rect 11069 11645 11103 11679
rect 13921 11645 13955 11679
rect 15761 11645 15795 11679
rect 20913 11645 20947 11679
rect 2237 11577 2271 11611
rect 5457 11577 5491 11611
rect 7021 11577 7055 11611
rect 7205 11577 7239 11611
rect 13277 11577 13311 11611
rect 15853 11577 15887 11611
rect 2605 11509 2639 11543
rect 4353 11509 4387 11543
rect 9045 11509 9079 11543
rect 13737 11509 13771 11543
rect 16221 11509 16255 11543
rect 20729 11509 20763 11543
rect 4261 11305 4295 11339
rect 5549 11305 5583 11339
rect 6377 11305 6411 11339
rect 11253 11305 11287 11339
rect 11621 11305 11655 11339
rect 13277 11305 13311 11339
rect 15117 11305 15151 11339
rect 15945 11305 15979 11339
rect 16773 11305 16807 11339
rect 5641 11237 5675 11271
rect 10333 11237 10367 11271
rect 2237 11169 2271 11203
rect 4261 11169 4295 11203
rect 4629 11169 4663 11203
rect 6561 11169 6595 11203
rect 7757 11169 7791 11203
rect 7849 11169 7883 11203
rect 8401 11169 8435 11203
rect 9597 11169 9631 11203
rect 9689 11169 9723 11203
rect 9873 11169 9907 11203
rect 11713 11169 11747 11203
rect 12909 11169 12943 11203
rect 13277 11169 13311 11203
rect 15577 11169 15611 11203
rect 16405 11169 16439 11203
rect 16773 11169 16807 11203
rect 17417 11169 17451 11203
rect 5733 11101 5767 11135
rect 6653 11101 6687 11135
rect 6745 11101 6779 11135
rect 6837 11101 6871 11135
rect 7389 11101 7423 11135
rect 7573 11101 7607 11135
rect 7665 11101 7699 11135
rect 11897 11101 11931 11135
rect 5181 11033 5215 11067
rect 15945 11033 15979 11067
rect 17233 11033 17267 11067
rect 2421 10965 2455 10999
rect 8493 10965 8527 10999
rect 15025 10965 15059 10999
rect 3801 10761 3835 10795
rect 8217 10761 8251 10795
rect 8953 10761 8987 10795
rect 9689 10761 9723 10795
rect 10517 10761 10551 10795
rect 14473 10761 14507 10795
rect 20729 10761 20763 10795
rect 9045 10693 9079 10727
rect 15117 10693 15151 10727
rect 16129 10693 16163 10727
rect 1869 10625 1903 10659
rect 3065 10625 3099 10659
rect 8401 10625 8435 10659
rect 9137 10625 9171 10659
rect 9873 10625 9907 10659
rect 13185 10625 13219 10659
rect 13369 10625 13403 10659
rect 2237 10557 2271 10591
rect 2697 10557 2731 10591
rect 3985 10557 4019 10591
rect 8125 10557 8159 10591
rect 8861 10557 8895 10591
rect 9597 10557 9631 10591
rect 12633 10557 12667 10591
rect 13461 10557 13495 10591
rect 14657 10557 14691 10591
rect 15485 10557 15519 10591
rect 15945 10557 15979 10591
rect 20913 10557 20947 10591
rect 9873 10489 9907 10523
rect 10496 10489 10530 10523
rect 10701 10489 10735 10523
rect 16313 10489 16347 10523
rect 2237 10421 2271 10455
rect 2697 10421 2731 10455
rect 8401 10421 8435 10455
rect 10333 10421 10367 10455
rect 12541 10421 12575 10455
rect 13829 10421 13863 10455
rect 15117 10421 15151 10455
rect 1501 10217 1535 10251
rect 2329 10217 2363 10251
rect 2973 10217 3007 10251
rect 6009 10217 6043 10251
rect 7113 10217 7147 10251
rect 7481 10217 7515 10251
rect 15945 10217 15979 10251
rect 20913 10217 20947 10251
rect 13001 10149 13035 10183
rect 1593 10081 1627 10115
rect 2513 10081 2547 10115
rect 5917 10081 5951 10115
rect 8125 10081 8159 10115
rect 8401 10081 8435 10115
rect 9505 10081 9539 10115
rect 10517 10081 10551 10115
rect 10701 10081 10735 10115
rect 15761 10081 15795 10115
rect 21097 10081 21131 10115
rect 6101 10013 6135 10047
rect 6837 10013 6871 10047
rect 7021 10013 7055 10047
rect 8217 10013 8251 10047
rect 8309 10013 8343 10047
rect 10425 10013 10459 10047
rect 12633 10013 12667 10047
rect 10885 9945 10919 9979
rect 3065 9877 3099 9911
rect 5549 9877 5583 9911
rect 7941 9877 7975 9911
rect 9597 9877 9631 9911
rect 12909 9877 12943 9911
rect 8861 9673 8895 9707
rect 10057 9673 10091 9707
rect 15485 9673 15519 9707
rect 12909 9605 12943 9639
rect 2697 9537 2731 9571
rect 4169 9537 4203 9571
rect 5549 9537 5583 9571
rect 10149 9537 10183 9571
rect 15117 9537 15151 9571
rect 2145 9469 2179 9503
rect 5181 9469 5215 9503
rect 7481 9469 7515 9503
rect 7665 9469 7699 9503
rect 7757 9469 7791 9503
rect 8953 9469 8987 9503
rect 9873 9469 9907 9503
rect 12265 9469 12299 9503
rect 13277 9469 13311 9503
rect 2605 9401 2639 9435
rect 4629 9401 4663 9435
rect 4721 9401 4755 9435
rect 12081 9401 12115 9435
rect 15485 9401 15519 9435
rect 5181 9333 5215 9367
rect 7297 9333 7331 9367
rect 9689 9333 9723 9367
rect 12449 9333 12483 9367
rect 12909 9333 12943 9367
rect 2053 9129 2087 9163
rect 2421 9129 2455 9163
rect 9965 9129 9999 9163
rect 13093 9129 13127 9163
rect 15669 9129 15703 9163
rect 7205 9061 7239 9095
rect 7389 9061 7423 9095
rect 1409 8993 1443 9027
rect 4261 8993 4295 9027
rect 4813 8993 4847 9027
rect 5641 8993 5675 9027
rect 6285 8993 6319 9027
rect 7113 8993 7147 9027
rect 9873 8993 9907 9027
rect 11069 8993 11103 9027
rect 12081 8993 12115 9027
rect 13185 8993 13219 9027
rect 16129 8993 16163 9027
rect 20913 8993 20947 9027
rect 2513 8925 2547 8959
rect 2697 8925 2731 8959
rect 4629 8925 4663 8959
rect 5273 8925 5307 8959
rect 10149 8925 10183 8959
rect 10977 8925 11011 8959
rect 13277 8925 13311 8959
rect 15301 8925 15335 8959
rect 6101 8857 6135 8891
rect 12725 8857 12759 8891
rect 15669 8857 15703 8891
rect 16221 8857 16255 8891
rect 1593 8789 1627 8823
rect 5273 8789 5307 8823
rect 7665 8789 7699 8823
rect 9505 8789 9539 8823
rect 10701 8789 10735 8823
rect 10885 8789 10919 8823
rect 11897 8789 11931 8823
rect 20729 8789 20763 8823
rect 1685 8585 1719 8619
rect 4905 8585 4939 8619
rect 9505 8585 9539 8619
rect 9873 8585 9907 8619
rect 20729 8585 20763 8619
rect 14933 8517 14967 8551
rect 15761 8517 15795 8551
rect 16221 8517 16255 8551
rect 9413 8449 9447 8483
rect 13093 8449 13127 8483
rect 13277 8449 13311 8483
rect 1501 8381 1535 8415
rect 2145 8381 2179 8415
rect 2697 8381 2731 8415
rect 3398 8381 3432 8415
rect 4997 8381 5031 8415
rect 9689 8381 9723 8415
rect 14565 8381 14599 8415
rect 15393 8381 15427 8415
rect 16405 8381 16439 8415
rect 20913 8381 20947 8415
rect 2605 8313 2639 8347
rect 14933 8313 14967 8347
rect 3295 8245 3329 8279
rect 10977 8245 11011 8279
rect 11069 8245 11103 8279
rect 12633 8245 12667 8279
rect 13001 8245 13035 8279
rect 15761 8245 15795 8279
rect 6101 8041 6135 8075
rect 9873 8041 9907 8075
rect 13001 8041 13035 8075
rect 15025 8041 15059 8075
rect 15485 8041 15519 8075
rect 15853 8041 15887 8075
rect 20913 8041 20947 8075
rect 11253 7973 11287 8007
rect 6285 7905 6319 7939
rect 7665 7905 7699 7939
rect 8217 7905 8251 7939
rect 10793 7905 10827 7939
rect 11345 7905 11379 7939
rect 11989 7905 12023 7939
rect 12817 7905 12851 7939
rect 14841 7905 14875 7939
rect 15945 7905 15979 7939
rect 21097 7905 21131 7939
rect 9597 7837 9631 7871
rect 9781 7837 9815 7871
rect 16037 7837 16071 7871
rect 10241 7701 10275 7735
rect 11805 7701 11839 7735
rect 13093 7497 13127 7531
rect 13737 7497 13771 7531
rect 10241 7429 10275 7463
rect 11069 7429 11103 7463
rect 9873 7361 9907 7395
rect 12081 7361 12115 7395
rect 13277 7361 13311 7395
rect 14105 7361 14139 7395
rect 2973 7293 3007 7327
rect 5181 7293 5215 7327
rect 5733 7293 5767 7327
rect 10701 7293 10735 7327
rect 12449 7293 12483 7327
rect 13737 7293 13771 7327
rect 17693 7293 17727 7327
rect 12909 7225 12943 7259
rect 17509 7225 17543 7259
rect 2881 7157 2915 7191
rect 4813 7157 4847 7191
rect 10241 7157 10275 7191
rect 11069 7157 11103 7191
rect 12081 7157 12115 7191
rect 4997 6953 5031 6987
rect 10885 6953 10919 6987
rect 11253 6953 11287 6987
rect 13185 6953 13219 6987
rect 1961 6817 1995 6851
rect 2605 6817 2639 6851
rect 6837 6817 6871 6851
rect 11345 6817 11379 6851
rect 13829 6817 13863 6851
rect 20729 6817 20763 6851
rect 4721 6749 4755 6783
rect 4905 6749 4939 6783
rect 11437 6749 11471 6783
rect 12817 6749 12851 6783
rect 1777 6681 1811 6715
rect 2421 6681 2455 6715
rect 5365 6681 5399 6715
rect 13185 6681 13219 6715
rect 13645 6681 13679 6715
rect 20913 6681 20947 6715
rect 6837 6613 6871 6647
rect 13185 6409 13219 6443
rect 13737 6409 13771 6443
rect 19717 6409 19751 6443
rect 20729 6409 20763 6443
rect 9597 6341 9631 6375
rect 14289 6341 14323 6375
rect 2421 6273 2455 6307
rect 8217 6273 8251 6307
rect 10241 6273 10275 6307
rect 12817 6273 12851 6307
rect 14749 6273 14783 6307
rect 14933 6273 14967 6307
rect 15485 6273 15519 6307
rect 15669 6273 15703 6307
rect 17969 6273 18003 6307
rect 4445 6205 4479 6239
rect 7665 6205 7699 6239
rect 9137 6205 9171 6239
rect 12173 6205 12207 6239
rect 13645 6205 13679 6239
rect 15853 6205 15887 6239
rect 16129 6205 16163 6239
rect 17693 6205 17727 6239
rect 20913 6205 20947 6239
rect 2697 6137 2731 6171
rect 7481 6137 7515 6171
rect 8861 6137 8895 6171
rect 13185 6137 13219 6171
rect 7297 6069 7331 6103
rect 9965 6069 9999 6103
rect 10057 6069 10091 6103
rect 12357 6069 12391 6103
rect 14657 6069 14691 6103
rect 9873 5865 9907 5899
rect 10425 5865 10459 5899
rect 14841 5865 14875 5899
rect 15209 5865 15243 5899
rect 16129 5865 16163 5899
rect 16497 5865 16531 5899
rect 17325 5865 17359 5899
rect 17785 5865 17819 5899
rect 20729 5865 20763 5899
rect 6561 5797 6595 5831
rect 8309 5797 8343 5831
rect 1593 5729 1627 5763
rect 5917 5729 5951 5763
rect 6653 5729 6687 5763
rect 7665 5729 7699 5763
rect 8585 5729 8619 5763
rect 9505 5729 9539 5763
rect 10333 5729 10367 5763
rect 11897 5729 11931 5763
rect 17693 5729 17727 5763
rect 20913 5729 20947 5763
rect 12265 5661 12299 5695
rect 15301 5661 15335 5695
rect 15485 5661 15519 5695
rect 16589 5661 16623 5695
rect 16681 5661 16715 5695
rect 17877 5661 17911 5695
rect 9873 5593 9907 5627
rect 1501 5525 1535 5559
rect 12265 5525 12299 5559
rect 1777 5321 1811 5355
rect 5641 5321 5675 5355
rect 6929 5321 6963 5355
rect 8953 5321 8987 5355
rect 9781 5321 9815 5355
rect 18153 5321 18187 5355
rect 20913 5321 20947 5355
rect 12449 5253 12483 5287
rect 12909 5253 12943 5287
rect 2789 5185 2823 5219
rect 9137 5185 9171 5219
rect 12081 5185 12115 5219
rect 15669 5185 15703 5219
rect 19901 5185 19935 5219
rect 20177 5185 20211 5219
rect 1961 5117 1995 5151
rect 2513 5117 2547 5151
rect 4537 5117 4571 5151
rect 5733 5117 5767 5151
rect 7113 5117 7147 5151
rect 9597 5117 9631 5151
rect 13093 5117 13127 5151
rect 15853 5117 15887 5151
rect 16037 5117 16071 5151
rect 16221 5117 16255 5151
rect 17509 5117 17543 5151
rect 21097 5117 21131 5151
rect 5917 5049 5951 5083
rect 8769 5049 8803 5083
rect 12449 4981 12483 5015
rect 17417 4981 17451 5015
rect 5825 4777 5859 4811
rect 6653 4777 6687 4811
rect 10517 4777 10551 4811
rect 11713 4777 11747 4811
rect 12541 4777 12575 4811
rect 16405 4777 16439 4811
rect 17785 4709 17819 4743
rect 5917 4641 5951 4675
rect 12541 4641 12575 4675
rect 13277 4641 13311 4675
rect 16405 4641 16439 4675
rect 16681 4641 16715 4675
rect 17233 4641 17267 4675
rect 17417 4641 17451 4675
rect 10241 4573 10275 4607
rect 10425 4573 10459 4607
rect 11345 4573 11379 4607
rect 12173 4573 12207 4607
rect 16221 4573 16255 4607
rect 17601 4573 17635 4607
rect 10885 4505 10919 4539
rect 11713 4505 11747 4539
rect 13093 4505 13127 4539
rect 12173 4233 12207 4267
rect 13277 4233 13311 4267
rect 16313 4233 16347 4267
rect 3525 4097 3559 4131
rect 13277 4097 13311 4131
rect 2053 4029 2087 4063
rect 3341 4029 3375 4063
rect 8033 4029 8067 4063
rect 10793 4029 10827 4063
rect 12265 4029 12299 4063
rect 13645 4029 13679 4063
rect 16221 4029 16255 4063
rect 20269 4029 20303 4063
rect 8677 3961 8711 3995
rect 8953 3961 8987 3995
rect 14105 3961 14139 3995
rect 1869 3893 1903 3927
rect 10701 3893 10735 3927
rect 14197 3893 14231 3927
rect 20453 3893 20487 3927
rect 13369 3689 13403 3723
rect 15117 3689 15151 3723
rect 20913 3689 20947 3723
rect 6009 3621 6043 3655
rect 8309 3621 8343 3655
rect 1409 3553 1443 3587
rect 6193 3553 6227 3587
rect 7665 3553 7699 3587
rect 8585 3553 8619 3587
rect 9505 3553 9539 3587
rect 10517 3553 10551 3587
rect 11437 3553 11471 3587
rect 12173 3553 12207 3587
rect 13369 3553 13403 3587
rect 15209 3553 15243 3587
rect 21097 3553 21131 3587
rect 9873 3485 9907 3519
rect 13737 3485 13771 3519
rect 15393 3485 15427 3519
rect 11989 3417 12023 3451
rect 14749 3417 14783 3451
rect 1593 3349 1627 3383
rect 9505 3349 9539 3383
rect 10333 3349 10367 3383
rect 11253 3349 11287 3383
rect 2053 3145 2087 3179
rect 4629 3145 4663 3179
rect 7021 3145 7055 3179
rect 8769 3145 8803 3179
rect 9321 3145 9355 3179
rect 18061 3145 18095 3179
rect 20729 3145 20763 3179
rect 10241 3077 10275 3111
rect 13921 3077 13955 3111
rect 14565 3077 14599 3111
rect 17325 3077 17359 3111
rect 20269 3077 20303 3111
rect 9321 3009 9355 3043
rect 9689 3009 9723 3043
rect 10701 3009 10735 3043
rect 10885 3009 10919 3043
rect 12725 3009 12759 3043
rect 12817 3009 12851 3043
rect 15393 3009 15427 3043
rect 1869 2941 1903 2975
rect 2513 2941 2547 2975
rect 4445 2941 4479 2975
rect 6837 2941 6871 2975
rect 8861 2941 8895 2975
rect 10609 2941 10643 2975
rect 13737 2941 13771 2975
rect 14749 2941 14783 2975
rect 16129 2941 16163 2975
rect 18245 2941 18279 2975
rect 20085 2941 20119 2975
rect 20913 2941 20947 2975
rect 12909 2873 12943 2907
rect 14105 2873 14139 2907
rect 17509 2873 17543 2907
rect 2697 2805 2731 2839
rect 13277 2805 13311 2839
rect 2605 2601 2639 2635
rect 4445 2601 4479 2635
rect 5733 2601 5767 2635
rect 6929 2601 6963 2635
rect 9781 2601 9815 2635
rect 10701 2601 10735 2635
rect 13185 2601 13219 2635
rect 16129 2601 16163 2635
rect 17601 2601 17635 2635
rect 18889 2601 18923 2635
rect 2053 2533 2087 2567
rect 15301 2533 15335 2567
rect 15485 2533 15519 2567
rect 20913 2533 20947 2567
rect 2789 2465 2823 2499
rect 4261 2465 4295 2499
rect 5549 2465 5583 2499
rect 7113 2465 7147 2499
rect 8493 2465 8527 2499
rect 9597 2465 9631 2499
rect 10517 2465 10551 2499
rect 11161 2465 11195 2499
rect 12817 2465 12851 2499
rect 13829 2465 13863 2499
rect 15945 2465 15979 2499
rect 17785 2465 17819 2499
rect 19073 2465 19107 2499
rect 1869 2329 1903 2363
rect 8677 2329 8711 2363
rect 13185 2329 13219 2363
rect 13645 2329 13679 2363
rect 20729 2329 20763 2363
rect 11345 2261 11379 2295
<< metal1 >>
rect 1104 22874 21804 22896
rect 1104 22822 4432 22874
rect 4484 22822 4496 22874
rect 4548 22822 4560 22874
rect 4612 22822 4624 22874
rect 4676 22822 11332 22874
rect 11384 22822 11396 22874
rect 11448 22822 11460 22874
rect 11512 22822 11524 22874
rect 11576 22822 18232 22874
rect 18284 22822 18296 22874
rect 18348 22822 18360 22874
rect 18412 22822 18424 22874
rect 18476 22822 21804 22874
rect 1104 22800 21804 22822
rect 1486 22760 1492 22772
rect 1447 22732 1492 22760
rect 1486 22720 1492 22732
rect 1544 22720 1550 22772
rect 12253 22695 12311 22701
rect 12253 22661 12265 22695
rect 12299 22661 12311 22695
rect 12253 22655 12311 22661
rect 934 22516 940 22568
rect 992 22556 998 22568
rect 2317 22559 2375 22565
rect 2317 22556 2329 22559
rect 992 22528 2329 22556
rect 992 22516 998 22528
rect 2317 22525 2329 22528
rect 2363 22525 2375 22559
rect 2774 22556 2780 22568
rect 2735 22528 2780 22556
rect 2317 22519 2375 22525
rect 2774 22516 2780 22528
rect 2832 22516 2838 22568
rect 4617 22559 4675 22565
rect 4617 22525 4629 22559
rect 4663 22556 4675 22559
rect 4798 22556 4804 22568
rect 4663 22528 4804 22556
rect 4663 22525 4675 22528
rect 4617 22519 4675 22525
rect 4798 22516 4804 22528
rect 4856 22516 4862 22568
rect 5994 22556 6000 22568
rect 5955 22528 6000 22556
rect 5994 22516 6000 22528
rect 6052 22516 6058 22568
rect 7834 22556 7840 22568
rect 7795 22528 7840 22556
rect 7834 22516 7840 22528
rect 7892 22516 7898 22568
rect 9674 22516 9680 22568
rect 9732 22556 9738 22568
rect 9861 22559 9919 22565
rect 9861 22556 9873 22559
rect 9732 22528 9873 22556
rect 9732 22516 9738 22528
rect 9861 22525 9873 22528
rect 9907 22525 9919 22559
rect 9861 22519 9919 22525
rect 10873 22559 10931 22565
rect 10873 22525 10885 22559
rect 10919 22556 10931 22559
rect 12268 22556 12296 22655
rect 10919 22528 12296 22556
rect 12437 22559 12495 22565
rect 10919 22525 10931 22528
rect 10873 22519 10931 22525
rect 12437 22525 12449 22559
rect 12483 22525 12495 22559
rect 12894 22556 12900 22568
rect 12855 22528 12900 22556
rect 12437 22519 12495 22525
rect 1578 22488 1584 22500
rect 1539 22460 1584 22488
rect 1578 22448 1584 22460
rect 1636 22448 1642 22500
rect 11698 22448 11704 22500
rect 11756 22488 11762 22500
rect 12452 22488 12480 22519
rect 12894 22516 12900 22528
rect 12952 22516 12958 22568
rect 14734 22516 14740 22568
rect 14792 22556 14798 22568
rect 14921 22559 14979 22565
rect 14921 22556 14933 22559
rect 14792 22528 14933 22556
rect 14792 22516 14798 22528
rect 14921 22525 14933 22528
rect 14967 22525 14979 22559
rect 14921 22519 14979 22525
rect 16574 22516 16580 22568
rect 16632 22556 16638 22568
rect 16669 22559 16727 22565
rect 16669 22556 16681 22559
rect 16632 22528 16681 22556
rect 16632 22516 16638 22528
rect 16669 22525 16681 22528
rect 16715 22525 16727 22559
rect 16669 22519 16727 22525
rect 17954 22516 17960 22568
rect 18012 22556 18018 22568
rect 18141 22559 18199 22565
rect 18141 22556 18153 22559
rect 18012 22528 18153 22556
rect 18012 22516 18018 22528
rect 18141 22525 18153 22528
rect 18187 22525 18199 22559
rect 18141 22519 18199 22525
rect 19794 22516 19800 22568
rect 19852 22556 19858 22568
rect 20441 22559 20499 22565
rect 20441 22556 20453 22559
rect 19852 22528 20453 22556
rect 19852 22516 19858 22528
rect 20441 22525 20453 22528
rect 20487 22525 20499 22559
rect 21082 22556 21088 22568
rect 21043 22528 21088 22556
rect 20441 22519 20499 22525
rect 21082 22516 21088 22528
rect 21140 22516 21146 22568
rect 11756 22460 12480 22488
rect 11756 22448 11762 22460
rect 1670 22380 1676 22432
rect 1728 22420 1734 22432
rect 2133 22423 2191 22429
rect 2133 22420 2145 22423
rect 1728 22392 2145 22420
rect 1728 22380 1734 22392
rect 2133 22389 2145 22392
rect 2179 22389 2191 22423
rect 2133 22383 2191 22389
rect 2961 22423 3019 22429
rect 2961 22389 2973 22423
rect 3007 22420 3019 22423
rect 3418 22420 3424 22432
rect 3007 22392 3424 22420
rect 3007 22389 3019 22392
rect 2961 22383 3019 22389
rect 3418 22380 3424 22392
rect 3476 22380 3482 22432
rect 4801 22423 4859 22429
rect 4801 22389 4813 22423
rect 4847 22420 4859 22423
rect 5074 22420 5080 22432
rect 4847 22392 5080 22420
rect 4847 22389 4859 22392
rect 4801 22383 4859 22389
rect 5074 22380 5080 22392
rect 5132 22380 5138 22432
rect 5718 22380 5724 22432
rect 5776 22420 5782 22432
rect 5813 22423 5871 22429
rect 5813 22420 5825 22423
rect 5776 22392 5825 22420
rect 5776 22380 5782 22392
rect 5813 22389 5825 22392
rect 5859 22389 5871 22423
rect 5813 22383 5871 22389
rect 8021 22423 8079 22429
rect 8021 22389 8033 22423
rect 8067 22420 8079 22423
rect 8202 22420 8208 22432
rect 8067 22392 8208 22420
rect 8067 22389 8079 22392
rect 8021 22383 8079 22389
rect 8202 22380 8208 22392
rect 8260 22380 8266 22432
rect 9674 22420 9680 22432
rect 9635 22392 9680 22420
rect 9674 22380 9680 22392
rect 9732 22380 9738 22432
rect 10318 22380 10324 22432
rect 10376 22420 10382 22432
rect 10689 22423 10747 22429
rect 10689 22420 10701 22423
rect 10376 22392 10701 22420
rect 10376 22380 10382 22392
rect 10689 22389 10701 22392
rect 10735 22389 10747 22423
rect 13078 22420 13084 22432
rect 13039 22392 13084 22420
rect 10689 22383 10747 22389
rect 13078 22380 13084 22392
rect 13136 22380 13142 22432
rect 15105 22423 15163 22429
rect 15105 22389 15117 22423
rect 15151 22420 15163 22423
rect 15378 22420 15384 22432
rect 15151 22392 15384 22420
rect 15151 22389 15163 22392
rect 15105 22383 15163 22389
rect 15378 22380 15384 22392
rect 15436 22380 15442 22432
rect 16022 22380 16028 22432
rect 16080 22420 16086 22432
rect 16485 22423 16543 22429
rect 16485 22420 16497 22423
rect 16080 22392 16497 22420
rect 16080 22380 16086 22392
rect 16485 22389 16497 22392
rect 16531 22389 16543 22423
rect 16485 22383 16543 22389
rect 16666 22380 16672 22432
rect 16724 22420 16730 22432
rect 17957 22423 18015 22429
rect 17957 22420 17969 22423
rect 16724 22392 17969 22420
rect 16724 22380 16730 22392
rect 17957 22389 17969 22392
rect 18003 22389 18015 22423
rect 17957 22383 18015 22389
rect 20162 22380 20168 22432
rect 20220 22420 20226 22432
rect 20257 22423 20315 22429
rect 20257 22420 20269 22423
rect 20220 22392 20269 22420
rect 20220 22380 20226 22392
rect 20257 22389 20269 22392
rect 20303 22389 20315 22423
rect 20257 22383 20315 22389
rect 20901 22423 20959 22429
rect 20901 22389 20913 22423
rect 20947 22420 20959 22423
rect 21358 22420 21364 22432
rect 20947 22392 21364 22420
rect 20947 22389 20959 22392
rect 20901 22383 20959 22389
rect 21358 22380 21364 22392
rect 21416 22380 21422 22432
rect 1104 22330 21804 22352
rect 1104 22278 7882 22330
rect 7934 22278 7946 22330
rect 7998 22278 8010 22330
rect 8062 22278 8074 22330
rect 8126 22278 14782 22330
rect 14834 22278 14846 22330
rect 14898 22278 14910 22330
rect 14962 22278 14974 22330
rect 15026 22278 21804 22330
rect 1104 22256 21804 22278
rect 19981 22219 20039 22225
rect 19981 22216 19993 22219
rect 18800 22188 19993 22216
rect 6822 22148 6828 22160
rect 6670 22120 6828 22148
rect 6822 22108 6828 22120
rect 6880 22108 6886 22160
rect 18800 22134 18828 22188
rect 19981 22185 19993 22188
rect 20027 22185 20039 22219
rect 19981 22179 20039 22185
rect 7006 22040 7012 22092
rect 7064 22080 7070 22092
rect 8389 22083 8447 22089
rect 8389 22080 8401 22083
rect 7064 22052 8401 22080
rect 7064 22040 7070 22052
rect 8389 22049 8401 22052
rect 8435 22049 8447 22083
rect 8389 22043 8447 22049
rect 9493 22083 9551 22089
rect 9493 22049 9505 22083
rect 9539 22080 9551 22083
rect 9674 22080 9680 22092
rect 9539 22052 9680 22080
rect 9539 22049 9551 22052
rect 9493 22043 9551 22049
rect 5166 22012 5172 22024
rect 5127 21984 5172 22012
rect 5166 21972 5172 21984
rect 5224 21972 5230 22024
rect 5445 22015 5503 22021
rect 5445 21981 5457 22015
rect 5491 22012 5503 22015
rect 5810 22012 5816 22024
rect 5491 21984 5816 22012
rect 5491 21981 5503 21984
rect 5445 21975 5503 21981
rect 5810 21972 5816 21984
rect 5868 21972 5874 22024
rect 8404 22012 8432 22043
rect 9674 22040 9680 22052
rect 9732 22040 9738 22092
rect 12066 22040 12072 22092
rect 12124 22040 12130 22092
rect 13078 22080 13084 22092
rect 13039 22052 13084 22080
rect 13078 22040 13084 22052
rect 13136 22040 13142 22092
rect 14921 22083 14979 22089
rect 14921 22049 14933 22083
rect 14967 22049 14979 22083
rect 16666 22080 16672 22092
rect 16627 22052 16672 22080
rect 14921 22043 14979 22049
rect 9766 22012 9772 22024
rect 8404 21984 9772 22012
rect 9766 21972 9772 21984
rect 9824 21972 9830 22024
rect 10686 22012 10692 22024
rect 10647 21984 10692 22012
rect 10686 21972 10692 21984
rect 10744 21972 10750 22024
rect 10965 22015 11023 22021
rect 10965 21981 10977 22015
rect 11011 22012 11023 22015
rect 11054 22012 11060 22024
rect 11011 21984 11060 22012
rect 11011 21981 11023 21984
rect 10965 21975 11023 21981
rect 11054 21972 11060 21984
rect 11112 21972 11118 22024
rect 12250 21972 12256 22024
rect 12308 22012 12314 22024
rect 14936 22012 14964 22043
rect 16666 22040 16672 22052
rect 16724 22040 16730 22092
rect 20165 22083 20223 22089
rect 20165 22049 20177 22083
rect 20211 22080 20223 22083
rect 20806 22080 20812 22092
rect 20211 22052 20812 22080
rect 20211 22049 20223 22052
rect 20165 22043 20223 22049
rect 20806 22040 20812 22052
rect 20864 22040 20870 22092
rect 21085 22083 21143 22089
rect 21085 22049 21097 22083
rect 21131 22080 21143 22083
rect 21634 22080 21640 22092
rect 21131 22052 21640 22080
rect 21131 22049 21143 22052
rect 21085 22043 21143 22049
rect 21634 22040 21640 22052
rect 21692 22040 21698 22092
rect 12308 21984 14964 22012
rect 17313 22015 17371 22021
rect 12308 21972 12314 21984
rect 17313 21981 17325 22015
rect 17359 21981 17371 22015
rect 17586 22012 17592 22024
rect 17547 21984 17592 22012
rect 17313 21975 17371 21981
rect 15194 21904 15200 21956
rect 15252 21944 15258 21956
rect 17328 21944 17356 21975
rect 17586 21972 17592 21984
rect 17644 21972 17650 22024
rect 17678 21972 17684 22024
rect 17736 22012 17742 22024
rect 17736 21984 20944 22012
rect 17736 21972 17742 21984
rect 20916 21953 20944 21984
rect 15252 21916 17356 21944
rect 20901 21947 20959 21953
rect 15252 21904 15258 21916
rect 20901 21913 20913 21947
rect 20947 21913 20959 21947
rect 20901 21907 20959 21913
rect 6454 21836 6460 21888
rect 6512 21876 6518 21888
rect 6917 21879 6975 21885
rect 6917 21876 6929 21879
rect 6512 21848 6929 21876
rect 6512 21836 6518 21848
rect 6917 21845 6929 21848
rect 6963 21845 6975 21879
rect 6917 21839 6975 21845
rect 8478 21836 8484 21888
rect 8536 21876 8542 21888
rect 8573 21879 8631 21885
rect 8573 21876 8585 21879
rect 8536 21848 8585 21876
rect 8536 21836 8542 21848
rect 8573 21845 8585 21848
rect 8619 21845 8631 21879
rect 8573 21839 8631 21845
rect 9677 21879 9735 21885
rect 9677 21845 9689 21879
rect 9723 21876 9735 21879
rect 10226 21876 10232 21888
rect 9723 21848 10232 21876
rect 9723 21845 9735 21848
rect 9677 21839 9735 21845
rect 10226 21836 10232 21848
rect 10284 21836 10290 21888
rect 10962 21836 10968 21888
rect 11020 21876 11026 21888
rect 12437 21879 12495 21885
rect 12437 21876 12449 21879
rect 11020 21848 12449 21876
rect 11020 21836 11026 21848
rect 12437 21845 12449 21848
rect 12483 21845 12495 21879
rect 12437 21839 12495 21845
rect 13265 21879 13323 21885
rect 13265 21845 13277 21879
rect 13311 21876 13323 21879
rect 13354 21876 13360 21888
rect 13311 21848 13360 21876
rect 13311 21845 13323 21848
rect 13265 21839 13323 21845
rect 13354 21836 13360 21848
rect 13412 21836 13418 21888
rect 14642 21836 14648 21888
rect 14700 21876 14706 21888
rect 14737 21879 14795 21885
rect 14737 21876 14749 21879
rect 14700 21848 14749 21876
rect 14700 21836 14706 21848
rect 14737 21845 14749 21848
rect 14783 21845 14795 21879
rect 16850 21876 16856 21888
rect 16811 21848 16856 21876
rect 14737 21839 14795 21845
rect 16850 21836 16856 21848
rect 16908 21836 16914 21888
rect 19061 21879 19119 21885
rect 19061 21845 19073 21879
rect 19107 21876 19119 21879
rect 19978 21876 19984 21888
rect 19107 21848 19984 21876
rect 19107 21845 19119 21848
rect 19061 21839 19119 21845
rect 19978 21836 19984 21848
rect 20036 21836 20042 21888
rect 1104 21786 21804 21808
rect 1104 21734 4432 21786
rect 4484 21734 4496 21786
rect 4548 21734 4560 21786
rect 4612 21734 4624 21786
rect 4676 21734 11332 21786
rect 11384 21734 11396 21786
rect 11448 21734 11460 21786
rect 11512 21734 11524 21786
rect 11576 21734 18232 21786
rect 18284 21734 18296 21786
rect 18348 21734 18360 21786
rect 18412 21734 18424 21786
rect 18476 21734 21804 21786
rect 1104 21712 21804 21734
rect 1578 21632 1584 21684
rect 1636 21672 1642 21684
rect 1765 21675 1823 21681
rect 1765 21672 1777 21675
rect 1636 21644 1777 21672
rect 1636 21632 1642 21644
rect 1765 21641 1777 21644
rect 1811 21641 1823 21675
rect 6822 21672 6828 21684
rect 6783 21644 6828 21672
rect 1765 21635 1823 21641
rect 6822 21632 6828 21644
rect 6880 21632 6886 21684
rect 8386 21672 8392 21684
rect 7484 21644 8392 21672
rect 2501 21607 2559 21613
rect 2501 21573 2513 21607
rect 2547 21573 2559 21607
rect 3234 21604 3240 21616
rect 2501 21567 2559 21573
rect 2746 21576 3240 21604
rect 1949 21471 2007 21477
rect 1949 21437 1961 21471
rect 1995 21468 2007 21471
rect 2516 21468 2544 21567
rect 2746 21536 2774 21576
rect 3234 21564 3240 21576
rect 3292 21604 3298 21616
rect 5166 21604 5172 21616
rect 3292 21576 5172 21604
rect 3292 21564 3298 21576
rect 5166 21564 5172 21576
rect 5224 21604 5230 21616
rect 7484 21604 7512 21644
rect 8386 21632 8392 21644
rect 8444 21672 8450 21684
rect 11054 21672 11060 21684
rect 8444 21644 9674 21672
rect 11015 21644 11060 21672
rect 8444 21632 8450 21644
rect 5224 21576 7512 21604
rect 9646 21604 9674 21644
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 12066 21672 12072 21684
rect 12027 21644 12072 21672
rect 12066 21632 12072 21644
rect 12124 21632 12130 21684
rect 17313 21675 17371 21681
rect 17313 21641 17325 21675
rect 17359 21672 17371 21675
rect 17586 21672 17592 21684
rect 17359 21644 17592 21672
rect 17359 21641 17371 21644
rect 17313 21635 17371 21641
rect 17586 21632 17592 21644
rect 17644 21632 17650 21684
rect 10686 21604 10692 21616
rect 9646 21576 10692 21604
rect 5224 21564 5230 21576
rect 7484 21545 7512 21576
rect 10686 21564 10692 21576
rect 10744 21604 10750 21616
rect 10744 21576 13032 21604
rect 10744 21564 10750 21576
rect 2700 21508 2774 21536
rect 7469 21539 7527 21545
rect 2700 21477 2728 21508
rect 7469 21505 7481 21539
rect 7515 21505 7527 21539
rect 7469 21499 7527 21505
rect 7745 21539 7803 21545
rect 7745 21505 7757 21539
rect 7791 21536 7803 21539
rect 9677 21539 9735 21545
rect 9677 21536 9689 21539
rect 7791 21508 9689 21536
rect 7791 21505 7803 21508
rect 7745 21499 7803 21505
rect 9677 21505 9689 21508
rect 9723 21505 9735 21539
rect 11054 21536 11060 21548
rect 9677 21499 9735 21505
rect 10520 21508 11060 21536
rect 1995 21440 2544 21468
rect 2685 21471 2743 21477
rect 1995 21437 2007 21440
rect 1949 21431 2007 21437
rect 2685 21437 2697 21471
rect 2731 21437 2743 21471
rect 3418 21468 3424 21480
rect 3379 21440 3424 21468
rect 2685 21431 2743 21437
rect 3418 21428 3424 21440
rect 3476 21428 3482 21480
rect 5074 21468 5080 21480
rect 5035 21440 5080 21468
rect 5074 21428 5080 21440
rect 5132 21428 5138 21480
rect 5718 21468 5724 21480
rect 5679 21440 5724 21468
rect 5718 21428 5724 21440
rect 5776 21428 5782 21480
rect 7006 21468 7012 21480
rect 6919 21440 7012 21468
rect 7006 21428 7012 21440
rect 7064 21428 7070 21480
rect 10520 21477 10548 21508
rect 11054 21496 11060 21508
rect 11112 21496 11118 21548
rect 10045 21471 10103 21477
rect 10045 21437 10057 21471
rect 10091 21468 10103 21471
rect 10505 21471 10563 21477
rect 10505 21468 10517 21471
rect 10091 21440 10517 21468
rect 10091 21437 10103 21440
rect 10045 21431 10103 21437
rect 10505 21437 10517 21440
rect 10551 21437 10563 21471
rect 10505 21431 10563 21437
rect 10873 21471 10931 21477
rect 10873 21437 10885 21471
rect 10919 21468 10931 21471
rect 11146 21468 11152 21480
rect 10919 21440 11152 21468
rect 10919 21437 10931 21440
rect 10873 21431 10931 21437
rect 11146 21428 11152 21440
rect 11204 21428 11210 21480
rect 12250 21468 12256 21480
rect 12163 21440 12256 21468
rect 12250 21428 12256 21440
rect 12308 21428 12314 21480
rect 13004 21477 13032 21576
rect 14274 21564 14280 21616
rect 14332 21604 14338 21616
rect 15197 21607 15255 21613
rect 15197 21604 15209 21607
rect 14332 21576 15209 21604
rect 14332 21564 14338 21576
rect 15197 21573 15209 21576
rect 15243 21573 15255 21607
rect 15197 21567 15255 21573
rect 19978 21564 19984 21616
rect 20036 21604 20042 21616
rect 20036 21576 21036 21604
rect 20036 21564 20042 21576
rect 13265 21539 13323 21545
rect 13265 21505 13277 21539
rect 13311 21536 13323 21539
rect 13998 21536 14004 21548
rect 13311 21508 14004 21536
rect 13311 21505 13323 21508
rect 13265 21499 13323 21505
rect 13998 21496 14004 21508
rect 14056 21496 14062 21548
rect 14737 21539 14795 21545
rect 14737 21505 14749 21539
rect 14783 21536 14795 21539
rect 15102 21536 15108 21548
rect 14783 21508 15108 21536
rect 14783 21505 14795 21508
rect 14737 21499 14795 21505
rect 15102 21496 15108 21508
rect 15160 21496 15166 21548
rect 16850 21496 16856 21548
rect 16908 21536 16914 21548
rect 21008 21545 21036 21576
rect 18785 21539 18843 21545
rect 18785 21536 18797 21539
rect 16908 21508 18797 21536
rect 16908 21496 16914 21508
rect 18785 21505 18797 21508
rect 18831 21505 18843 21539
rect 18785 21499 18843 21505
rect 20993 21539 21051 21545
rect 20993 21505 21005 21539
rect 21039 21505 21051 21539
rect 20993 21499 21051 21505
rect 12989 21471 13047 21477
rect 12989 21437 13001 21471
rect 13035 21437 13047 21471
rect 15378 21468 15384 21480
rect 15339 21440 15384 21468
rect 12989 21431 13047 21437
rect 5350 21360 5356 21412
rect 5408 21400 5414 21412
rect 7024 21400 7052 21428
rect 5408 21372 7052 21400
rect 5408 21360 5414 21372
rect 8478 21360 8484 21412
rect 8536 21360 8542 21412
rect 9861 21403 9919 21409
rect 9861 21369 9873 21403
rect 9907 21369 9919 21403
rect 9861 21363 9919 21369
rect 10689 21403 10747 21409
rect 10689 21369 10701 21403
rect 10735 21369 10747 21403
rect 10689 21363 10747 21369
rect 10781 21403 10839 21409
rect 10781 21369 10793 21403
rect 10827 21400 10839 21403
rect 10962 21400 10968 21412
rect 10827 21372 10968 21400
rect 10827 21369 10839 21372
rect 10781 21363 10839 21369
rect 3605 21335 3663 21341
rect 3605 21301 3617 21335
rect 3651 21332 3663 21335
rect 3694 21332 3700 21344
rect 3651 21304 3700 21332
rect 3651 21301 3663 21304
rect 3605 21295 3663 21301
rect 3694 21292 3700 21304
rect 3752 21292 3758 21344
rect 5261 21335 5319 21341
rect 5261 21301 5273 21335
rect 5307 21332 5319 21335
rect 5442 21332 5448 21344
rect 5307 21304 5448 21332
rect 5307 21301 5319 21304
rect 5261 21295 5319 21301
rect 5442 21292 5448 21304
rect 5500 21292 5506 21344
rect 5902 21332 5908 21344
rect 5863 21304 5908 21332
rect 5902 21292 5908 21304
rect 5960 21292 5966 21344
rect 9217 21335 9275 21341
rect 9217 21301 9229 21335
rect 9263 21332 9275 21335
rect 9876 21332 9904 21363
rect 10594 21332 10600 21344
rect 9263 21304 10600 21332
rect 9263 21301 9275 21304
rect 9217 21295 9275 21301
rect 10594 21292 10600 21304
rect 10652 21332 10658 21344
rect 10704 21332 10732 21363
rect 10962 21360 10968 21372
rect 11020 21360 11026 21412
rect 10652 21304 10732 21332
rect 10652 21292 10658 21304
rect 10870 21292 10876 21344
rect 10928 21332 10934 21344
rect 12268 21332 12296 21428
rect 10928 21304 12296 21332
rect 13004 21332 13032 21431
rect 15378 21428 15384 21440
rect 15436 21428 15442 21480
rect 16022 21468 16028 21480
rect 15983 21440 16028 21468
rect 16022 21428 16028 21440
rect 16080 21428 16086 21480
rect 19061 21471 19119 21477
rect 19061 21437 19073 21471
rect 19107 21468 19119 21471
rect 19334 21468 19340 21480
rect 19107 21440 19340 21468
rect 19107 21437 19119 21440
rect 19061 21431 19119 21437
rect 19334 21428 19340 21440
rect 19392 21428 19398 21480
rect 19978 21428 19984 21480
rect 20036 21468 20042 21480
rect 20165 21471 20223 21477
rect 20165 21468 20177 21471
rect 20036 21440 20177 21468
rect 20036 21428 20042 21440
rect 20165 21437 20177 21440
rect 20211 21437 20223 21471
rect 20165 21431 20223 21437
rect 20349 21471 20407 21477
rect 20349 21437 20361 21471
rect 20395 21437 20407 21471
rect 20349 21431 20407 21437
rect 20901 21471 20959 21477
rect 20901 21437 20913 21471
rect 20947 21468 20959 21471
rect 21082 21468 21088 21480
rect 20947 21440 21088 21468
rect 20947 21437 20959 21440
rect 20901 21431 20959 21437
rect 14642 21400 14648 21412
rect 14490 21372 14648 21400
rect 14642 21360 14648 21372
rect 14700 21360 14706 21412
rect 18138 21360 18144 21412
rect 18196 21360 18202 21412
rect 20364 21400 20392 21431
rect 20916 21400 20944 21431
rect 21082 21428 21088 21440
rect 21140 21428 21146 21480
rect 20364 21372 20944 21400
rect 15194 21332 15200 21344
rect 13004 21304 15200 21332
rect 10928 21292 10934 21304
rect 15194 21292 15200 21304
rect 15252 21292 15258 21344
rect 15838 21332 15844 21344
rect 15799 21304 15844 21332
rect 15838 21292 15844 21304
rect 15896 21292 15902 21344
rect 19886 21332 19892 21344
rect 19847 21304 19892 21332
rect 19886 21292 19892 21304
rect 19944 21292 19950 21344
rect 1104 21242 21804 21264
rect 1104 21190 7882 21242
rect 7934 21190 7946 21242
rect 7998 21190 8010 21242
rect 8062 21190 8074 21242
rect 8126 21190 14782 21242
rect 14834 21190 14846 21242
rect 14898 21190 14910 21242
rect 14962 21190 14974 21242
rect 15026 21190 21804 21242
rect 1104 21168 21804 21190
rect 5810 21128 5816 21140
rect 5771 21100 5816 21128
rect 5810 21088 5816 21100
rect 5868 21088 5874 21140
rect 9766 21088 9772 21140
rect 9824 21128 9830 21140
rect 10870 21128 10876 21140
rect 9824 21100 10876 21128
rect 9824 21088 9830 21100
rect 10870 21088 10876 21100
rect 10928 21088 10934 21140
rect 17497 21131 17555 21137
rect 17497 21097 17509 21131
rect 17543 21097 17555 21131
rect 18138 21128 18144 21140
rect 18099 21100 18144 21128
rect 17497 21091 17555 21097
rect 5718 21020 5724 21072
rect 5776 21060 5782 21072
rect 6181 21063 6239 21069
rect 6181 21060 6193 21063
rect 5776 21032 6193 21060
rect 5776 21020 5782 21032
rect 6181 21029 6193 21032
rect 6227 21029 6239 21063
rect 6181 21023 6239 21029
rect 6319 21063 6377 21069
rect 6319 21029 6331 21063
rect 6365 21060 6377 21063
rect 6454 21060 6460 21072
rect 6365 21032 6460 21060
rect 6365 21029 6377 21032
rect 6319 21023 6377 21029
rect 6454 21020 6460 21032
rect 6512 21020 6518 21072
rect 10962 21020 10968 21072
rect 11020 21060 11026 21072
rect 15562 21060 15568 21072
rect 11020 21032 11468 21060
rect 11020 21020 11026 21032
rect 5810 20952 5816 21004
rect 5868 20992 5874 21004
rect 6006 20995 6064 21001
rect 6006 20992 6018 20995
rect 5868 20964 6018 20992
rect 5868 20952 5874 20964
rect 6006 20961 6018 20964
rect 6052 20961 6064 20995
rect 6006 20955 6064 20961
rect 6100 20995 6158 21001
rect 6100 20961 6112 20995
rect 6146 20961 6158 20995
rect 8202 20992 8208 21004
rect 8163 20964 8208 20992
rect 6100 20955 6158 20961
rect 6115 20868 6143 20955
rect 8202 20952 8208 20964
rect 8260 20952 8266 21004
rect 10594 20992 10600 21004
rect 10555 20964 10600 20992
rect 10594 20952 10600 20964
rect 10652 20952 10658 21004
rect 10778 20992 10784 21004
rect 10739 20964 10784 20992
rect 10778 20952 10784 20964
rect 10836 20952 10842 21004
rect 11054 20992 11060 21004
rect 11015 20964 11060 20992
rect 11054 20952 11060 20964
rect 11112 20952 11118 21004
rect 11440 21001 11468 21032
rect 15212 21032 15568 21060
rect 15212 21004 15240 21032
rect 15562 21020 15568 21032
rect 15620 21020 15626 21072
rect 17512 21060 17540 21091
rect 18138 21088 18144 21100
rect 18196 21088 18202 21140
rect 16698 21032 17540 21060
rect 11425 20995 11483 21001
rect 11425 20961 11437 20995
rect 11471 20961 11483 20995
rect 15194 20992 15200 21004
rect 15155 20964 15200 20992
rect 11425 20955 11483 20961
rect 15194 20952 15200 20964
rect 15252 20952 15258 21004
rect 17494 20952 17500 21004
rect 17552 20992 17558 21004
rect 17681 20995 17739 21001
rect 17681 20992 17693 20995
rect 17552 20964 17693 20992
rect 17552 20952 17558 20964
rect 17681 20961 17693 20964
rect 17727 20992 17739 20995
rect 18325 20995 18383 21001
rect 18325 20992 18337 20995
rect 17727 20964 18337 20992
rect 17727 20961 17739 20964
rect 17681 20955 17739 20961
rect 18325 20961 18337 20964
rect 18371 20961 18383 20995
rect 20162 20992 20168 21004
rect 20123 20964 20168 20992
rect 18325 20955 18383 20961
rect 20162 20952 20168 20964
rect 20220 20952 20226 21004
rect 20901 20995 20959 21001
rect 20901 20961 20913 20995
rect 20947 20992 20959 20995
rect 21174 20992 21180 21004
rect 20947 20964 21180 20992
rect 20947 20961 20959 20964
rect 20901 20955 20959 20961
rect 21174 20952 21180 20964
rect 21232 20952 21238 21004
rect 6457 20927 6515 20933
rect 6457 20893 6469 20927
rect 6503 20924 6515 20927
rect 6546 20924 6552 20936
rect 6503 20896 6552 20924
rect 6503 20893 6515 20896
rect 6457 20887 6515 20893
rect 6546 20884 6552 20896
rect 6604 20884 6610 20936
rect 11241 20927 11299 20933
rect 11241 20893 11253 20927
rect 11287 20924 11299 20927
rect 12342 20924 12348 20936
rect 11287 20896 12348 20924
rect 11287 20893 11299 20896
rect 11241 20887 11299 20893
rect 12342 20884 12348 20896
rect 12400 20884 12406 20936
rect 15470 20924 15476 20936
rect 15431 20896 15476 20924
rect 15470 20884 15476 20896
rect 15528 20884 15534 20936
rect 6086 20816 6092 20868
rect 6144 20816 6150 20868
rect 8389 20791 8447 20797
rect 8389 20757 8401 20791
rect 8435 20788 8447 20791
rect 11790 20788 11796 20800
rect 8435 20760 11796 20788
rect 8435 20757 8447 20760
rect 8389 20751 8447 20757
rect 11790 20748 11796 20760
rect 11848 20748 11854 20800
rect 16942 20788 16948 20800
rect 16903 20760 16948 20788
rect 16942 20748 16948 20760
rect 17000 20748 17006 20800
rect 19610 20748 19616 20800
rect 19668 20788 19674 20800
rect 19981 20791 20039 20797
rect 19981 20788 19993 20791
rect 19668 20760 19993 20788
rect 19668 20748 19674 20760
rect 19981 20757 19993 20760
rect 20027 20757 20039 20791
rect 19981 20751 20039 20757
rect 20622 20748 20628 20800
rect 20680 20788 20686 20800
rect 20993 20791 21051 20797
rect 20993 20788 21005 20791
rect 20680 20760 21005 20788
rect 20680 20748 20686 20760
rect 20993 20757 21005 20760
rect 21039 20757 21051 20791
rect 20993 20751 21051 20757
rect 1104 20698 21804 20720
rect 1104 20646 4432 20698
rect 4484 20646 4496 20698
rect 4548 20646 4560 20698
rect 4612 20646 4624 20698
rect 4676 20646 11332 20698
rect 11384 20646 11396 20698
rect 11448 20646 11460 20698
rect 11512 20646 11524 20698
rect 11576 20646 18232 20698
rect 18284 20646 18296 20698
rect 18348 20646 18360 20698
rect 18412 20646 18424 20698
rect 18476 20646 21804 20698
rect 1104 20624 21804 20646
rect 13998 20584 14004 20596
rect 13959 20556 14004 20584
rect 13998 20544 14004 20556
rect 14056 20544 14062 20596
rect 21082 20584 21088 20596
rect 21043 20556 21088 20584
rect 21082 20544 21088 20556
rect 21140 20544 21146 20596
rect 6914 20516 6920 20528
rect 6875 20488 6920 20516
rect 6914 20476 6920 20488
rect 6972 20476 6978 20528
rect 10597 20519 10655 20525
rect 10597 20485 10609 20519
rect 10643 20485 10655 20519
rect 11054 20516 11060 20528
rect 10597 20479 10655 20485
rect 10796 20488 11060 20516
rect 3234 20448 3240 20460
rect 3195 20420 3240 20448
rect 3234 20408 3240 20420
rect 3292 20448 3298 20460
rect 4062 20448 4068 20460
rect 3292 20420 4068 20448
rect 3292 20408 3298 20420
rect 4062 20408 4068 20420
rect 4120 20408 4126 20460
rect 4985 20451 5043 20457
rect 4985 20417 4997 20451
rect 5031 20417 5043 20451
rect 4985 20411 5043 20417
rect 1394 20380 1400 20392
rect 1355 20352 1400 20380
rect 1394 20340 1400 20352
rect 1452 20340 1458 20392
rect 5000 20380 5028 20411
rect 6086 20408 6092 20460
rect 6144 20448 6150 20460
rect 6825 20451 6883 20457
rect 6825 20448 6837 20451
rect 6144 20420 6837 20448
rect 6144 20408 6150 20420
rect 6825 20417 6837 20420
rect 6871 20417 6883 20451
rect 8386 20448 8392 20460
rect 8347 20420 8392 20448
rect 6825 20411 6883 20417
rect 8386 20408 8392 20420
rect 8444 20408 8450 20460
rect 8665 20451 8723 20457
rect 8665 20417 8677 20451
rect 8711 20448 8723 20451
rect 10612 20448 10640 20479
rect 8711 20420 10640 20448
rect 8711 20417 8723 20420
rect 8665 20411 8723 20417
rect 5626 20380 5632 20392
rect 5000 20352 5632 20380
rect 5626 20340 5632 20352
rect 5684 20340 5690 20392
rect 7006 20380 7012 20392
rect 6967 20352 7012 20380
rect 7006 20340 7012 20352
rect 7064 20340 7070 20392
rect 7098 20340 7104 20392
rect 7156 20380 7162 20392
rect 10796 20389 10824 20488
rect 11054 20476 11060 20488
rect 11112 20516 11118 20528
rect 13909 20519 13967 20525
rect 13909 20516 13921 20519
rect 11112 20488 13921 20516
rect 11112 20476 11118 20488
rect 13909 20485 13921 20488
rect 13955 20485 13967 20519
rect 14550 20516 14556 20528
rect 13909 20479 13967 20485
rect 14200 20488 14556 20516
rect 10962 20448 10968 20460
rect 10888 20420 10968 20448
rect 10888 20389 10916 20420
rect 10962 20408 10968 20420
rect 11020 20408 11026 20460
rect 10781 20383 10839 20389
rect 7156 20352 7201 20380
rect 7156 20340 7162 20352
rect 10781 20349 10793 20383
rect 10827 20349 10839 20383
rect 10781 20343 10839 20349
rect 10873 20383 10931 20389
rect 10873 20349 10885 20383
rect 10919 20349 10931 20383
rect 11146 20380 11152 20392
rect 11107 20352 11152 20380
rect 10873 20343 10931 20349
rect 11146 20340 11152 20352
rect 11204 20340 11210 20392
rect 11238 20340 11244 20392
rect 11296 20380 11302 20392
rect 14200 20389 14228 20488
rect 14550 20476 14556 20488
rect 14608 20476 14614 20528
rect 19613 20451 19671 20457
rect 14292 20420 15056 20448
rect 14292 20389 14320 20420
rect 15028 20389 15056 20420
rect 19613 20417 19625 20451
rect 19659 20448 19671 20451
rect 19978 20448 19984 20460
rect 19659 20420 19984 20448
rect 19659 20417 19671 20420
rect 19613 20411 19671 20417
rect 19978 20408 19984 20420
rect 20036 20408 20042 20460
rect 14185 20383 14243 20389
rect 14185 20380 14197 20383
rect 11296 20352 14197 20380
rect 11296 20340 11302 20352
rect 14185 20349 14197 20352
rect 14231 20349 14243 20383
rect 14185 20343 14243 20349
rect 14277 20383 14335 20389
rect 14277 20349 14289 20383
rect 14323 20349 14335 20383
rect 14277 20343 14335 20349
rect 14553 20383 14611 20389
rect 14553 20349 14565 20383
rect 14599 20349 14611 20383
rect 14553 20343 14611 20349
rect 15013 20383 15071 20389
rect 15013 20349 15025 20383
rect 15059 20380 15071 20383
rect 15102 20380 15108 20392
rect 15059 20352 15108 20380
rect 15059 20349 15071 20352
rect 15013 20343 15071 20349
rect 3510 20312 3516 20324
rect 3471 20284 3516 20312
rect 3510 20272 3516 20284
rect 3568 20272 3574 20324
rect 4246 20272 4252 20324
rect 4304 20272 4310 20324
rect 9398 20272 9404 20324
rect 9456 20272 9462 20324
rect 10965 20315 11023 20321
rect 10965 20281 10977 20315
rect 11011 20281 11023 20315
rect 10965 20275 11023 20281
rect 14369 20315 14427 20321
rect 14369 20281 14381 20315
rect 14415 20312 14427 20315
rect 14458 20312 14464 20324
rect 14415 20284 14464 20312
rect 14415 20281 14427 20284
rect 14369 20275 14427 20281
rect 1581 20247 1639 20253
rect 1581 20213 1593 20247
rect 1627 20244 1639 20247
rect 2406 20244 2412 20256
rect 1627 20216 2412 20244
rect 1627 20213 1639 20216
rect 1581 20207 1639 20213
rect 2406 20204 2412 20216
rect 2464 20204 2470 20256
rect 5534 20244 5540 20256
rect 5495 20216 5540 20244
rect 5534 20204 5540 20216
rect 5592 20204 5598 20256
rect 10137 20247 10195 20253
rect 10137 20213 10149 20247
rect 10183 20244 10195 20247
rect 10778 20244 10784 20256
rect 10183 20216 10784 20244
rect 10183 20213 10195 20216
rect 10137 20207 10195 20213
rect 10778 20204 10784 20216
rect 10836 20244 10842 20256
rect 10980 20244 11008 20275
rect 14458 20272 14464 20284
rect 14516 20272 14522 20324
rect 14568 20312 14596 20343
rect 15102 20340 15108 20352
rect 15160 20340 15166 20392
rect 19334 20380 19340 20392
rect 19295 20352 19340 20380
rect 19334 20340 19340 20352
rect 19392 20340 19398 20392
rect 15746 20312 15752 20324
rect 14568 20284 15752 20312
rect 10836 20216 11008 20244
rect 13909 20247 13967 20253
rect 10836 20204 10842 20216
rect 13909 20213 13921 20247
rect 13955 20244 13967 20247
rect 14568 20244 14596 20284
rect 15746 20272 15752 20284
rect 15804 20272 15810 20324
rect 20622 20272 20628 20324
rect 20680 20272 20686 20324
rect 13955 20216 14596 20244
rect 13955 20213 13967 20216
rect 13909 20207 13967 20213
rect 14642 20204 14648 20256
rect 14700 20244 14706 20256
rect 15105 20247 15163 20253
rect 15105 20244 15117 20247
rect 14700 20216 15117 20244
rect 14700 20204 14706 20216
rect 15105 20213 15117 20216
rect 15151 20213 15163 20247
rect 15105 20207 15163 20213
rect 1104 20154 21804 20176
rect 1104 20102 7882 20154
rect 7934 20102 7946 20154
rect 7998 20102 8010 20154
rect 8062 20102 8074 20154
rect 8126 20102 14782 20154
rect 14834 20102 14846 20154
rect 14898 20102 14910 20154
rect 14962 20102 14974 20154
rect 15026 20102 21804 20154
rect 1104 20080 21804 20102
rect 3510 20000 3516 20052
rect 3568 20040 3574 20052
rect 4801 20043 4859 20049
rect 4801 20040 4813 20043
rect 3568 20012 4813 20040
rect 3568 20000 3574 20012
rect 4801 20009 4813 20012
rect 4847 20009 4859 20043
rect 4801 20003 4859 20009
rect 5810 20000 5816 20052
rect 5868 20040 5874 20052
rect 7561 20043 7619 20049
rect 7561 20040 7573 20043
rect 5868 20012 7573 20040
rect 5868 20000 5874 20012
rect 7561 20009 7573 20012
rect 7607 20009 7619 20043
rect 7561 20003 7619 20009
rect 9398 20000 9404 20052
rect 9456 20040 9462 20052
rect 9493 20043 9551 20049
rect 9493 20040 9505 20043
rect 9456 20012 9505 20040
rect 9456 20000 9462 20012
rect 9493 20009 9505 20012
rect 9539 20009 9551 20043
rect 9493 20003 9551 20009
rect 14458 20000 14464 20052
rect 14516 20040 14522 20052
rect 20622 20040 20628 20052
rect 14516 20012 15056 20040
rect 20583 20012 20628 20040
rect 14516 20000 14522 20012
rect 5534 19972 5540 19984
rect 5000 19944 5540 19972
rect 5000 19913 5028 19944
rect 5534 19932 5540 19944
rect 5592 19932 5598 19984
rect 6178 19972 6184 19984
rect 6091 19944 6184 19972
rect 6178 19932 6184 19944
rect 6236 19972 6242 19984
rect 15028 19981 15056 20012
rect 20622 20000 20628 20012
rect 20680 20000 20686 20052
rect 7193 19975 7251 19981
rect 7193 19972 7205 19975
rect 6236 19944 7205 19972
rect 6236 19932 6242 19944
rect 7193 19941 7205 19944
rect 7239 19941 7251 19975
rect 7193 19935 7251 19941
rect 15013 19975 15071 19981
rect 15013 19941 15025 19975
rect 15059 19941 15071 19975
rect 15013 19935 15071 19941
rect 15105 19975 15163 19981
rect 15105 19941 15117 19975
rect 15151 19972 15163 19975
rect 15194 19972 15200 19984
rect 15151 19944 15200 19972
rect 15151 19941 15163 19944
rect 15105 19935 15163 19941
rect 15194 19932 15200 19944
rect 15252 19972 15258 19984
rect 15933 19975 15991 19981
rect 15933 19972 15945 19975
rect 15252 19944 15945 19972
rect 15252 19932 15258 19944
rect 15933 19941 15945 19944
rect 15979 19941 15991 19975
rect 15933 19935 15991 19941
rect 4985 19907 5043 19913
rect 4985 19873 4997 19907
rect 5031 19873 5043 19907
rect 4985 19867 5043 19873
rect 5077 19907 5135 19913
rect 5077 19873 5089 19907
rect 5123 19904 5135 19907
rect 5353 19907 5411 19913
rect 5123 19876 5304 19904
rect 5123 19873 5135 19876
rect 5077 19867 5135 19873
rect 5276 19768 5304 19876
rect 5353 19873 5365 19907
rect 5399 19873 5411 19907
rect 6362 19904 6368 19916
rect 6323 19876 6368 19904
rect 5353 19867 5411 19873
rect 5368 19836 5396 19867
rect 6362 19864 6368 19876
rect 6420 19864 6426 19916
rect 6457 19907 6515 19913
rect 6457 19873 6469 19907
rect 6503 19904 6515 19907
rect 6638 19904 6644 19916
rect 6503 19876 6644 19904
rect 6503 19873 6515 19876
rect 6457 19867 6515 19873
rect 6638 19864 6644 19876
rect 6696 19864 6702 19916
rect 6733 19907 6791 19913
rect 6733 19873 6745 19907
rect 6779 19904 6791 19907
rect 7098 19904 7104 19916
rect 6779 19876 7104 19904
rect 6779 19873 6791 19876
rect 6733 19867 6791 19873
rect 7098 19864 7104 19876
rect 7156 19864 7162 19916
rect 7377 19907 7435 19913
rect 7377 19873 7389 19907
rect 7423 19873 7435 19907
rect 8018 19904 8024 19916
rect 7979 19876 8024 19904
rect 7377 19867 7435 19873
rect 5626 19836 5632 19848
rect 5368 19808 5632 19836
rect 5626 19796 5632 19808
rect 5684 19836 5690 19848
rect 7392 19836 7420 19867
rect 8018 19864 8024 19876
rect 8076 19864 8082 19916
rect 9677 19907 9735 19913
rect 9677 19873 9689 19907
rect 9723 19904 9735 19907
rect 9766 19904 9772 19916
rect 9723 19876 9772 19904
rect 9723 19873 9735 19876
rect 9677 19867 9735 19873
rect 9766 19864 9772 19876
rect 9824 19864 9830 19916
rect 11885 19907 11943 19913
rect 11885 19873 11897 19907
rect 11931 19904 11943 19907
rect 12434 19904 12440 19916
rect 11931 19876 12440 19904
rect 11931 19873 11943 19876
rect 11885 19867 11943 19873
rect 12434 19864 12440 19876
rect 12492 19864 12498 19916
rect 14918 19904 14924 19916
rect 14879 19876 14924 19904
rect 14918 19864 14924 19876
rect 14976 19864 14982 19916
rect 15289 19907 15347 19913
rect 15289 19873 15301 19907
rect 15335 19873 15347 19907
rect 15746 19904 15752 19916
rect 15707 19876 15752 19904
rect 15289 19867 15347 19873
rect 13170 19836 13176 19848
rect 5684 19808 7420 19836
rect 13131 19808 13176 19836
rect 5684 19796 5690 19808
rect 13170 19796 13176 19808
rect 13228 19796 13234 19848
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19805 13599 19839
rect 13541 19799 13599 19805
rect 13633 19839 13691 19845
rect 13633 19805 13645 19839
rect 13679 19836 13691 19839
rect 13814 19836 13820 19848
rect 13679 19808 13820 19836
rect 13679 19805 13691 19808
rect 13633 19799 13691 19805
rect 6546 19768 6552 19780
rect 5276 19740 6552 19768
rect 6546 19728 6552 19740
rect 6604 19768 6610 19780
rect 8018 19768 8024 19780
rect 6604 19740 8024 19768
rect 6604 19728 6610 19740
rect 8018 19728 8024 19740
rect 8076 19728 8082 19780
rect 13556 19768 13584 19799
rect 13814 19796 13820 19808
rect 13872 19796 13878 19848
rect 14182 19796 14188 19848
rect 14240 19836 14246 19848
rect 14642 19836 14648 19848
rect 14240 19808 14648 19836
rect 14240 19796 14246 19808
rect 14642 19796 14648 19808
rect 14700 19836 14706 19848
rect 15304 19836 15332 19867
rect 15746 19864 15752 19876
rect 15804 19864 15810 19916
rect 16022 19904 16028 19916
rect 15983 19876 16028 19904
rect 16022 19864 16028 19876
rect 16080 19864 16086 19916
rect 20806 19904 20812 19916
rect 20767 19876 20812 19904
rect 20806 19864 20812 19876
rect 20864 19864 20870 19916
rect 14700 19808 15332 19836
rect 14700 19796 14706 19808
rect 13722 19768 13728 19780
rect 13556 19740 13728 19768
rect 13722 19728 13728 19740
rect 13780 19768 13786 19780
rect 14737 19771 14795 19777
rect 14737 19768 14749 19771
rect 13780 19740 14749 19768
rect 13780 19728 13786 19740
rect 14737 19737 14749 19740
rect 14783 19737 14795 19771
rect 14737 19731 14795 19737
rect 15470 19728 15476 19780
rect 15528 19768 15534 19780
rect 15749 19771 15807 19777
rect 15749 19768 15761 19771
rect 15528 19740 15761 19768
rect 15528 19728 15534 19740
rect 15749 19737 15761 19740
rect 15795 19737 15807 19771
rect 15749 19731 15807 19737
rect 5261 19703 5319 19709
rect 5261 19669 5273 19703
rect 5307 19700 5319 19703
rect 5534 19700 5540 19712
rect 5307 19672 5540 19700
rect 5307 19669 5319 19672
rect 5261 19663 5319 19669
rect 5534 19660 5540 19672
rect 5592 19700 5598 19712
rect 5718 19700 5724 19712
rect 5592 19672 5724 19700
rect 5592 19660 5598 19672
rect 5718 19660 5724 19672
rect 5776 19660 5782 19712
rect 6641 19703 6699 19709
rect 6641 19669 6653 19703
rect 6687 19700 6699 19703
rect 7006 19700 7012 19712
rect 6687 19672 7012 19700
rect 6687 19669 6699 19672
rect 6641 19663 6699 19669
rect 7006 19660 7012 19672
rect 7064 19700 7070 19712
rect 7742 19700 7748 19712
rect 7064 19672 7748 19700
rect 7064 19660 7070 19672
rect 7742 19660 7748 19672
rect 7800 19660 7806 19712
rect 8113 19703 8171 19709
rect 8113 19669 8125 19703
rect 8159 19700 8171 19703
rect 8202 19700 8208 19712
rect 8159 19672 8208 19700
rect 8159 19669 8171 19672
rect 8113 19663 8171 19669
rect 8202 19660 8208 19672
rect 8260 19660 8266 19712
rect 11698 19660 11704 19712
rect 11756 19700 11762 19712
rect 11793 19703 11851 19709
rect 11793 19700 11805 19703
rect 11756 19672 11805 19700
rect 11756 19660 11762 19672
rect 11793 19669 11805 19672
rect 11839 19669 11851 19703
rect 11793 19663 11851 19669
rect 13817 19703 13875 19709
rect 13817 19669 13829 19703
rect 13863 19700 13875 19703
rect 14090 19700 14096 19712
rect 13863 19672 14096 19700
rect 13863 19669 13875 19672
rect 13817 19663 13875 19669
rect 14090 19660 14096 19672
rect 14148 19660 14154 19712
rect 1104 19610 21804 19632
rect 1104 19558 4432 19610
rect 4484 19558 4496 19610
rect 4548 19558 4560 19610
rect 4612 19558 4624 19610
rect 4676 19558 11332 19610
rect 11384 19558 11396 19610
rect 11448 19558 11460 19610
rect 11512 19558 11524 19610
rect 11576 19558 18232 19610
rect 18284 19558 18296 19610
rect 18348 19558 18360 19610
rect 18412 19558 18424 19610
rect 18476 19558 21804 19610
rect 1104 19536 21804 19558
rect 4246 19456 4252 19508
rect 4304 19496 4310 19508
rect 4433 19499 4491 19505
rect 4433 19496 4445 19499
rect 4304 19468 4445 19496
rect 4304 19456 4310 19468
rect 4433 19465 4445 19468
rect 4479 19465 4491 19499
rect 4433 19459 4491 19465
rect 5813 19499 5871 19505
rect 5813 19465 5825 19499
rect 5859 19496 5871 19499
rect 6086 19496 6092 19508
rect 5859 19468 6092 19496
rect 5859 19465 5871 19468
rect 5813 19459 5871 19465
rect 6086 19456 6092 19468
rect 6144 19456 6150 19508
rect 6917 19499 6975 19505
rect 6917 19465 6929 19499
rect 6963 19496 6975 19499
rect 7098 19496 7104 19508
rect 6963 19468 7104 19496
rect 6963 19465 6975 19468
rect 6917 19459 6975 19465
rect 7098 19456 7104 19468
rect 7156 19456 7162 19508
rect 14366 19456 14372 19508
rect 14424 19496 14430 19508
rect 15105 19499 15163 19505
rect 15105 19496 15117 19499
rect 14424 19468 15117 19496
rect 14424 19456 14430 19468
rect 15105 19465 15117 19468
rect 15151 19496 15163 19499
rect 15194 19496 15200 19508
rect 15151 19468 15200 19496
rect 15151 19465 15163 19468
rect 15105 19459 15163 19465
rect 15194 19456 15200 19468
rect 15252 19456 15258 19508
rect 16298 19456 16304 19508
rect 16356 19496 16362 19508
rect 16393 19499 16451 19505
rect 16393 19496 16405 19499
rect 16356 19468 16405 19496
rect 16356 19456 16362 19468
rect 16393 19465 16405 19468
rect 16439 19465 16451 19499
rect 16393 19459 16451 19465
rect 16114 19388 16120 19440
rect 16172 19388 16178 19440
rect 12618 19360 12624 19372
rect 12579 19332 12624 19360
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 14090 19360 14096 19372
rect 14051 19332 14096 19360
rect 14090 19320 14096 19332
rect 14148 19320 14154 19372
rect 14182 19320 14188 19372
rect 14240 19360 14246 19372
rect 14240 19332 14285 19360
rect 14240 19320 14246 19332
rect 14458 19320 14464 19372
rect 14516 19360 14522 19372
rect 15933 19363 15991 19369
rect 14516 19332 15056 19360
rect 14516 19320 14522 19332
rect 2406 19292 2412 19304
rect 2367 19264 2412 19292
rect 2406 19252 2412 19264
rect 2464 19252 2470 19304
rect 4617 19295 4675 19301
rect 4617 19261 4629 19295
rect 4663 19292 4675 19295
rect 4890 19292 4896 19304
rect 4663 19264 4896 19292
rect 4663 19261 4675 19264
rect 4617 19255 4675 19261
rect 4890 19252 4896 19264
rect 4948 19292 4954 19304
rect 5350 19292 5356 19304
rect 4948 19264 5356 19292
rect 4948 19252 4954 19264
rect 5350 19252 5356 19264
rect 5408 19252 5414 19304
rect 5626 19252 5632 19304
rect 5684 19292 5690 19304
rect 5721 19295 5779 19301
rect 5721 19292 5733 19295
rect 5684 19264 5733 19292
rect 5684 19252 5690 19264
rect 5721 19261 5733 19264
rect 5767 19261 5779 19295
rect 5721 19255 5779 19261
rect 5905 19295 5963 19301
rect 5905 19261 5917 19295
rect 5951 19292 5963 19295
rect 6178 19292 6184 19304
rect 5951 19264 6184 19292
rect 5951 19261 5963 19264
rect 5905 19255 5963 19261
rect 6178 19252 6184 19264
rect 6236 19252 6242 19304
rect 6454 19252 6460 19304
rect 6512 19292 6518 19304
rect 6825 19295 6883 19301
rect 6825 19292 6837 19295
rect 6512 19264 6837 19292
rect 6512 19252 6518 19264
rect 6825 19261 6837 19264
rect 6871 19261 6883 19295
rect 7742 19292 7748 19304
rect 7703 19264 7748 19292
rect 6825 19255 6883 19261
rect 7742 19252 7748 19264
rect 7800 19252 7806 19304
rect 8018 19252 8024 19304
rect 8076 19292 8082 19304
rect 12161 19295 12219 19301
rect 12161 19292 12173 19295
rect 8076 19264 12173 19292
rect 8076 19252 8082 19264
rect 12161 19261 12173 19264
rect 12207 19261 12219 19295
rect 12342 19292 12348 19304
rect 12303 19264 12348 19292
rect 12161 19255 12219 19261
rect 12342 19252 12348 19264
rect 12400 19252 12406 19304
rect 12434 19252 12440 19304
rect 12492 19292 12498 19304
rect 12492 19264 12585 19292
rect 12492 19252 12498 19264
rect 13170 19252 13176 19304
rect 13228 19292 13234 19304
rect 13817 19295 13875 19301
rect 13817 19292 13829 19295
rect 13228 19264 13829 19292
rect 13228 19252 13234 19264
rect 13817 19261 13829 19264
rect 13863 19261 13875 19295
rect 13817 19255 13875 19261
rect 14001 19295 14059 19301
rect 14001 19261 14013 19295
rect 14047 19292 14059 19295
rect 14274 19292 14280 19304
rect 14047 19264 14280 19292
rect 14047 19261 14059 19264
rect 14001 19255 14059 19261
rect 14274 19252 14280 19264
rect 14332 19252 14338 19304
rect 14366 19252 14372 19304
rect 14424 19292 14430 19304
rect 15028 19301 15056 19332
rect 15488 19332 15792 19360
rect 15933 19346 15945 19363
rect 15979 19346 15991 19363
rect 15013 19295 15071 19301
rect 14424 19264 14469 19292
rect 14424 19252 14430 19264
rect 15013 19261 15025 19295
rect 15059 19292 15071 19295
rect 15102 19292 15108 19304
rect 15059 19264 15108 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 15102 19252 15108 19264
rect 15160 19292 15166 19304
rect 15488 19292 15516 19332
rect 15654 19292 15660 19304
rect 15160 19264 15516 19292
rect 15615 19264 15660 19292
rect 15160 19252 15166 19264
rect 15654 19252 15660 19264
rect 15712 19252 15718 19304
rect 15764 19292 15792 19332
rect 15841 19295 15899 19301
rect 15841 19292 15853 19295
rect 15764 19264 15853 19292
rect 15841 19261 15853 19264
rect 15887 19261 15899 19295
rect 15930 19294 15936 19346
rect 15988 19294 15994 19346
rect 16025 19295 16083 19301
rect 15841 19255 15899 19261
rect 16025 19261 16037 19295
rect 16071 19292 16083 19295
rect 16132 19292 16160 19388
rect 17678 19360 17684 19372
rect 16316 19332 16712 19360
rect 17639 19332 17684 19360
rect 16071 19264 16160 19292
rect 16209 19295 16267 19301
rect 16071 19261 16083 19264
rect 16025 19255 16083 19261
rect 16209 19261 16221 19295
rect 16255 19292 16267 19295
rect 16316 19292 16344 19332
rect 16255 19264 16344 19292
rect 16684 19292 16712 19332
rect 17678 19320 17684 19332
rect 17736 19320 17742 19372
rect 17586 19292 17592 19304
rect 16684 19264 17592 19292
rect 16255 19261 16267 19264
rect 16209 19255 16267 19261
rect 17586 19252 17592 19264
rect 17644 19252 17650 19304
rect 17862 19292 17868 19304
rect 17823 19264 17868 19292
rect 17862 19252 17868 19264
rect 17920 19252 17926 19304
rect 17954 19252 17960 19304
rect 18012 19292 18018 19304
rect 18509 19295 18567 19301
rect 18509 19292 18521 19295
rect 18012 19264 18057 19292
rect 18156 19264 18521 19292
rect 18012 19252 18018 19264
rect 6638 19184 6644 19236
rect 6696 19224 6702 19236
rect 7837 19227 7895 19233
rect 7837 19224 7849 19227
rect 6696 19196 7849 19224
rect 6696 19184 6702 19196
rect 7837 19193 7849 19196
rect 7883 19193 7895 19227
rect 7837 19187 7895 19193
rect 2590 19156 2596 19168
rect 2551 19128 2596 19156
rect 2590 19116 2596 19128
rect 2648 19116 2654 19168
rect 7650 19116 7656 19168
rect 7708 19156 7714 19168
rect 8036 19156 8064 19252
rect 7708 19128 8064 19156
rect 12452 19156 12480 19252
rect 12710 19224 12716 19236
rect 12671 19196 12716 19224
rect 12710 19184 12716 19196
rect 12768 19184 12774 19236
rect 12802 19184 12808 19236
rect 12860 19224 12866 19236
rect 12860 19196 12905 19224
rect 12860 19184 12866 19196
rect 12986 19184 12992 19236
rect 13044 19224 13050 19236
rect 17681 19227 17739 19233
rect 17681 19224 17693 19227
rect 13044 19196 17693 19224
rect 13044 19184 13050 19196
rect 17681 19193 17693 19196
rect 17727 19193 17739 19227
rect 17681 19187 17739 19193
rect 14553 19159 14611 19165
rect 14553 19156 14565 19159
rect 12452 19128 14565 19156
rect 7708 19116 7714 19128
rect 14553 19125 14565 19128
rect 14599 19125 14611 19159
rect 14553 19119 14611 19125
rect 15654 19116 15660 19168
rect 15712 19156 15718 19168
rect 18156 19156 18184 19264
rect 18509 19261 18521 19264
rect 18555 19261 18567 19295
rect 18509 19255 18567 19261
rect 18524 19224 18552 19255
rect 19150 19252 19156 19304
rect 19208 19292 19214 19304
rect 19429 19295 19487 19301
rect 19429 19292 19441 19295
rect 19208 19264 19441 19292
rect 19208 19252 19214 19264
rect 19429 19261 19441 19264
rect 19475 19261 19487 19295
rect 19610 19292 19616 19304
rect 19571 19264 19616 19292
rect 19429 19255 19487 19261
rect 19610 19252 19616 19264
rect 19668 19252 19674 19304
rect 19886 19224 19892 19236
rect 18524 19196 19892 19224
rect 19886 19184 19892 19196
rect 19944 19224 19950 19236
rect 20438 19224 20444 19236
rect 19944 19196 20444 19224
rect 19944 19184 19950 19196
rect 20438 19184 20444 19196
rect 20496 19184 20502 19236
rect 18598 19156 18604 19168
rect 15712 19128 18184 19156
rect 18559 19128 18604 19156
rect 15712 19116 15718 19128
rect 18598 19116 18604 19128
rect 18656 19116 18662 19168
rect 19518 19156 19524 19168
rect 19479 19128 19524 19156
rect 19518 19116 19524 19128
rect 19576 19116 19582 19168
rect 1104 19066 21804 19088
rect 1104 19014 7882 19066
rect 7934 19014 7946 19066
rect 7998 19014 8010 19066
rect 8062 19014 8074 19066
rect 8126 19014 14782 19066
rect 14834 19014 14846 19066
rect 14898 19014 14910 19066
rect 14962 19014 14974 19066
rect 15026 19014 21804 19066
rect 1104 18992 21804 19014
rect 12710 18912 12716 18964
rect 12768 18952 12774 18964
rect 12768 18924 13124 18952
rect 12768 18912 12774 18924
rect 5813 18887 5871 18893
rect 5813 18853 5825 18887
rect 5859 18884 5871 18887
rect 12802 18884 12808 18896
rect 5859 18856 6500 18884
rect 5859 18853 5871 18856
rect 5813 18847 5871 18853
rect 5994 18816 6000 18828
rect 5955 18788 6000 18816
rect 5994 18776 6000 18788
rect 6052 18776 6058 18828
rect 6472 18825 6500 18856
rect 11808 18856 12808 18884
rect 6457 18819 6515 18825
rect 6457 18785 6469 18819
rect 6503 18816 6515 18819
rect 6914 18816 6920 18828
rect 6503 18788 6920 18816
rect 6503 18785 6515 18788
rect 6457 18779 6515 18785
rect 6914 18776 6920 18788
rect 6972 18776 6978 18828
rect 7374 18816 7380 18828
rect 7335 18788 7380 18816
rect 7374 18776 7380 18788
rect 7432 18776 7438 18828
rect 7558 18776 7564 18828
rect 7616 18816 7622 18828
rect 7837 18819 7895 18825
rect 7837 18816 7849 18819
rect 7616 18788 7849 18816
rect 7616 18776 7622 18788
rect 7837 18785 7849 18788
rect 7883 18785 7895 18819
rect 11698 18816 11704 18828
rect 11659 18788 11704 18816
rect 7837 18779 7895 18785
rect 11698 18776 11704 18788
rect 11756 18776 11762 18828
rect 11808 18825 11836 18856
rect 12802 18844 12808 18856
rect 12860 18844 12866 18896
rect 13096 18884 13124 18924
rect 13170 18912 13176 18964
rect 13228 18952 13234 18964
rect 13449 18955 13507 18961
rect 13449 18952 13461 18955
rect 13228 18924 13461 18952
rect 13228 18912 13234 18924
rect 13449 18921 13461 18924
rect 13495 18921 13507 18955
rect 18877 18955 18935 18961
rect 18877 18952 18889 18955
rect 13449 18915 13507 18921
rect 13556 18924 18889 18952
rect 13556 18884 13584 18924
rect 18877 18921 18889 18924
rect 18923 18921 18935 18955
rect 18877 18915 18935 18921
rect 13096 18856 13584 18884
rect 13633 18887 13691 18893
rect 13633 18853 13645 18887
rect 13679 18884 13691 18887
rect 13722 18884 13728 18896
rect 13679 18856 13728 18884
rect 13679 18853 13691 18856
rect 13633 18847 13691 18853
rect 13722 18844 13728 18856
rect 13780 18844 13786 18896
rect 16209 18887 16267 18893
rect 16209 18853 16221 18887
rect 16255 18884 16267 18887
rect 16298 18884 16304 18896
rect 16255 18856 16304 18884
rect 16255 18853 16267 18856
rect 16209 18847 16267 18853
rect 16298 18844 16304 18856
rect 16356 18844 16362 18896
rect 18969 18887 19027 18893
rect 18969 18853 18981 18887
rect 19015 18884 19027 18887
rect 20714 18884 20720 18896
rect 19015 18856 20720 18884
rect 19015 18853 19027 18856
rect 18969 18847 19027 18853
rect 20714 18844 20720 18856
rect 20772 18844 20778 18896
rect 11793 18819 11851 18825
rect 11793 18785 11805 18819
rect 11839 18785 11851 18819
rect 11974 18816 11980 18828
rect 11935 18788 11980 18816
rect 11793 18779 11851 18785
rect 11974 18776 11980 18788
rect 12032 18776 12038 18828
rect 12250 18816 12256 18828
rect 12211 18788 12256 18816
rect 12250 18776 12256 18788
rect 12308 18776 12314 18828
rect 12529 18819 12587 18825
rect 12529 18785 12541 18819
rect 12575 18816 12587 18819
rect 12986 18816 12992 18828
rect 12575 18788 12992 18816
rect 12575 18785 12587 18788
rect 12529 18779 12587 18785
rect 12986 18776 12992 18788
rect 13044 18776 13050 18828
rect 13814 18816 13820 18828
rect 13775 18788 13820 18816
rect 13814 18776 13820 18788
rect 13872 18776 13878 18828
rect 17310 18776 17316 18828
rect 17368 18776 17374 18828
rect 17862 18776 17868 18828
rect 17920 18816 17926 18828
rect 18601 18819 18659 18825
rect 18601 18816 18613 18819
rect 17920 18788 18613 18816
rect 17920 18776 17926 18788
rect 18601 18785 18613 18788
rect 18647 18816 18659 18819
rect 18782 18816 18788 18828
rect 18647 18788 18788 18816
rect 18647 18785 18659 18788
rect 18601 18779 18659 18785
rect 18782 18776 18788 18788
rect 18840 18776 18846 18828
rect 19058 18816 19064 18828
rect 19019 18788 19064 18816
rect 19058 18776 19064 18788
rect 19116 18776 19122 18828
rect 7742 18708 7748 18760
rect 7800 18748 7806 18760
rect 8110 18748 8116 18760
rect 7800 18720 8116 18748
rect 7800 18708 7806 18720
rect 8110 18708 8116 18720
rect 8168 18748 8174 18760
rect 11149 18751 11207 18757
rect 11149 18748 11161 18751
rect 8168 18720 11161 18748
rect 8168 18708 8174 18720
rect 11149 18717 11161 18720
rect 11195 18717 11207 18751
rect 11149 18711 11207 18717
rect 15562 18708 15568 18760
rect 15620 18748 15626 18760
rect 15933 18751 15991 18757
rect 15933 18748 15945 18751
rect 15620 18720 15945 18748
rect 15620 18708 15626 18720
rect 15933 18717 15945 18720
rect 15979 18717 15991 18751
rect 15933 18711 15991 18717
rect 5350 18572 5356 18624
rect 5408 18612 5414 18624
rect 5629 18615 5687 18621
rect 5629 18612 5641 18615
rect 5408 18584 5641 18612
rect 5408 18572 5414 18584
rect 5629 18581 5641 18584
rect 5675 18581 5687 18615
rect 5629 18575 5687 18581
rect 6549 18615 6607 18621
rect 6549 18581 6561 18615
rect 6595 18612 6607 18615
rect 7006 18612 7012 18624
rect 6595 18584 7012 18612
rect 6595 18581 6607 18584
rect 6549 18575 6607 18581
rect 7006 18572 7012 18584
rect 7064 18572 7070 18624
rect 7285 18615 7343 18621
rect 7285 18581 7297 18615
rect 7331 18612 7343 18615
rect 7742 18612 7748 18624
rect 7331 18584 7748 18612
rect 7331 18581 7343 18584
rect 7285 18575 7343 18581
rect 7742 18572 7748 18584
rect 7800 18572 7806 18624
rect 7929 18615 7987 18621
rect 7929 18581 7941 18615
rect 7975 18612 7987 18615
rect 8202 18612 8208 18624
rect 7975 18584 8208 18612
rect 7975 18581 7987 18584
rect 7929 18575 7987 18581
rect 8202 18572 8208 18584
rect 8260 18572 8266 18624
rect 15102 18572 15108 18624
rect 15160 18612 15166 18624
rect 16942 18612 16948 18624
rect 15160 18584 16948 18612
rect 15160 18572 15166 18584
rect 16942 18572 16948 18584
rect 17000 18612 17006 18624
rect 17402 18612 17408 18624
rect 17000 18584 17408 18612
rect 17000 18572 17006 18584
rect 17402 18572 17408 18584
rect 17460 18572 17466 18624
rect 17678 18612 17684 18624
rect 17639 18584 17684 18612
rect 17678 18572 17684 18584
rect 17736 18572 17742 18624
rect 1104 18522 21804 18544
rect 1104 18470 4432 18522
rect 4484 18470 4496 18522
rect 4548 18470 4560 18522
rect 4612 18470 4624 18522
rect 4676 18470 11332 18522
rect 11384 18470 11396 18522
rect 11448 18470 11460 18522
rect 11512 18470 11524 18522
rect 11576 18470 18232 18522
rect 18284 18470 18296 18522
rect 18348 18470 18360 18522
rect 18412 18470 18424 18522
rect 18476 18470 21804 18522
rect 1104 18448 21804 18470
rect 6638 18368 6644 18420
rect 6696 18408 6702 18420
rect 8297 18411 8355 18417
rect 8297 18408 8309 18411
rect 6696 18380 8309 18408
rect 6696 18368 6702 18380
rect 8297 18377 8309 18380
rect 8343 18377 8355 18411
rect 12066 18408 12072 18420
rect 12027 18380 12072 18408
rect 8297 18371 8355 18377
rect 12066 18368 12072 18380
rect 12124 18368 12130 18420
rect 12250 18368 12256 18420
rect 12308 18408 12314 18420
rect 12437 18411 12495 18417
rect 12437 18408 12449 18411
rect 12308 18380 12449 18408
rect 12308 18368 12314 18380
rect 12437 18377 12449 18380
rect 12483 18377 12495 18411
rect 12437 18371 12495 18377
rect 12802 18368 12808 18420
rect 12860 18408 12866 18420
rect 13817 18411 13875 18417
rect 13817 18408 13829 18411
rect 12860 18380 13829 18408
rect 12860 18368 12866 18380
rect 13817 18377 13829 18380
rect 13863 18377 13875 18411
rect 13817 18371 13875 18377
rect 16022 18368 16028 18420
rect 16080 18408 16086 18420
rect 16301 18411 16359 18417
rect 16301 18408 16313 18411
rect 16080 18380 16313 18408
rect 16080 18368 16086 18380
rect 16301 18377 16313 18380
rect 16347 18377 16359 18411
rect 17310 18408 17316 18420
rect 17271 18380 17316 18408
rect 16301 18371 16359 18377
rect 17310 18368 17316 18380
rect 17368 18368 17374 18420
rect 17954 18368 17960 18420
rect 18012 18408 18018 18420
rect 18233 18411 18291 18417
rect 18233 18408 18245 18411
rect 18012 18380 18245 18408
rect 18012 18368 18018 18380
rect 18233 18377 18245 18380
rect 18279 18377 18291 18411
rect 18782 18408 18788 18420
rect 18743 18380 18788 18408
rect 18233 18371 18291 18377
rect 18782 18368 18788 18380
rect 18840 18368 18846 18420
rect 6178 18340 6184 18352
rect 5460 18312 6184 18340
rect 4525 18207 4583 18213
rect 4525 18173 4537 18207
rect 4571 18204 4583 18207
rect 4890 18204 4896 18216
rect 4571 18176 4896 18204
rect 4571 18173 4583 18176
rect 4525 18167 4583 18173
rect 4890 18164 4896 18176
rect 4948 18164 4954 18216
rect 5350 18204 5356 18216
rect 5311 18176 5356 18204
rect 5350 18164 5356 18176
rect 5408 18164 5414 18216
rect 5460 18213 5488 18312
rect 6178 18300 6184 18312
rect 6236 18300 6242 18352
rect 6273 18343 6331 18349
rect 6273 18309 6285 18343
rect 6319 18340 6331 18343
rect 7650 18340 7656 18352
rect 6319 18312 7656 18340
rect 6319 18309 6331 18312
rect 6273 18303 6331 18309
rect 7650 18300 7656 18312
rect 7708 18300 7714 18352
rect 12084 18340 12112 18368
rect 12989 18343 13047 18349
rect 12989 18340 13001 18343
rect 8312 18312 9076 18340
rect 12084 18312 13001 18340
rect 8312 18284 8340 18312
rect 8294 18272 8300 18284
rect 5736 18244 8300 18272
rect 5445 18207 5503 18213
rect 5445 18173 5457 18207
rect 5491 18173 5503 18207
rect 5736 18204 5764 18244
rect 8294 18232 8300 18244
rect 8352 18232 8358 18284
rect 8846 18272 8852 18284
rect 8807 18244 8852 18272
rect 8846 18232 8852 18244
rect 8904 18232 8910 18284
rect 9048 18281 9076 18312
rect 12989 18309 13001 18312
rect 13035 18309 13047 18343
rect 12989 18303 13047 18309
rect 19239 18300 19245 18352
rect 19297 18340 19303 18352
rect 19518 18340 19524 18352
rect 19297 18312 19524 18340
rect 19297 18300 19303 18312
rect 19518 18300 19524 18312
rect 19576 18300 19582 18352
rect 9033 18275 9091 18281
rect 9033 18241 9045 18275
rect 9079 18272 9091 18275
rect 9582 18272 9588 18284
rect 9079 18244 9588 18272
rect 9079 18241 9091 18244
rect 9033 18235 9091 18241
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 11057 18275 11115 18281
rect 11057 18241 11069 18275
rect 11103 18272 11115 18275
rect 11974 18272 11980 18284
rect 11103 18244 11980 18272
rect 11103 18241 11115 18244
rect 11057 18235 11115 18241
rect 11974 18232 11980 18244
rect 12032 18272 12038 18284
rect 12161 18275 12219 18281
rect 12161 18272 12173 18275
rect 12032 18244 12173 18272
rect 12032 18232 12038 18244
rect 12161 18241 12173 18244
rect 12207 18241 12219 18275
rect 14090 18272 14096 18284
rect 12161 18235 12219 18241
rect 13740 18244 14096 18272
rect 5445 18167 5503 18173
rect 5598 18176 5764 18204
rect 5813 18207 5871 18213
rect 5598 18148 5626 18176
rect 5813 18173 5825 18207
rect 5859 18204 5871 18207
rect 6273 18207 6331 18213
rect 6273 18204 6285 18207
rect 5859 18176 6285 18204
rect 5859 18173 5871 18176
rect 5813 18167 5871 18173
rect 6273 18173 6285 18176
rect 6319 18173 6331 18207
rect 7006 18204 7012 18216
rect 6967 18176 7012 18204
rect 6273 18167 6331 18173
rect 7006 18164 7012 18176
rect 7064 18164 7070 18216
rect 8021 18207 8079 18213
rect 8021 18173 8033 18207
rect 8067 18173 8079 18207
rect 8021 18167 8079 18173
rect 4614 18096 4620 18148
rect 4672 18136 4678 18148
rect 5169 18139 5227 18145
rect 5169 18136 5181 18139
rect 4672 18108 5181 18136
rect 4672 18096 4678 18108
rect 5169 18105 5181 18108
rect 5215 18105 5227 18139
rect 5534 18136 5540 18148
rect 5447 18108 5540 18136
rect 5169 18099 5227 18105
rect 5534 18096 5540 18108
rect 5592 18108 5626 18148
rect 5675 18139 5733 18145
rect 5592 18096 5598 18108
rect 5675 18105 5687 18139
rect 5721 18136 5733 18139
rect 6086 18136 6092 18148
rect 5721 18108 6092 18136
rect 5721 18105 5733 18108
rect 5675 18099 5733 18105
rect 6086 18096 6092 18108
rect 6144 18096 6150 18148
rect 6730 18096 6736 18148
rect 6788 18136 6794 18148
rect 6825 18139 6883 18145
rect 6825 18136 6837 18139
rect 6788 18108 6837 18136
rect 6788 18096 6794 18108
rect 6825 18105 6837 18108
rect 6871 18105 6883 18139
rect 6825 18099 6883 18105
rect 4709 18071 4767 18077
rect 4709 18037 4721 18071
rect 4755 18068 4767 18071
rect 4982 18068 4988 18080
rect 4755 18040 4988 18068
rect 4755 18037 4767 18040
rect 4709 18031 4767 18037
rect 4982 18028 4988 18040
rect 5040 18028 5046 18080
rect 6178 18028 6184 18080
rect 6236 18068 6242 18080
rect 7193 18071 7251 18077
rect 7193 18068 7205 18071
rect 6236 18040 7205 18068
rect 6236 18028 6242 18040
rect 7193 18037 7205 18040
rect 7239 18068 7251 18071
rect 7282 18068 7288 18080
rect 7239 18040 7288 18068
rect 7239 18037 7251 18040
rect 7193 18031 7251 18037
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 7558 18028 7564 18080
rect 7616 18068 7622 18080
rect 7837 18071 7895 18077
rect 7837 18068 7849 18071
rect 7616 18040 7849 18068
rect 7616 18028 7622 18040
rect 7837 18037 7849 18040
rect 7883 18037 7895 18071
rect 8036 18068 8064 18167
rect 8110 18164 8116 18216
rect 8168 18204 8174 18216
rect 8386 18204 8392 18216
rect 8168 18176 8213 18204
rect 8347 18176 8392 18204
rect 8168 18164 8174 18176
rect 8386 18164 8392 18176
rect 8444 18164 8450 18216
rect 9125 18207 9183 18213
rect 9125 18173 9137 18207
rect 9171 18173 9183 18207
rect 9125 18167 9183 18173
rect 8128 18136 8156 18164
rect 8294 18136 8300 18148
rect 8128 18108 8300 18136
rect 8294 18096 8300 18108
rect 8352 18096 8358 18148
rect 8404 18136 8432 18164
rect 9140 18136 9168 18167
rect 9766 18164 9772 18216
rect 9824 18204 9830 18216
rect 9861 18207 9919 18213
rect 9861 18204 9873 18207
rect 9824 18176 9873 18204
rect 9824 18164 9830 18176
rect 9861 18173 9873 18176
rect 9907 18204 9919 18207
rect 10502 18204 10508 18216
rect 9907 18176 10508 18204
rect 9907 18173 9919 18176
rect 9861 18167 9919 18173
rect 10502 18164 10508 18176
rect 10560 18164 10566 18216
rect 10965 18207 11023 18213
rect 10965 18173 10977 18207
rect 11011 18204 11023 18207
rect 11790 18204 11796 18216
rect 11011 18176 11796 18204
rect 11011 18173 11023 18176
rect 10965 18167 11023 18173
rect 11790 18164 11796 18176
rect 11848 18164 11854 18216
rect 13740 18213 13768 18244
rect 14090 18232 14096 18244
rect 14148 18232 14154 18284
rect 17678 18272 17684 18284
rect 16224 18244 17684 18272
rect 16224 18216 16252 18244
rect 17678 18232 17684 18244
rect 17736 18232 17742 18284
rect 19610 18272 19616 18284
rect 18984 18244 19616 18272
rect 12069 18207 12127 18213
rect 12069 18173 12081 18207
rect 12115 18204 12127 18207
rect 13081 18207 13139 18213
rect 12115 18176 12204 18204
rect 12115 18173 12127 18176
rect 12069 18167 12127 18173
rect 12176 18148 12204 18176
rect 13081 18173 13093 18207
rect 13127 18173 13139 18207
rect 13081 18167 13139 18173
rect 13725 18207 13783 18213
rect 13725 18173 13737 18207
rect 13771 18173 13783 18207
rect 13725 18167 13783 18173
rect 13909 18207 13967 18213
rect 13909 18173 13921 18207
rect 13955 18204 13967 18207
rect 14274 18204 14280 18216
rect 13955 18176 14280 18204
rect 13955 18173 13967 18176
rect 13909 18167 13967 18173
rect 8404 18108 9168 18136
rect 12158 18096 12164 18148
rect 12216 18096 12222 18148
rect 13096 18136 13124 18167
rect 14274 18164 14280 18176
rect 14332 18164 14338 18216
rect 16206 18204 16212 18216
rect 16119 18176 16212 18204
rect 16206 18164 16212 18176
rect 16264 18164 16270 18216
rect 16393 18207 16451 18213
rect 16393 18173 16405 18207
rect 16439 18173 16451 18207
rect 17494 18204 17500 18216
rect 17455 18176 17500 18204
rect 16393 18167 16451 18173
rect 14090 18136 14096 18148
rect 13096 18108 14096 18136
rect 14090 18096 14096 18108
rect 14148 18096 14154 18148
rect 16114 18096 16120 18148
rect 16172 18136 16178 18148
rect 16408 18136 16436 18167
rect 17494 18164 17500 18176
rect 17552 18164 17558 18216
rect 18984 18213 19012 18244
rect 19610 18232 19616 18244
rect 19668 18232 19674 18284
rect 18325 18207 18383 18213
rect 18325 18173 18337 18207
rect 18371 18173 18383 18207
rect 18325 18167 18383 18173
rect 18969 18207 19027 18213
rect 18969 18173 18981 18207
rect 19015 18173 19027 18207
rect 19150 18204 19156 18216
rect 19111 18176 19156 18204
rect 18969 18167 19027 18173
rect 17586 18136 17592 18148
rect 16172 18108 17592 18136
rect 16172 18096 16178 18108
rect 17586 18096 17592 18108
rect 17644 18096 17650 18148
rect 8662 18068 8668 18080
rect 8036 18040 8668 18068
rect 7837 18031 7895 18037
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 8849 18071 8907 18077
rect 8849 18037 8861 18071
rect 8895 18068 8907 18071
rect 9766 18068 9772 18080
rect 8895 18040 9772 18068
rect 8895 18037 8907 18040
rect 8849 18031 8907 18037
rect 9766 18028 9772 18040
rect 9824 18028 9830 18080
rect 10042 18068 10048 18080
rect 10003 18040 10048 18068
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 18340 18068 18368 18167
rect 19150 18164 19156 18176
rect 19208 18164 19214 18216
rect 19245 18207 19303 18213
rect 19245 18173 19257 18207
rect 19291 18173 19303 18207
rect 19245 18167 19303 18173
rect 19337 18207 19395 18213
rect 19337 18173 19349 18207
rect 19383 18173 19395 18207
rect 19518 18204 19524 18216
rect 19479 18176 19524 18204
rect 19337 18167 19395 18173
rect 19058 18096 19064 18148
rect 19116 18136 19122 18148
rect 19260 18136 19288 18167
rect 19116 18108 19288 18136
rect 19116 18096 19122 18108
rect 19242 18068 19248 18080
rect 18340 18040 19248 18068
rect 19242 18028 19248 18040
rect 19300 18028 19306 18080
rect 19352 18068 19380 18167
rect 19518 18164 19524 18176
rect 19576 18164 19582 18216
rect 20622 18164 20628 18216
rect 20680 18204 20686 18216
rect 21085 18207 21143 18213
rect 21085 18204 21097 18207
rect 20680 18176 21097 18204
rect 20680 18164 20686 18176
rect 21085 18173 21097 18176
rect 21131 18173 21143 18207
rect 21085 18167 21143 18173
rect 20714 18068 20720 18080
rect 19352 18040 20720 18068
rect 20714 18028 20720 18040
rect 20772 18028 20778 18080
rect 20806 18028 20812 18080
rect 20864 18068 20870 18080
rect 20901 18071 20959 18077
rect 20901 18068 20913 18071
rect 20864 18040 20913 18068
rect 20864 18028 20870 18040
rect 20901 18037 20913 18040
rect 20947 18037 20959 18071
rect 20901 18031 20959 18037
rect 1104 17978 21804 18000
rect 1104 17926 7882 17978
rect 7934 17926 7946 17978
rect 7998 17926 8010 17978
rect 8062 17926 8074 17978
rect 8126 17926 14782 17978
rect 14834 17926 14846 17978
rect 14898 17926 14910 17978
rect 14962 17926 14974 17978
rect 15026 17926 21804 17978
rect 1104 17904 21804 17926
rect 5994 17824 6000 17876
rect 6052 17864 6058 17876
rect 6549 17867 6607 17873
rect 6549 17864 6561 17867
rect 6052 17836 6561 17864
rect 6052 17824 6058 17836
rect 6549 17833 6561 17836
rect 6595 17833 6607 17867
rect 8202 17864 8208 17876
rect 6549 17827 6607 17833
rect 8036 17836 8208 17864
rect 4525 17799 4583 17805
rect 4525 17765 4537 17799
rect 4571 17796 4583 17799
rect 4614 17796 4620 17808
rect 4571 17768 4620 17796
rect 4571 17765 4583 17768
rect 4525 17759 4583 17765
rect 4614 17756 4620 17768
rect 4672 17756 4678 17808
rect 4982 17756 4988 17808
rect 5040 17756 5046 17808
rect 6638 17756 6644 17808
rect 6696 17796 6702 17808
rect 6696 17768 6868 17796
rect 6696 17756 6702 17768
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 4154 17688 4160 17740
rect 4212 17728 4218 17740
rect 4249 17731 4307 17737
rect 4249 17728 4261 17731
rect 4212 17700 4261 17728
rect 4212 17688 4218 17700
rect 4249 17697 4261 17700
rect 4295 17697 4307 17731
rect 4249 17691 4307 17697
rect 6086 17688 6092 17740
rect 6144 17728 6150 17740
rect 6840 17737 6868 17768
rect 7190 17756 7196 17808
rect 7248 17796 7254 17808
rect 7558 17796 7564 17808
rect 7248 17768 7564 17796
rect 7248 17756 7254 17768
rect 7558 17756 7564 17768
rect 7616 17796 7622 17808
rect 8036 17805 8064 17836
rect 8202 17824 8208 17836
rect 8260 17824 8266 17876
rect 8297 17867 8355 17873
rect 8297 17833 8309 17867
rect 8343 17864 8355 17867
rect 8846 17864 8852 17876
rect 8343 17836 8852 17864
rect 8343 17833 8355 17836
rect 8297 17827 8355 17833
rect 8846 17824 8852 17836
rect 8904 17824 8910 17876
rect 12618 17824 12624 17876
rect 12676 17864 12682 17876
rect 12713 17867 12771 17873
rect 12713 17864 12725 17867
rect 12676 17836 12725 17864
rect 12676 17824 12682 17836
rect 12713 17833 12725 17836
rect 12759 17833 12771 17867
rect 12713 17827 12771 17833
rect 13906 17824 13912 17876
rect 13964 17864 13970 17876
rect 15197 17867 15255 17873
rect 15197 17864 15209 17867
rect 13964 17836 15209 17864
rect 13964 17824 13970 17836
rect 15197 17833 15209 17836
rect 15243 17833 15255 17867
rect 15197 17827 15255 17833
rect 15381 17867 15439 17873
rect 15381 17833 15393 17867
rect 15427 17833 15439 17867
rect 15381 17827 15439 17833
rect 7929 17799 7987 17805
rect 7929 17796 7941 17799
rect 7616 17768 7941 17796
rect 7616 17756 7622 17768
rect 7929 17765 7941 17768
rect 7975 17765 7987 17799
rect 7929 17759 7987 17765
rect 8021 17799 8079 17805
rect 8021 17765 8033 17799
rect 8067 17765 8079 17799
rect 9766 17796 9772 17808
rect 9727 17768 9772 17796
rect 8021 17759 8079 17765
rect 9766 17756 9772 17768
rect 9824 17756 9830 17808
rect 10042 17756 10048 17808
rect 10100 17796 10106 17808
rect 10100 17768 10258 17796
rect 10100 17756 10106 17768
rect 11790 17756 11796 17808
rect 11848 17796 11854 17808
rect 11848 17768 12112 17796
rect 11848 17756 11854 17768
rect 6733 17731 6791 17737
rect 6733 17728 6745 17731
rect 6144 17700 6745 17728
rect 6144 17688 6150 17700
rect 6733 17697 6745 17700
rect 6779 17697 6791 17731
rect 6733 17691 6791 17697
rect 6825 17731 6883 17737
rect 6825 17697 6837 17731
rect 6871 17697 6883 17731
rect 6825 17691 6883 17697
rect 7101 17731 7159 17737
rect 7101 17697 7113 17731
rect 7147 17697 7159 17731
rect 7650 17728 7656 17740
rect 7101 17691 7159 17697
rect 7208 17700 7656 17728
rect 7116 17592 7144 17691
rect 7208 17672 7236 17700
rect 7650 17688 7656 17700
rect 7708 17688 7714 17740
rect 7742 17688 7748 17740
rect 7800 17728 7806 17740
rect 8118 17731 8176 17737
rect 8118 17728 8130 17731
rect 7800 17700 7845 17728
rect 7944 17700 8130 17728
rect 7800 17688 7806 17700
rect 7190 17620 7196 17672
rect 7248 17620 7254 17672
rect 7374 17620 7380 17672
rect 7432 17660 7438 17672
rect 7944 17660 7972 17700
rect 8118 17697 8130 17700
rect 8164 17697 8176 17731
rect 8118 17691 8176 17697
rect 8478 17688 8484 17740
rect 8536 17728 8542 17740
rect 9490 17728 9496 17740
rect 8536 17700 9496 17728
rect 8536 17688 8542 17700
rect 9490 17688 9496 17700
rect 9548 17688 9554 17740
rect 11974 17728 11980 17740
rect 11935 17700 11980 17728
rect 11974 17688 11980 17700
rect 12032 17688 12038 17740
rect 12084 17728 12112 17768
rect 12158 17756 12164 17808
rect 12216 17796 12222 17808
rect 12216 17768 12848 17796
rect 12216 17756 12222 17768
rect 12820 17737 12848 17768
rect 13814 17756 13820 17808
rect 13872 17796 13878 17808
rect 15396 17796 15424 17827
rect 13872 17768 15424 17796
rect 19076 17768 20300 17796
rect 13872 17756 13878 17768
rect 12345 17731 12403 17737
rect 12345 17728 12357 17731
rect 12084 17700 12357 17728
rect 12345 17697 12357 17700
rect 12391 17697 12403 17731
rect 12345 17691 12403 17697
rect 12805 17731 12863 17737
rect 12805 17697 12817 17731
rect 12851 17697 12863 17731
rect 12805 17691 12863 17697
rect 13630 17688 13636 17740
rect 13688 17728 13694 17740
rect 15256 17731 15314 17737
rect 15256 17728 15268 17731
rect 13688 17700 15268 17728
rect 13688 17688 13694 17700
rect 15256 17697 15268 17700
rect 15302 17728 15314 17731
rect 16206 17728 16212 17740
rect 15302 17700 16212 17728
rect 15302 17697 15314 17700
rect 15256 17691 15314 17697
rect 16206 17688 16212 17700
rect 16264 17688 16270 17740
rect 16390 17688 16396 17740
rect 16448 17728 16454 17740
rect 17494 17728 17500 17740
rect 16448 17700 17500 17728
rect 16448 17688 16454 17700
rect 17494 17688 17500 17700
rect 17552 17728 17558 17740
rect 19076 17737 19104 17768
rect 20272 17740 20300 17768
rect 17589 17731 17647 17737
rect 17589 17728 17601 17731
rect 17552 17700 17601 17728
rect 17552 17688 17558 17700
rect 17589 17697 17601 17700
rect 17635 17697 17647 17731
rect 17589 17691 17647 17697
rect 19061 17731 19119 17737
rect 19061 17697 19073 17731
rect 19107 17697 19119 17731
rect 19061 17691 19119 17697
rect 19334 17688 19340 17740
rect 19392 17728 19398 17740
rect 19981 17731 20039 17737
rect 19981 17728 19993 17731
rect 19392 17700 19993 17728
rect 19392 17688 19398 17700
rect 19981 17697 19993 17700
rect 20027 17697 20039 17731
rect 19981 17691 20039 17697
rect 20165 17731 20223 17737
rect 20165 17697 20177 17731
rect 20211 17697 20223 17731
rect 20165 17691 20223 17697
rect 8018 17660 8024 17672
rect 7432 17632 8024 17660
rect 7432 17620 7438 17632
rect 8018 17620 8024 17632
rect 8076 17620 8082 17672
rect 12066 17660 12072 17672
rect 12027 17632 12072 17660
rect 12066 17620 12072 17632
rect 12124 17620 12130 17672
rect 12529 17663 12587 17669
rect 12529 17629 12541 17663
rect 12575 17660 12587 17663
rect 12575 17632 13492 17660
rect 12575 17629 12587 17632
rect 12529 17623 12587 17629
rect 7650 17592 7656 17604
rect 7116 17564 7656 17592
rect 7650 17552 7656 17564
rect 7708 17552 7714 17604
rect 13464 17592 13492 17632
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14737 17663 14795 17669
rect 14737 17660 14749 17663
rect 13872 17632 14749 17660
rect 13872 17620 13878 17632
rect 14737 17629 14749 17632
rect 14783 17629 14795 17663
rect 14737 17623 14795 17629
rect 18874 17620 18880 17672
rect 18932 17660 18938 17672
rect 20180 17660 20208 17691
rect 20254 17688 20260 17740
rect 20312 17728 20318 17740
rect 20438 17737 20444 17740
rect 20395 17731 20444 17737
rect 20312 17700 20357 17728
rect 20312 17688 20318 17700
rect 20395 17697 20407 17731
rect 20441 17697 20444 17731
rect 20395 17691 20444 17697
rect 20438 17688 20444 17691
rect 20496 17688 20502 17740
rect 18932 17632 20208 17660
rect 18932 17620 18938 17632
rect 14090 17592 14096 17604
rect 13464 17564 14096 17592
rect 14090 17552 14096 17564
rect 14148 17552 14154 17604
rect 1581 17527 1639 17533
rect 1581 17493 1593 17527
rect 1627 17524 1639 17527
rect 2314 17524 2320 17536
rect 1627 17496 2320 17524
rect 1627 17493 1639 17496
rect 1581 17487 1639 17493
rect 2314 17484 2320 17496
rect 2372 17484 2378 17536
rect 5997 17527 6055 17533
rect 5997 17493 6009 17527
rect 6043 17524 6055 17527
rect 6086 17524 6092 17536
rect 6043 17496 6092 17524
rect 6043 17493 6055 17496
rect 5997 17487 6055 17493
rect 6086 17484 6092 17496
rect 6144 17484 6150 17536
rect 7009 17527 7067 17533
rect 7009 17493 7021 17527
rect 7055 17524 7067 17527
rect 8294 17524 8300 17536
rect 7055 17496 8300 17524
rect 7055 17493 7067 17496
rect 7009 17487 7067 17493
rect 8294 17484 8300 17496
rect 8352 17484 8358 17536
rect 8662 17484 8668 17536
rect 8720 17524 8726 17536
rect 9582 17524 9588 17536
rect 8720 17496 9588 17524
rect 8720 17484 8726 17496
rect 9582 17484 9588 17496
rect 9640 17524 9646 17536
rect 11241 17527 11299 17533
rect 11241 17524 11253 17527
rect 9640 17496 11253 17524
rect 9640 17484 9646 17496
rect 11241 17493 11253 17496
rect 11287 17493 11299 17527
rect 11241 17487 11299 17493
rect 13998 17484 14004 17536
rect 14056 17524 14062 17536
rect 14829 17527 14887 17533
rect 14829 17524 14841 17527
rect 14056 17496 14841 17524
rect 14056 17484 14062 17496
rect 14829 17493 14841 17496
rect 14875 17493 14887 17527
rect 14829 17487 14887 17493
rect 17310 17484 17316 17536
rect 17368 17524 17374 17536
rect 17405 17527 17463 17533
rect 17405 17524 17417 17527
rect 17368 17496 17417 17524
rect 17368 17484 17374 17496
rect 17405 17493 17417 17496
rect 17451 17493 17463 17527
rect 18966 17524 18972 17536
rect 18927 17496 18972 17524
rect 17405 17487 17463 17493
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 19610 17484 19616 17536
rect 19668 17524 19674 17536
rect 20533 17527 20591 17533
rect 20533 17524 20545 17527
rect 19668 17496 20545 17524
rect 19668 17484 19674 17496
rect 20533 17493 20545 17496
rect 20579 17493 20591 17527
rect 20533 17487 20591 17493
rect 1104 17434 21804 17456
rect 1104 17382 4432 17434
rect 4484 17382 4496 17434
rect 4548 17382 4560 17434
rect 4612 17382 4624 17434
rect 4676 17382 11332 17434
rect 11384 17382 11396 17434
rect 11448 17382 11460 17434
rect 11512 17382 11524 17434
rect 11576 17382 18232 17434
rect 18284 17382 18296 17434
rect 18348 17382 18360 17434
rect 18412 17382 18424 17434
rect 18476 17382 21804 17434
rect 1104 17360 21804 17382
rect 8018 17320 8024 17332
rect 7979 17292 8024 17320
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 8113 17323 8171 17329
rect 8113 17289 8125 17323
rect 8159 17320 8171 17323
rect 8294 17320 8300 17332
rect 8159 17292 8300 17320
rect 8159 17289 8171 17292
rect 8113 17283 8171 17289
rect 7006 17212 7012 17264
rect 7064 17252 7070 17264
rect 7064 17224 7236 17252
rect 7064 17212 7070 17224
rect 7098 17184 7104 17196
rect 7059 17156 7104 17184
rect 7098 17144 7104 17156
rect 7156 17144 7162 17196
rect 7208 17193 7236 17224
rect 7282 17212 7288 17264
rect 7340 17212 7346 17264
rect 7193 17187 7251 17193
rect 7193 17153 7205 17187
rect 7239 17153 7251 17187
rect 7300 17184 7328 17212
rect 7929 17187 7987 17193
rect 7929 17184 7941 17187
rect 7300 17156 7941 17184
rect 7193 17147 7251 17153
rect 7929 17153 7941 17156
rect 7975 17153 7987 17187
rect 7929 17147 7987 17153
rect 5905 17119 5963 17125
rect 5905 17085 5917 17119
rect 5951 17116 5963 17119
rect 5994 17116 6000 17128
rect 5951 17088 6000 17116
rect 5951 17085 5963 17088
rect 5905 17079 5963 17085
rect 5994 17076 6000 17088
rect 6052 17076 6058 17128
rect 7009 17119 7067 17125
rect 7009 17085 7021 17119
rect 7055 17085 7067 17119
rect 7009 17079 7067 17085
rect 7285 17119 7343 17125
rect 7285 17085 7297 17119
rect 7331 17116 7343 17119
rect 7374 17116 7380 17128
rect 7331 17088 7380 17116
rect 7331 17085 7343 17088
rect 7285 17079 7343 17085
rect 5813 17051 5871 17057
rect 5813 17017 5825 17051
rect 5859 17048 5871 17051
rect 6730 17048 6736 17060
rect 5859 17020 6736 17048
rect 5859 17017 5871 17020
rect 5813 17011 5871 17017
rect 6730 17008 6736 17020
rect 6788 17048 6794 17060
rect 7024 17048 7052 17079
rect 7374 17076 7380 17088
rect 7432 17076 7438 17128
rect 7469 17119 7527 17125
rect 7469 17085 7481 17119
rect 7515 17116 7527 17119
rect 7558 17116 7564 17128
rect 7515 17088 7564 17116
rect 7515 17085 7527 17088
rect 7469 17079 7527 17085
rect 7558 17076 7564 17088
rect 7616 17116 7622 17128
rect 8128 17116 8156 17283
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 11882 17280 11888 17332
rect 11940 17320 11946 17332
rect 12069 17323 12127 17329
rect 12069 17320 12081 17323
rect 11940 17292 12081 17320
rect 11940 17280 11946 17292
rect 12069 17289 12081 17292
rect 12115 17289 12127 17323
rect 12069 17283 12127 17289
rect 18877 17323 18935 17329
rect 18877 17289 18889 17323
rect 18923 17320 18935 17323
rect 19058 17320 19064 17332
rect 18923 17292 19064 17320
rect 18923 17289 18935 17292
rect 18877 17283 18935 17289
rect 19058 17280 19064 17292
rect 19116 17280 19122 17332
rect 20254 17280 20260 17332
rect 20312 17320 20318 17332
rect 21085 17323 21143 17329
rect 21085 17320 21097 17323
rect 20312 17292 21097 17320
rect 20312 17280 20318 17292
rect 21085 17289 21097 17292
rect 21131 17289 21143 17323
rect 21085 17283 21143 17289
rect 18598 17184 18604 17196
rect 17972 17156 18604 17184
rect 7616 17088 8156 17116
rect 8205 17119 8263 17125
rect 7616 17076 7622 17088
rect 8205 17085 8217 17119
rect 8251 17085 8263 17119
rect 8662 17116 8668 17128
rect 8623 17088 8668 17116
rect 8205 17079 8263 17085
rect 6788 17020 7052 17048
rect 6788 17008 6794 17020
rect 7650 17008 7656 17060
rect 7708 17048 7714 17060
rect 8220 17048 8248 17079
rect 8662 17076 8668 17088
rect 8720 17076 8726 17128
rect 15473 17119 15531 17125
rect 15473 17085 15485 17119
rect 15519 17116 15531 17119
rect 15562 17116 15568 17128
rect 15519 17088 15568 17116
rect 15519 17085 15531 17088
rect 15473 17079 15531 17085
rect 15562 17076 15568 17088
rect 15620 17076 15626 17128
rect 17402 17076 17408 17128
rect 17460 17116 17466 17128
rect 17497 17119 17555 17125
rect 17497 17116 17509 17119
rect 17460 17088 17509 17116
rect 17460 17076 17466 17088
rect 17497 17085 17509 17088
rect 17543 17085 17555 17119
rect 17497 17079 17555 17085
rect 17586 17076 17592 17128
rect 17644 17116 17650 17128
rect 17972 17125 18000 17156
rect 18598 17144 18604 17156
rect 18656 17184 18662 17196
rect 19242 17184 19248 17196
rect 18656 17156 19248 17184
rect 18656 17144 18662 17156
rect 19242 17144 19248 17156
rect 19300 17144 19306 17196
rect 19610 17184 19616 17196
rect 19571 17156 19616 17184
rect 19610 17144 19616 17156
rect 19668 17144 19674 17196
rect 17865 17119 17923 17125
rect 17644 17088 17689 17116
rect 17644 17076 17650 17088
rect 17865 17085 17877 17119
rect 17911 17085 17923 17119
rect 17865 17079 17923 17085
rect 17957 17119 18015 17125
rect 17957 17085 17969 17119
rect 18003 17085 18015 17119
rect 17957 17079 18015 17085
rect 18417 17119 18475 17125
rect 18417 17085 18429 17119
rect 18463 17085 18475 17119
rect 18690 17116 18696 17128
rect 18651 17088 18696 17116
rect 18417 17079 18475 17085
rect 7708 17020 8248 17048
rect 7708 17008 7714 17020
rect 11790 17008 11796 17060
rect 11848 17048 11854 17060
rect 12253 17051 12311 17057
rect 12253 17048 12265 17051
rect 11848 17020 12265 17048
rect 11848 17008 11854 17020
rect 12253 17017 12265 17020
rect 12299 17017 12311 17051
rect 12253 17011 12311 17017
rect 12434 17008 12440 17060
rect 12492 17048 12498 17060
rect 15197 17051 15255 17057
rect 12492 17020 12537 17048
rect 12492 17008 12498 17020
rect 6822 16980 6828 16992
rect 6783 16952 6828 16980
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 8386 16940 8392 16992
rect 8444 16980 8450 16992
rect 8757 16983 8815 16989
rect 8757 16980 8769 16983
rect 8444 16952 8769 16980
rect 8444 16940 8450 16952
rect 8757 16949 8769 16952
rect 8803 16949 8815 16983
rect 8757 16943 8815 16949
rect 13725 16983 13783 16989
rect 13725 16949 13737 16983
rect 13771 16980 13783 16983
rect 13906 16980 13912 16992
rect 13771 16952 13912 16980
rect 13771 16949 13783 16952
rect 13725 16943 13783 16949
rect 13906 16940 13912 16952
rect 13964 16940 13970 16992
rect 14752 16980 14780 17034
rect 15197 17017 15209 17051
rect 15243 17048 15255 17051
rect 15286 17048 15292 17060
rect 15243 17020 15292 17048
rect 15243 17017 15255 17020
rect 15197 17011 15255 17017
rect 15286 17008 15292 17020
rect 15344 17008 15350 17060
rect 17678 17048 17684 17060
rect 17639 17020 17684 17048
rect 17678 17008 17684 17020
rect 17736 17008 17742 17060
rect 15746 16980 15752 16992
rect 14752 16952 15752 16980
rect 15746 16940 15752 16952
rect 15804 16980 15810 16992
rect 16390 16980 16396 16992
rect 15804 16952 16396 16980
rect 15804 16940 15810 16952
rect 16390 16940 16396 16952
rect 16448 16940 16454 16992
rect 16574 16940 16580 16992
rect 16632 16980 16638 16992
rect 17313 16983 17371 16989
rect 17313 16980 17325 16983
rect 16632 16952 17325 16980
rect 16632 16940 16638 16952
rect 17313 16949 17325 16952
rect 17359 16949 17371 16983
rect 17313 16943 17371 16949
rect 17494 16940 17500 16992
rect 17552 16980 17558 16992
rect 17880 16980 17908 17079
rect 18432 17048 18460 17079
rect 18690 17076 18696 17088
rect 18748 17076 18754 17128
rect 19334 17116 19340 17128
rect 19295 17088 19340 17116
rect 19334 17076 19340 17088
rect 19392 17076 19398 17128
rect 18966 17048 18972 17060
rect 18432 17020 18972 17048
rect 18966 17008 18972 17020
rect 19024 17008 19030 17060
rect 20622 17008 20628 17060
rect 20680 17008 20686 17060
rect 18509 16983 18567 16989
rect 18509 16980 18521 16983
rect 17552 16952 18521 16980
rect 17552 16940 17558 16952
rect 18509 16949 18521 16952
rect 18555 16980 18567 16983
rect 19058 16980 19064 16992
rect 18555 16952 19064 16980
rect 18555 16949 18567 16952
rect 18509 16943 18567 16949
rect 19058 16940 19064 16952
rect 19116 16940 19122 16992
rect 1104 16890 21804 16912
rect 1104 16838 7882 16890
rect 7934 16838 7946 16890
rect 7998 16838 8010 16890
rect 8062 16838 8074 16890
rect 8126 16838 14782 16890
rect 14834 16838 14846 16890
rect 14898 16838 14910 16890
rect 14962 16838 14974 16890
rect 15026 16838 21804 16890
rect 1104 16816 21804 16838
rect 1857 16779 1915 16785
rect 1857 16745 1869 16779
rect 1903 16776 1915 16779
rect 2406 16776 2412 16788
rect 1903 16748 2412 16776
rect 1903 16745 1915 16748
rect 1857 16739 1915 16745
rect 2406 16736 2412 16748
rect 2464 16736 2470 16788
rect 2501 16779 2559 16785
rect 2501 16745 2513 16779
rect 2547 16776 2559 16779
rect 4246 16776 4252 16788
rect 2547 16748 4252 16776
rect 2547 16745 2559 16748
rect 2501 16739 2559 16745
rect 4246 16736 4252 16748
rect 4304 16736 4310 16788
rect 11425 16779 11483 16785
rect 11425 16745 11437 16779
rect 11471 16776 11483 16779
rect 11882 16776 11888 16788
rect 11471 16748 11888 16776
rect 11471 16745 11483 16748
rect 11425 16739 11483 16745
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 12069 16779 12127 16785
rect 12069 16745 12081 16779
rect 12115 16776 12127 16779
rect 12158 16776 12164 16788
rect 12115 16748 12164 16776
rect 12115 16745 12127 16748
rect 12069 16739 12127 16745
rect 12158 16736 12164 16748
rect 12216 16736 12222 16788
rect 13630 16736 13636 16788
rect 13688 16776 13694 16788
rect 15286 16776 15292 16788
rect 13688 16748 14964 16776
rect 15247 16748 15292 16776
rect 13688 16736 13694 16748
rect 12434 16708 12440 16720
rect 12406 16668 12440 16708
rect 12492 16708 12498 16720
rect 12802 16708 12808 16720
rect 12492 16680 12808 16708
rect 12492 16668 12498 16680
rect 12802 16668 12808 16680
rect 12860 16668 12866 16720
rect 14936 16717 14964 16748
rect 15286 16736 15292 16748
rect 15344 16736 15350 16788
rect 18049 16779 18107 16785
rect 18049 16745 18061 16779
rect 18095 16745 18107 16779
rect 18049 16739 18107 16745
rect 14921 16711 14979 16717
rect 14921 16677 14933 16711
rect 14967 16677 14979 16711
rect 16574 16708 16580 16720
rect 16535 16680 16580 16708
rect 14921 16671 14979 16677
rect 16574 16668 16580 16680
rect 16632 16668 16638 16720
rect 17310 16668 17316 16720
rect 17368 16668 17374 16720
rect 18064 16708 18092 16739
rect 18690 16736 18696 16788
rect 18748 16776 18754 16788
rect 20073 16779 20131 16785
rect 20073 16776 20085 16779
rect 18748 16748 20085 16776
rect 18748 16736 18754 16748
rect 20073 16745 20085 16748
rect 20119 16745 20131 16779
rect 20073 16739 20131 16745
rect 20622 16736 20628 16788
rect 20680 16776 20686 16788
rect 20809 16779 20867 16785
rect 20809 16776 20821 16779
rect 20680 16748 20821 16776
rect 20680 16736 20686 16748
rect 20809 16745 20821 16748
rect 20855 16745 20867 16779
rect 20809 16739 20867 16745
rect 18064 16680 18920 16708
rect 1670 16640 1676 16652
rect 1631 16612 1676 16640
rect 1670 16600 1676 16612
rect 1728 16600 1734 16652
rect 2314 16640 2320 16652
rect 2275 16612 2320 16640
rect 2314 16600 2320 16612
rect 2372 16600 2378 16652
rect 6086 16600 6092 16652
rect 6144 16640 6150 16652
rect 7285 16643 7343 16649
rect 7285 16640 7297 16643
rect 6144 16612 7297 16640
rect 6144 16600 6150 16612
rect 7285 16609 7297 16612
rect 7331 16609 7343 16643
rect 7285 16603 7343 16609
rect 7377 16643 7435 16649
rect 7377 16609 7389 16643
rect 7423 16640 7435 16643
rect 7650 16640 7656 16652
rect 7423 16612 7656 16640
rect 7423 16609 7435 16612
rect 7377 16603 7435 16609
rect 7650 16600 7656 16612
rect 7708 16600 7714 16652
rect 11790 16640 11796 16652
rect 11751 16612 11796 16640
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16640 11943 16643
rect 12406 16640 12434 16668
rect 18892 16652 18920 16680
rect 18966 16668 18972 16720
rect 19024 16708 19030 16720
rect 19024 16680 20208 16708
rect 19024 16668 19030 16680
rect 13630 16640 13636 16652
rect 11931 16612 12434 16640
rect 13591 16612 13636 16640
rect 11931 16609 11943 16612
rect 11885 16603 11943 16609
rect 13630 16600 13636 16612
rect 13688 16600 13694 16652
rect 13817 16643 13875 16649
rect 13817 16609 13829 16643
rect 13863 16640 13875 16643
rect 13906 16640 13912 16652
rect 13863 16612 13912 16640
rect 13863 16609 13875 16612
rect 13817 16603 13875 16609
rect 13906 16600 13912 16612
rect 13964 16640 13970 16652
rect 14366 16640 14372 16652
rect 13964 16612 14372 16640
rect 13964 16600 13970 16612
rect 14366 16600 14372 16612
rect 14424 16600 14430 16652
rect 14642 16600 14648 16652
rect 14700 16640 14706 16652
rect 15194 16649 15200 16652
rect 14737 16643 14795 16649
rect 14737 16640 14749 16643
rect 14700 16612 14749 16640
rect 14700 16600 14706 16612
rect 14737 16609 14749 16612
rect 14783 16609 14795 16643
rect 14737 16603 14795 16609
rect 15009 16643 15067 16649
rect 15009 16609 15021 16643
rect 15055 16609 15067 16643
rect 15009 16603 15067 16609
rect 15151 16643 15200 16649
rect 15151 16609 15163 16643
rect 15197 16609 15200 16643
rect 15151 16603 15200 16609
rect 14384 16572 14412 16600
rect 15028 16572 15056 16603
rect 15194 16600 15200 16603
rect 15252 16640 15258 16652
rect 15470 16640 15476 16652
rect 15252 16612 15476 16640
rect 15252 16600 15258 16612
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 15562 16600 15568 16652
rect 15620 16640 15626 16652
rect 16301 16643 16359 16649
rect 16301 16640 16313 16643
rect 15620 16612 16313 16640
rect 15620 16600 15626 16612
rect 16301 16609 16313 16612
rect 16347 16609 16359 16643
rect 18874 16640 18880 16652
rect 18835 16612 18880 16640
rect 16301 16603 16359 16609
rect 18874 16600 18880 16612
rect 18932 16600 18938 16652
rect 19058 16640 19064 16652
rect 18984 16612 19064 16640
rect 18984 16581 19012 16612
rect 19058 16600 19064 16612
rect 19116 16640 19122 16652
rect 20180 16649 20208 16680
rect 19981 16643 20039 16649
rect 19981 16640 19993 16643
rect 19116 16612 19993 16640
rect 19116 16600 19122 16612
rect 19981 16609 19993 16612
rect 20027 16609 20039 16643
rect 19981 16603 20039 16609
rect 20165 16643 20223 16649
rect 20165 16609 20177 16643
rect 20211 16609 20223 16643
rect 20165 16603 20223 16609
rect 20898 16600 20904 16652
rect 20956 16640 20962 16652
rect 20993 16643 21051 16649
rect 20993 16640 21005 16643
rect 20956 16612 21005 16640
rect 20956 16600 20962 16612
rect 20993 16609 21005 16612
rect 21039 16609 21051 16643
rect 20993 16603 21051 16609
rect 14384 16544 15056 16572
rect 18969 16575 19027 16581
rect 18969 16541 18981 16575
rect 19015 16541 19027 16575
rect 18969 16535 19027 16541
rect 13814 16504 13820 16516
rect 13775 16476 13820 16504
rect 13814 16464 13820 16476
rect 13872 16464 13878 16516
rect 1104 16346 21804 16368
rect 1104 16294 4432 16346
rect 4484 16294 4496 16346
rect 4548 16294 4560 16346
rect 4612 16294 4624 16346
rect 4676 16294 11332 16346
rect 11384 16294 11396 16346
rect 11448 16294 11460 16346
rect 11512 16294 11524 16346
rect 11576 16294 18232 16346
rect 18284 16294 18296 16346
rect 18348 16294 18360 16346
rect 18412 16294 18424 16346
rect 18476 16294 21804 16346
rect 1104 16272 21804 16294
rect 2685 16235 2743 16241
rect 2685 16201 2697 16235
rect 2731 16232 2743 16235
rect 11790 16232 11796 16244
rect 2731 16204 11796 16232
rect 2731 16201 2743 16204
rect 2685 16195 2743 16201
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 12802 16232 12808 16244
rect 12763 16204 12808 16232
rect 12802 16192 12808 16204
rect 12860 16192 12866 16244
rect 19150 16232 19156 16244
rect 19111 16204 19156 16232
rect 19150 16192 19156 16204
rect 19208 16192 19214 16244
rect 20714 16232 20720 16244
rect 20675 16204 20720 16232
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 7009 16167 7067 16173
rect 7009 16133 7021 16167
rect 7055 16164 7067 16167
rect 7558 16164 7564 16176
rect 7055 16136 7564 16164
rect 7055 16133 7067 16136
rect 7009 16127 7067 16133
rect 7558 16124 7564 16136
rect 7616 16124 7622 16176
rect 17313 16167 17371 16173
rect 17313 16133 17325 16167
rect 17359 16164 17371 16167
rect 17678 16164 17684 16176
rect 17359 16136 17684 16164
rect 17359 16133 17371 16136
rect 17313 16127 17371 16133
rect 17678 16124 17684 16136
rect 17736 16124 17742 16176
rect 3329 16099 3387 16105
rect 3329 16065 3341 16099
rect 3375 16096 3387 16099
rect 4154 16096 4160 16108
rect 3375 16068 4160 16096
rect 3375 16065 3387 16068
rect 3329 16059 3387 16065
rect 4154 16056 4160 16068
rect 4212 16056 4218 16108
rect 5718 16056 5724 16108
rect 5776 16096 5782 16108
rect 6825 16099 6883 16105
rect 6825 16096 6837 16099
rect 5776 16068 6837 16096
rect 5776 16056 5782 16068
rect 6825 16065 6837 16068
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 7466 16056 7472 16108
rect 7524 16096 7530 16108
rect 8757 16099 8815 16105
rect 8757 16096 8769 16099
rect 7524 16068 8769 16096
rect 7524 16056 7530 16068
rect 8757 16065 8769 16068
rect 8803 16065 8815 16099
rect 8757 16059 8815 16065
rect 8846 16056 8852 16108
rect 8904 16096 8910 16108
rect 8941 16099 8999 16105
rect 8941 16096 8953 16099
rect 8904 16068 8953 16096
rect 8904 16056 8910 16068
rect 8941 16065 8953 16068
rect 8987 16096 8999 16099
rect 9674 16096 9680 16108
rect 8987 16068 9680 16096
rect 8987 16065 8999 16068
rect 8941 16059 8999 16065
rect 9674 16056 9680 16068
rect 9732 16056 9738 16108
rect 13357 16099 13415 16105
rect 13357 16096 13369 16099
rect 12912 16068 13369 16096
rect 2130 15988 2136 16040
rect 2188 16028 2194 16040
rect 2593 16031 2651 16037
rect 2593 16028 2605 16031
rect 2188 16000 2605 16028
rect 2188 15988 2194 16000
rect 2593 15997 2605 16000
rect 2639 15997 2651 16031
rect 2593 15991 2651 15997
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 9030 16028 9036 16040
rect 7156 16000 7201 16028
rect 8991 16000 9036 16028
rect 7156 15988 7162 16000
rect 9030 15988 9036 16000
rect 9088 15988 9094 16040
rect 10502 16028 10508 16040
rect 10463 16000 10508 16028
rect 10502 15988 10508 16000
rect 10560 16028 10566 16040
rect 10962 16028 10968 16040
rect 10560 16000 10968 16028
rect 10560 15988 10566 16000
rect 10962 15988 10968 16000
rect 11020 15988 11026 16040
rect 3605 15963 3663 15969
rect 3605 15929 3617 15963
rect 3651 15929 3663 15963
rect 3605 15923 3663 15929
rect 3620 15892 3648 15923
rect 4338 15920 4344 15972
rect 4396 15920 4402 15972
rect 4982 15892 4988 15904
rect 3620 15864 4988 15892
rect 4982 15852 4988 15864
rect 5040 15852 5046 15904
rect 5077 15895 5135 15901
rect 5077 15861 5089 15895
rect 5123 15892 5135 15895
rect 5626 15892 5632 15904
rect 5123 15864 5632 15892
rect 5123 15861 5135 15864
rect 5077 15855 5135 15861
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 6362 15852 6368 15904
rect 6420 15892 6426 15904
rect 6825 15895 6883 15901
rect 6825 15892 6837 15895
rect 6420 15864 6837 15892
rect 6420 15852 6426 15864
rect 6825 15861 6837 15864
rect 6871 15892 6883 15895
rect 7282 15892 7288 15904
rect 6871 15864 7288 15892
rect 6871 15861 6883 15864
rect 6825 15855 6883 15861
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 8757 15895 8815 15901
rect 8757 15861 8769 15895
rect 8803 15892 8815 15895
rect 9766 15892 9772 15904
rect 8803 15864 9772 15892
rect 8803 15861 8815 15864
rect 8757 15855 8815 15861
rect 9766 15852 9772 15864
rect 9824 15852 9830 15904
rect 10689 15895 10747 15901
rect 10689 15861 10701 15895
rect 10735 15892 10747 15895
rect 10778 15892 10784 15904
rect 10735 15864 10784 15892
rect 10735 15861 10747 15864
rect 10689 15855 10747 15861
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 12912 15892 12940 16068
rect 13357 16065 13369 16068
rect 13403 16096 13415 16099
rect 13909 16099 13967 16105
rect 13909 16096 13921 16099
rect 13403 16068 13921 16096
rect 13403 16065 13415 16068
rect 13357 16059 13415 16065
rect 13909 16065 13921 16068
rect 13955 16065 13967 16099
rect 13909 16059 13967 16065
rect 16942 16056 16948 16108
rect 17000 16096 17006 16108
rect 17865 16099 17923 16105
rect 17865 16096 17877 16099
rect 17000 16068 17877 16096
rect 17000 16056 17006 16068
rect 17865 16065 17877 16068
rect 17911 16065 17923 16099
rect 17865 16059 17923 16065
rect 18984 16068 19564 16096
rect 12986 16031 13044 16037
rect 12986 15997 12998 16031
rect 13032 16028 13044 16031
rect 13449 16031 13507 16037
rect 13449 16028 13461 16031
rect 13032 16000 13461 16028
rect 13032 15997 13044 16000
rect 12986 15991 13044 15997
rect 13449 15997 13461 16000
rect 13495 15997 13507 16031
rect 13449 15991 13507 15997
rect 13464 15960 13492 15991
rect 13814 15988 13820 16040
rect 13872 16028 13878 16040
rect 14093 16031 14151 16037
rect 14093 16028 14105 16031
rect 13872 16000 14105 16028
rect 13872 15988 13878 16000
rect 14093 15997 14105 16000
rect 14139 15997 14151 16031
rect 14366 16028 14372 16040
rect 14327 16000 14372 16028
rect 14093 15991 14151 15997
rect 14366 15988 14372 16000
rect 14424 15988 14430 16040
rect 17497 16031 17555 16037
rect 17497 15997 17509 16031
rect 17543 16028 17555 16031
rect 17586 16028 17592 16040
rect 17543 16000 17592 16028
rect 17543 15997 17555 16000
rect 17497 15991 17555 15997
rect 17586 15988 17592 16000
rect 17644 15988 17650 16040
rect 18690 15988 18696 16040
rect 18748 16028 18754 16040
rect 18984 16037 19012 16068
rect 19536 16037 19564 16068
rect 18969 16031 19027 16037
rect 18969 16028 18981 16031
rect 18748 16000 18981 16028
rect 18748 15988 18754 16000
rect 18969 15997 18981 16000
rect 19015 15997 19027 16031
rect 18969 15991 19027 15997
rect 19153 16031 19211 16037
rect 19153 15997 19165 16031
rect 19199 16028 19211 16031
rect 19521 16031 19579 16037
rect 19199 16000 19472 16028
rect 19199 15997 19211 16000
rect 19153 15991 19211 15997
rect 13998 15960 14004 15972
rect 13464 15932 14004 15960
rect 13998 15920 14004 15932
rect 14056 15920 14062 15972
rect 15470 15920 15476 15972
rect 15528 15960 15534 15972
rect 17681 15963 17739 15969
rect 17681 15960 17693 15963
rect 15528 15932 17693 15960
rect 15528 15920 15534 15932
rect 17681 15929 17693 15932
rect 17727 15960 17739 15963
rect 18598 15960 18604 15972
rect 17727 15932 18604 15960
rect 17727 15929 17739 15932
rect 17681 15923 17739 15929
rect 18598 15920 18604 15932
rect 18656 15920 18662 15972
rect 12989 15895 13047 15901
rect 12989 15892 13001 15895
rect 12912 15864 13001 15892
rect 12989 15861 13001 15864
rect 13035 15861 13047 15895
rect 12989 15855 13047 15861
rect 13630 15852 13636 15904
rect 13688 15892 13694 15904
rect 14277 15895 14335 15901
rect 14277 15892 14289 15895
rect 13688 15864 14289 15892
rect 13688 15852 13694 15864
rect 14277 15861 14289 15864
rect 14323 15861 14335 15895
rect 14277 15855 14335 15861
rect 17402 15852 17408 15904
rect 17460 15892 17466 15904
rect 19444 15901 19472 16000
rect 19521 15997 19533 16031
rect 19567 15997 19579 16031
rect 20898 16028 20904 16040
rect 20859 16000 20904 16028
rect 19521 15991 19579 15997
rect 20898 15988 20904 16000
rect 20956 15988 20962 16040
rect 17589 15895 17647 15901
rect 17589 15892 17601 15895
rect 17460 15864 17601 15892
rect 17460 15852 17466 15864
rect 17589 15861 17601 15864
rect 17635 15861 17647 15895
rect 17589 15855 17647 15861
rect 19429 15895 19487 15901
rect 19429 15861 19441 15895
rect 19475 15892 19487 15895
rect 19978 15892 19984 15904
rect 19475 15864 19984 15892
rect 19475 15861 19487 15864
rect 19429 15855 19487 15861
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 1104 15802 21804 15824
rect 1104 15750 7882 15802
rect 7934 15750 7946 15802
rect 7998 15750 8010 15802
rect 8062 15750 8074 15802
rect 8126 15750 14782 15802
rect 14834 15750 14846 15802
rect 14898 15750 14910 15802
rect 14962 15750 14974 15802
rect 15026 15750 21804 15802
rect 1104 15728 21804 15750
rect 4338 15648 4344 15700
rect 4396 15688 4402 15700
rect 4433 15691 4491 15697
rect 4433 15688 4445 15691
rect 4396 15660 4445 15688
rect 4396 15648 4402 15660
rect 4433 15657 4445 15660
rect 4479 15657 4491 15691
rect 4433 15651 4491 15657
rect 4982 15648 4988 15700
rect 5040 15688 5046 15700
rect 5077 15691 5135 15697
rect 5077 15688 5089 15691
rect 5040 15660 5089 15688
rect 5040 15648 5046 15660
rect 5077 15657 5089 15660
rect 5123 15657 5135 15691
rect 5077 15651 5135 15657
rect 7190 15648 7196 15700
rect 7248 15648 7254 15700
rect 14090 15648 14096 15700
rect 14148 15688 14154 15700
rect 14737 15691 14795 15697
rect 14737 15688 14749 15691
rect 14148 15660 14749 15688
rect 14148 15648 14154 15660
rect 14737 15657 14749 15660
rect 14783 15657 14795 15691
rect 14737 15651 14795 15657
rect 16945 15691 17003 15697
rect 16945 15657 16957 15691
rect 16991 15688 17003 15691
rect 17586 15688 17592 15700
rect 16991 15660 17592 15688
rect 16991 15657 17003 15660
rect 16945 15651 17003 15657
rect 17586 15648 17592 15660
rect 17644 15648 17650 15700
rect 20898 15688 20904 15700
rect 20859 15660 20904 15688
rect 20898 15648 20904 15660
rect 20956 15648 20962 15700
rect 5353 15623 5411 15629
rect 5353 15589 5365 15623
rect 5399 15620 5411 15623
rect 5718 15620 5724 15632
rect 5399 15592 5724 15620
rect 5399 15589 5411 15592
rect 5353 15583 5411 15589
rect 5718 15580 5724 15592
rect 5776 15580 5782 15632
rect 7208 15620 7236 15648
rect 9766 15620 9772 15632
rect 6196 15592 6500 15620
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15552 4675 15555
rect 4890 15552 4896 15564
rect 4663 15524 4896 15552
rect 4663 15521 4675 15524
rect 4617 15515 4675 15521
rect 4890 15512 4896 15524
rect 4948 15512 4954 15564
rect 5258 15552 5264 15564
rect 5219 15524 5264 15552
rect 5258 15512 5264 15524
rect 5316 15512 5322 15564
rect 5626 15561 5632 15564
rect 5445 15555 5503 15561
rect 5445 15521 5457 15555
rect 5491 15521 5503 15555
rect 5445 15515 5503 15521
rect 5583 15555 5632 15561
rect 5583 15521 5595 15555
rect 5629 15521 5632 15555
rect 5583 15515 5632 15521
rect 5460 15416 5488 15515
rect 5626 15512 5632 15515
rect 5684 15512 5690 15564
rect 5721 15487 5779 15493
rect 5721 15453 5733 15487
rect 5767 15484 5779 15487
rect 6196 15484 6224 15592
rect 6362 15552 6368 15564
rect 6323 15524 6368 15552
rect 6362 15512 6368 15524
rect 6420 15512 6426 15564
rect 6472 15552 6500 15592
rect 6840 15592 7972 15620
rect 9727 15592 9772 15620
rect 6840 15561 6868 15592
rect 6825 15555 6883 15561
rect 6825 15552 6837 15555
rect 6472 15524 6837 15552
rect 6825 15521 6837 15524
rect 6871 15521 6883 15555
rect 6825 15515 6883 15521
rect 6918 15555 6976 15561
rect 6918 15521 6930 15555
rect 6964 15521 6976 15555
rect 6918 15515 6976 15521
rect 5767 15456 6224 15484
rect 6273 15487 6331 15493
rect 5767 15453 5779 15456
rect 5721 15447 5779 15453
rect 6273 15453 6285 15487
rect 6319 15484 6331 15487
rect 6932 15484 6960 15515
rect 7006 15512 7012 15564
rect 7064 15561 7070 15564
rect 7064 15555 7113 15561
rect 7064 15521 7067 15555
rect 7101 15521 7113 15555
rect 7190 15552 7196 15564
rect 7151 15524 7196 15552
rect 7064 15515 7113 15521
rect 7064 15512 7070 15515
rect 7190 15512 7196 15524
rect 7248 15512 7254 15564
rect 7282 15512 7288 15564
rect 7340 15561 7346 15564
rect 7944 15561 7972 15592
rect 9766 15580 9772 15592
rect 9824 15580 9830 15632
rect 10778 15580 10784 15632
rect 10836 15580 10842 15632
rect 7340 15552 7348 15561
rect 7929 15555 7987 15561
rect 7340 15524 7385 15552
rect 7340 15515 7348 15524
rect 7929 15521 7941 15555
rect 7975 15521 7987 15555
rect 7929 15515 7987 15521
rect 8022 15555 8080 15561
rect 8022 15521 8034 15555
rect 8068 15521 8080 15555
rect 8202 15552 8208 15564
rect 8163 15524 8208 15552
rect 8022 15515 8080 15521
rect 7340 15512 7346 15515
rect 6319 15456 6960 15484
rect 8036 15484 8064 15515
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 8294 15512 8300 15564
rect 8352 15552 8358 15564
rect 8435 15555 8493 15561
rect 8352 15524 8397 15552
rect 8352 15512 8358 15524
rect 8435 15521 8447 15555
rect 8481 15552 8493 15555
rect 8938 15552 8944 15564
rect 8481 15524 8944 15552
rect 8481 15521 8493 15524
rect 8435 15515 8493 15521
rect 8938 15512 8944 15524
rect 8996 15512 9002 15564
rect 9490 15552 9496 15564
rect 9451 15524 9496 15552
rect 9490 15512 9496 15524
rect 9548 15512 9554 15564
rect 15013 15555 15071 15561
rect 15013 15521 15025 15555
rect 15059 15521 15071 15555
rect 17034 15552 17040 15564
rect 16995 15524 17040 15552
rect 15013 15515 15071 15521
rect 8570 15484 8576 15496
rect 8036 15456 8576 15484
rect 6319 15453 6331 15456
rect 6273 15447 6331 15453
rect 8570 15444 8576 15456
rect 8628 15444 8634 15496
rect 14921 15487 14979 15493
rect 14921 15453 14933 15487
rect 14967 15453 14979 15487
rect 15028 15484 15056 15515
rect 17034 15512 17040 15524
rect 17092 15512 17098 15564
rect 18325 15555 18383 15561
rect 18325 15521 18337 15555
rect 18371 15552 18383 15555
rect 18782 15552 18788 15564
rect 18371 15524 18788 15552
rect 18371 15521 18383 15524
rect 18325 15515 18383 15521
rect 18782 15512 18788 15524
rect 18840 15512 18846 15564
rect 21082 15552 21088 15564
rect 21043 15524 21088 15552
rect 21082 15512 21088 15524
rect 21140 15512 21146 15564
rect 15286 15484 15292 15496
rect 15028 15456 15292 15484
rect 14921 15447 14979 15453
rect 8846 15416 8852 15428
rect 5460 15388 8852 15416
rect 8846 15376 8852 15388
rect 8904 15376 8910 15428
rect 14936 15416 14964 15447
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 15378 15444 15384 15496
rect 15436 15484 15442 15496
rect 15436 15456 15481 15484
rect 15436 15444 15442 15456
rect 15396 15416 15424 15444
rect 14936 15388 15424 15416
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15348 1639 15351
rect 1854 15348 1860 15360
rect 1627 15320 1860 15348
rect 1627 15317 1639 15320
rect 1581 15311 1639 15317
rect 1854 15308 1860 15320
rect 1912 15308 1918 15360
rect 7466 15348 7472 15360
rect 7427 15320 7472 15348
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 8573 15351 8631 15357
rect 8573 15317 8585 15351
rect 8619 15348 8631 15351
rect 9950 15348 9956 15360
rect 8619 15320 9956 15348
rect 8619 15317 8631 15320
rect 8573 15311 8631 15317
rect 9950 15308 9956 15320
rect 10008 15308 10014 15360
rect 10134 15308 10140 15360
rect 10192 15348 10198 15360
rect 11241 15351 11299 15357
rect 11241 15348 11253 15351
rect 10192 15320 11253 15348
rect 10192 15308 10198 15320
rect 11241 15317 11253 15320
rect 11287 15317 11299 15351
rect 11241 15311 11299 15317
rect 14090 15308 14096 15360
rect 14148 15348 14154 15360
rect 15562 15348 15568 15360
rect 14148 15320 15568 15348
rect 14148 15308 14154 15320
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 17954 15308 17960 15360
rect 18012 15348 18018 15360
rect 18233 15351 18291 15357
rect 18233 15348 18245 15351
rect 18012 15320 18245 15348
rect 18012 15308 18018 15320
rect 18233 15317 18245 15320
rect 18279 15317 18291 15351
rect 18233 15311 18291 15317
rect 1104 15258 21804 15280
rect 1104 15206 4432 15258
rect 4484 15206 4496 15258
rect 4548 15206 4560 15258
rect 4612 15206 4624 15258
rect 4676 15206 11332 15258
rect 11384 15206 11396 15258
rect 11448 15206 11460 15258
rect 11512 15206 11524 15258
rect 11576 15206 18232 15258
rect 18284 15206 18296 15258
rect 18348 15206 18360 15258
rect 18412 15206 18424 15258
rect 18476 15206 21804 15258
rect 1104 15184 21804 15206
rect 4985 15147 5043 15153
rect 4985 15113 4997 15147
rect 5031 15144 5043 15147
rect 5258 15144 5264 15156
rect 5031 15116 5264 15144
rect 5031 15113 5043 15116
rect 4985 15107 5043 15113
rect 5258 15104 5264 15116
rect 5316 15104 5322 15156
rect 5537 15147 5595 15153
rect 5537 15113 5549 15147
rect 5583 15144 5595 15147
rect 5718 15144 5724 15156
rect 5583 15116 5724 15144
rect 5583 15113 5595 15116
rect 5537 15107 5595 15113
rect 5718 15104 5724 15116
rect 5776 15104 5782 15156
rect 6638 15104 6644 15156
rect 6696 15144 6702 15156
rect 8389 15147 8447 15153
rect 8389 15144 8401 15147
rect 6696 15116 8401 15144
rect 6696 15104 6702 15116
rect 8389 15113 8401 15116
rect 8435 15144 8447 15147
rect 8938 15144 8944 15156
rect 8435 15116 8616 15144
rect 8899 15116 8944 15144
rect 8435 15113 8447 15116
rect 8389 15107 8447 15113
rect 7006 15036 7012 15088
rect 7064 15076 7070 15088
rect 7193 15079 7251 15085
rect 7193 15076 7205 15079
rect 7064 15048 7205 15076
rect 7064 15036 7070 15048
rect 7193 15045 7205 15048
rect 7239 15076 7251 15079
rect 7929 15079 7987 15085
rect 7929 15076 7941 15079
rect 7239 15048 7941 15076
rect 7239 15045 7251 15048
rect 7193 15039 7251 15045
rect 7929 15045 7941 15048
rect 7975 15045 7987 15079
rect 8588 15076 8616 15116
rect 8938 15104 8944 15116
rect 8996 15104 9002 15156
rect 9674 15104 9680 15156
rect 9732 15144 9738 15156
rect 10137 15147 10195 15153
rect 10137 15144 10149 15147
rect 9732 15116 10149 15144
rect 9732 15104 9738 15116
rect 10137 15113 10149 15116
rect 10183 15113 10195 15147
rect 10137 15107 10195 15113
rect 13998 15104 14004 15156
rect 14056 15144 14062 15156
rect 14369 15147 14427 15153
rect 14369 15144 14381 15147
rect 14056 15116 14381 15144
rect 14056 15104 14062 15116
rect 14369 15113 14381 15116
rect 14415 15113 14427 15147
rect 14369 15107 14427 15113
rect 15286 15104 15292 15156
rect 15344 15144 15350 15156
rect 15473 15147 15531 15153
rect 15473 15144 15485 15147
rect 15344 15116 15485 15144
rect 15344 15104 15350 15116
rect 15473 15113 15485 15116
rect 15519 15113 15531 15147
rect 15473 15107 15531 15113
rect 17034 15104 17040 15156
rect 17092 15144 17098 15156
rect 17313 15147 17371 15153
rect 17313 15144 17325 15147
rect 17092 15116 17325 15144
rect 17092 15104 17098 15116
rect 17313 15113 17325 15116
rect 17359 15113 17371 15147
rect 17494 15144 17500 15156
rect 17455 15116 17500 15144
rect 17313 15107 17371 15113
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 9401 15079 9459 15085
rect 9401 15076 9413 15079
rect 8588 15048 9413 15076
rect 7929 15039 7987 15045
rect 9401 15045 9413 15048
rect 9447 15045 9459 15079
rect 9401 15039 9459 15045
rect 10962 15036 10968 15088
rect 11020 15076 11026 15088
rect 15194 15076 15200 15088
rect 11020 15048 15200 15076
rect 11020 15036 11026 15048
rect 6730 15008 6736 15020
rect 5736 14980 6736 15008
rect 1854 14940 1860 14952
rect 1815 14912 1860 14940
rect 1854 14900 1860 14912
rect 1912 14900 1918 14952
rect 5736 14949 5764 14980
rect 6730 14968 6736 14980
rect 6788 15008 6794 15020
rect 7101 15011 7159 15017
rect 7101 15008 7113 15011
rect 6788 14980 7113 15008
rect 6788 14968 6794 14980
rect 7101 14977 7113 14980
rect 7147 14977 7159 15011
rect 7466 15008 7472 15020
rect 7427 14980 7472 15008
rect 7101 14971 7159 14977
rect 7466 14968 7472 14980
rect 7524 14968 7530 15020
rect 7558 14968 7564 15020
rect 7616 15008 7622 15020
rect 9950 15008 9956 15020
rect 7616 14980 9260 15008
rect 9911 14980 9956 15008
rect 7616 14968 7622 14980
rect 4893 14943 4951 14949
rect 4893 14909 4905 14943
rect 4939 14909 4951 14943
rect 4893 14903 4951 14909
rect 5077 14943 5135 14949
rect 5077 14909 5089 14943
rect 5123 14940 5135 14943
rect 5721 14943 5779 14949
rect 5721 14940 5733 14943
rect 5123 14912 5733 14940
rect 5123 14909 5135 14912
rect 5077 14903 5135 14909
rect 5721 14909 5733 14912
rect 5767 14909 5779 14943
rect 6822 14940 6828 14952
rect 6783 14912 6828 14940
rect 5721 14903 5779 14909
rect 2038 14804 2044 14816
rect 1999 14776 2044 14804
rect 2038 14764 2044 14776
rect 2096 14764 2102 14816
rect 2314 14764 2320 14816
rect 2372 14804 2378 14816
rect 2685 14807 2743 14813
rect 2685 14804 2697 14807
rect 2372 14776 2697 14804
rect 2372 14764 2378 14776
rect 2685 14773 2697 14776
rect 2731 14773 2743 14807
rect 2685 14767 2743 14773
rect 2777 14807 2835 14813
rect 2777 14773 2789 14807
rect 2823 14804 2835 14807
rect 3510 14804 3516 14816
rect 2823 14776 3516 14804
rect 2823 14773 2835 14776
rect 2777 14767 2835 14773
rect 3510 14764 3516 14776
rect 3568 14764 3574 14816
rect 4908 14804 4936 14903
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 6914 14900 6920 14952
rect 6972 14940 6978 14952
rect 7009 14943 7067 14949
rect 7009 14940 7021 14943
rect 6972 14912 7021 14940
rect 6972 14900 6978 14912
rect 7009 14909 7021 14912
rect 7055 14909 7067 14943
rect 7009 14903 7067 14909
rect 7285 14943 7343 14949
rect 7285 14909 7297 14943
rect 7331 14909 7343 14943
rect 7285 14903 7343 14909
rect 5905 14875 5963 14881
rect 5905 14841 5917 14875
rect 5951 14872 5963 14875
rect 6178 14872 6184 14884
rect 5951 14844 6184 14872
rect 5951 14841 5963 14844
rect 5905 14835 5963 14841
rect 5920 14804 5948 14835
rect 6178 14832 6184 14844
rect 6236 14872 6242 14884
rect 7300 14872 7328 14903
rect 7742 14900 7748 14952
rect 7800 14940 7806 14952
rect 8220 14949 8248 14980
rect 8113 14943 8171 14949
rect 8113 14940 8125 14943
rect 7800 14912 8125 14940
rect 7800 14900 7806 14912
rect 8113 14909 8125 14912
rect 8159 14909 8171 14943
rect 8113 14903 8171 14909
rect 8205 14943 8263 14949
rect 8205 14909 8217 14943
rect 8251 14909 8263 14943
rect 8205 14903 8263 14909
rect 8481 14943 8539 14949
rect 8481 14909 8493 14943
rect 8527 14940 8539 14943
rect 9030 14940 9036 14952
rect 8527 14912 9036 14940
rect 8527 14909 8539 14912
rect 8481 14903 8539 14909
rect 9030 14900 9036 14912
rect 9088 14900 9094 14952
rect 9232 14949 9260 14980
rect 9950 14968 9956 14980
rect 10008 14968 10014 15020
rect 9125 14943 9183 14949
rect 9125 14909 9137 14943
rect 9171 14909 9183 14943
rect 9125 14903 9183 14909
rect 9217 14943 9275 14949
rect 9217 14909 9229 14943
rect 9263 14909 9275 14943
rect 9217 14903 9275 14909
rect 9493 14943 9551 14949
rect 9493 14909 9505 14943
rect 9539 14940 9551 14943
rect 9674 14940 9680 14952
rect 9539 14912 9680 14940
rect 9539 14909 9551 14912
rect 9493 14903 9551 14909
rect 6236 14844 7328 14872
rect 6236 14832 6242 14844
rect 4908 14776 5948 14804
rect 6822 14764 6828 14816
rect 6880 14804 6886 14816
rect 7558 14804 7564 14816
rect 6880 14776 7564 14804
rect 6880 14764 6886 14776
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 9140 14804 9168 14903
rect 9674 14900 9680 14912
rect 9732 14900 9738 14952
rect 12544 14949 12572 15048
rect 15194 15036 15200 15048
rect 15252 15036 15258 15088
rect 15378 15036 15384 15088
rect 15436 15076 15442 15088
rect 18325 15079 18383 15085
rect 18325 15076 18337 15079
rect 15436 15048 18337 15076
rect 15436 15036 15442 15048
rect 14921 15011 14979 15017
rect 14921 14977 14933 15011
rect 14967 15008 14979 15011
rect 16301 15011 16359 15017
rect 16301 15008 16313 15011
rect 14967 14980 16313 15008
rect 14967 14977 14979 14980
rect 14921 14971 14979 14977
rect 16301 14977 16313 14980
rect 16347 14977 16359 15011
rect 16301 14971 16359 14977
rect 10229 14943 10287 14949
rect 10229 14909 10241 14943
rect 10275 14909 10287 14943
rect 10229 14903 10287 14909
rect 12529 14943 12587 14949
rect 12529 14909 12541 14943
rect 12575 14909 12587 14943
rect 12529 14903 12587 14909
rect 14550 14943 14608 14949
rect 14550 14909 14562 14943
rect 14596 14940 14608 14943
rect 14642 14940 14648 14952
rect 14596 14912 14648 14940
rect 14596 14909 14608 14912
rect 14550 14903 14608 14909
rect 10244 14872 10272 14903
rect 14642 14900 14648 14912
rect 14700 14900 14706 14952
rect 15013 14943 15071 14949
rect 15013 14909 15025 14943
rect 15059 14940 15071 14943
rect 15102 14940 15108 14952
rect 15059 14912 15108 14940
rect 15059 14909 15071 14912
rect 15013 14903 15071 14909
rect 15102 14900 15108 14912
rect 15160 14940 15166 14952
rect 16408 14949 16436 15048
rect 18325 15045 18337 15048
rect 18371 15045 18383 15079
rect 18325 15039 18383 15045
rect 17589 15011 17647 15017
rect 17589 14977 17601 15011
rect 17635 15008 17647 15011
rect 17954 15008 17960 15020
rect 17635 14980 17960 15008
rect 17635 14977 17647 14980
rect 17589 14971 17647 14977
rect 17954 14968 17960 14980
rect 18012 14968 18018 15020
rect 19978 15008 19984 15020
rect 18892 14980 19984 15008
rect 15473 14943 15531 14949
rect 15473 14940 15485 14943
rect 15160 14912 15485 14940
rect 15160 14900 15166 14912
rect 15473 14909 15485 14912
rect 15519 14909 15531 14943
rect 15473 14903 15531 14909
rect 15749 14943 15807 14949
rect 15749 14909 15761 14943
rect 15795 14909 15807 14943
rect 15749 14903 15807 14909
rect 16393 14943 16451 14949
rect 16393 14909 16405 14943
rect 16439 14909 16451 14943
rect 16393 14903 16451 14909
rect 10594 14872 10600 14884
rect 9646 14844 10600 14872
rect 9646 14804 9674 14844
rect 10594 14832 10600 14844
rect 10652 14832 10658 14884
rect 15764 14872 15792 14903
rect 17310 14900 17316 14952
rect 17368 14940 17374 14952
rect 17681 14943 17739 14949
rect 17681 14940 17693 14943
rect 17368 14912 17693 14940
rect 17368 14900 17374 14912
rect 17681 14909 17693 14912
rect 17727 14909 17739 14943
rect 17681 14903 17739 14909
rect 18509 14943 18567 14949
rect 18509 14909 18521 14943
rect 18555 14909 18567 14943
rect 18690 14940 18696 14952
rect 18651 14912 18696 14940
rect 18509 14903 18567 14909
rect 14568 14844 15792 14872
rect 14568 14816 14596 14844
rect 9140 14776 9674 14804
rect 9953 14807 10011 14813
rect 9953 14773 9965 14807
rect 9999 14804 10011 14807
rect 11422 14804 11428 14816
rect 9999 14776 11428 14804
rect 9999 14773 10011 14776
rect 9953 14767 10011 14773
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 12342 14804 12348 14816
rect 12303 14776 12348 14804
rect 12342 14764 12348 14776
rect 12400 14764 12406 14816
rect 14550 14804 14556 14816
rect 14511 14776 14556 14804
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 15657 14807 15715 14813
rect 15657 14773 15669 14807
rect 15703 14804 15715 14807
rect 16206 14804 16212 14816
rect 15703 14776 16212 14804
rect 15703 14773 15715 14776
rect 15657 14767 15715 14773
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 18524 14804 18552 14903
rect 18690 14900 18696 14912
rect 18748 14900 18754 14952
rect 18892 14949 18920 14980
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 18877 14943 18935 14949
rect 18877 14909 18889 14943
rect 18923 14909 18935 14943
rect 19334 14940 19340 14952
rect 19295 14912 19340 14940
rect 18877 14903 18935 14909
rect 19334 14900 19340 14912
rect 19392 14900 19398 14952
rect 18601 14875 18659 14881
rect 18601 14841 18613 14875
rect 18647 14872 18659 14875
rect 18782 14872 18788 14884
rect 18647 14844 18788 14872
rect 18647 14841 18659 14844
rect 18601 14835 18659 14841
rect 18782 14832 18788 14844
rect 18840 14832 18846 14884
rect 19610 14872 19616 14884
rect 19571 14844 19616 14872
rect 19610 14832 19616 14844
rect 19668 14832 19674 14884
rect 20622 14832 20628 14884
rect 20680 14832 20686 14884
rect 19702 14804 19708 14816
rect 18524 14776 19708 14804
rect 19702 14764 19708 14776
rect 19760 14804 19766 14816
rect 20254 14804 20260 14816
rect 19760 14776 20260 14804
rect 19760 14764 19766 14776
rect 20254 14764 20260 14776
rect 20312 14804 20318 14816
rect 21085 14807 21143 14813
rect 21085 14804 21097 14807
rect 20312 14776 21097 14804
rect 20312 14764 20318 14776
rect 21085 14773 21097 14776
rect 21131 14773 21143 14807
rect 21085 14767 21143 14773
rect 1104 14714 21804 14736
rect 1104 14662 7882 14714
rect 7934 14662 7946 14714
rect 7998 14662 8010 14714
rect 8062 14662 8074 14714
rect 8126 14662 14782 14714
rect 14834 14662 14846 14714
rect 14898 14662 14910 14714
rect 14962 14662 14974 14714
rect 15026 14662 21804 14714
rect 1104 14640 21804 14662
rect 6178 14600 6184 14612
rect 6139 14572 6184 14600
rect 6178 14560 6184 14572
rect 6236 14560 6242 14612
rect 6822 14600 6828 14612
rect 6472 14572 6828 14600
rect 5626 14492 5632 14544
rect 5684 14532 5690 14544
rect 6472 14541 6500 14572
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 7190 14560 7196 14612
rect 7248 14600 7254 14612
rect 7285 14603 7343 14609
rect 7285 14600 7297 14603
rect 7248 14572 7297 14600
rect 7248 14560 7254 14572
rect 7285 14569 7297 14572
rect 7331 14569 7343 14603
rect 7285 14563 7343 14569
rect 8294 14560 8300 14612
rect 8352 14600 8358 14612
rect 8481 14603 8539 14609
rect 8481 14600 8493 14603
rect 8352 14572 8493 14600
rect 8352 14560 8358 14572
rect 8481 14569 8493 14572
rect 8527 14569 8539 14603
rect 8481 14563 8539 14569
rect 9030 14560 9036 14612
rect 9088 14600 9094 14612
rect 9490 14600 9496 14612
rect 9088 14572 9496 14600
rect 9088 14560 9094 14572
rect 9490 14560 9496 14572
rect 9548 14600 9554 14612
rect 9953 14603 10011 14609
rect 9953 14600 9965 14603
rect 9548 14572 9965 14600
rect 9548 14560 9554 14572
rect 9953 14569 9965 14572
rect 9999 14569 10011 14603
rect 10594 14600 10600 14612
rect 10555 14572 10600 14600
rect 9953 14563 10011 14569
rect 10594 14560 10600 14572
rect 10652 14560 10658 14612
rect 12342 14560 12348 14612
rect 12400 14560 12406 14612
rect 14642 14560 14648 14612
rect 14700 14600 14706 14612
rect 14700 14572 15148 14600
rect 14700 14560 14706 14572
rect 6457 14535 6515 14541
rect 6457 14532 6469 14535
rect 5684 14504 6469 14532
rect 5684 14492 5690 14504
rect 6457 14501 6469 14504
rect 6503 14501 6515 14535
rect 6457 14495 6515 14501
rect 6549 14535 6607 14541
rect 6549 14501 6561 14535
rect 6595 14532 6607 14535
rect 7098 14532 7104 14544
rect 6595 14504 7104 14532
rect 6595 14501 6607 14504
rect 6549 14495 6607 14501
rect 7098 14492 7104 14504
rect 7156 14492 7162 14544
rect 7558 14492 7564 14544
rect 7616 14532 7622 14544
rect 7742 14532 7748 14544
rect 7616 14504 7748 14532
rect 7616 14492 7622 14504
rect 7742 14492 7748 14504
rect 7800 14532 7806 14544
rect 7800 14504 8524 14532
rect 7800 14492 7806 14504
rect 2314 14464 2320 14476
rect 2275 14436 2320 14464
rect 2314 14424 2320 14436
rect 2372 14424 2378 14476
rect 6365 14467 6423 14473
rect 6365 14433 6377 14467
rect 6411 14433 6423 14467
rect 6730 14464 6736 14476
rect 6691 14436 6736 14464
rect 6365 14427 6423 14433
rect 1946 14396 1952 14408
rect 1907 14368 1952 14396
rect 1946 14356 1952 14368
rect 2004 14356 2010 14408
rect 2774 14356 2780 14408
rect 2832 14396 2838 14408
rect 3142 14396 3148 14408
rect 2832 14368 2877 14396
rect 3103 14368 3148 14396
rect 2832 14356 2838 14368
rect 3142 14356 3148 14368
rect 3200 14356 3206 14408
rect 6380 14396 6408 14427
rect 6730 14424 6736 14436
rect 6788 14424 6794 14476
rect 7006 14424 7012 14476
rect 7064 14464 7070 14476
rect 7377 14467 7435 14473
rect 7377 14464 7389 14467
rect 7064 14436 7389 14464
rect 7064 14424 7070 14436
rect 7377 14433 7389 14436
rect 7423 14433 7435 14467
rect 7377 14427 7435 14433
rect 7466 14424 7472 14476
rect 7524 14464 7530 14476
rect 8202 14464 8208 14476
rect 7524 14436 8208 14464
rect 7524 14424 7530 14436
rect 8202 14424 8208 14436
rect 8260 14464 8266 14476
rect 8389 14467 8447 14473
rect 8389 14464 8401 14467
rect 8260 14436 8401 14464
rect 8260 14424 8266 14436
rect 8389 14433 8401 14436
rect 8435 14433 8447 14467
rect 8496 14464 8524 14504
rect 9674 14492 9680 14544
rect 9732 14532 9738 14544
rect 11422 14532 11428 14544
rect 9732 14504 10548 14532
rect 11383 14504 11428 14532
rect 9732 14492 9738 14504
rect 9861 14467 9919 14473
rect 9861 14464 9873 14467
rect 8496 14436 9873 14464
rect 8389 14427 8447 14433
rect 9861 14433 9873 14436
rect 9907 14464 9919 14467
rect 10134 14464 10140 14476
rect 9907 14436 10140 14464
rect 9907 14433 9919 14436
rect 9861 14427 9919 14433
rect 10134 14424 10140 14436
rect 10192 14424 10198 14476
rect 10520 14473 10548 14504
rect 11422 14492 11428 14504
rect 11480 14492 11486 14544
rect 12360 14518 12388 14560
rect 14550 14492 14556 14544
rect 14608 14532 14614 14544
rect 15010 14532 15016 14544
rect 14608 14504 15016 14532
rect 14608 14492 14614 14504
rect 15010 14492 15016 14504
rect 15068 14492 15074 14544
rect 15120 14541 15148 14572
rect 15194 14560 15200 14612
rect 15252 14600 15258 14612
rect 15746 14600 15752 14612
rect 15252 14572 15752 14600
rect 15252 14560 15258 14572
rect 15746 14560 15752 14572
rect 15804 14560 15810 14612
rect 19978 14600 19984 14612
rect 19939 14572 19984 14600
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 20165 14603 20223 14609
rect 20165 14569 20177 14603
rect 20211 14600 20223 14603
rect 20254 14600 20260 14612
rect 20211 14572 20260 14600
rect 20211 14569 20223 14572
rect 20165 14563 20223 14569
rect 20254 14560 20260 14572
rect 20312 14600 20318 14612
rect 20312 14572 20576 14600
rect 20312 14560 20318 14572
rect 15105 14535 15163 14541
rect 15105 14501 15117 14535
rect 15151 14532 15163 14535
rect 15151 14504 16252 14532
rect 15151 14501 15163 14504
rect 15105 14495 15163 14501
rect 16224 14476 16252 14504
rect 17034 14492 17040 14544
rect 17092 14532 17098 14544
rect 18874 14532 18880 14544
rect 17092 14504 17172 14532
rect 17092 14492 17098 14504
rect 10505 14467 10563 14473
rect 10505 14433 10517 14467
rect 10551 14464 10563 14467
rect 10778 14464 10784 14476
rect 10551 14436 10784 14464
rect 10551 14433 10563 14436
rect 10505 14427 10563 14433
rect 10778 14424 10784 14436
rect 10836 14424 10842 14476
rect 14921 14467 14979 14473
rect 14921 14433 14933 14467
rect 14967 14433 14979 14467
rect 15286 14464 15292 14476
rect 15247 14436 15292 14464
rect 14921 14427 14979 14433
rect 6638 14396 6644 14408
rect 6380 14368 6644 14396
rect 6638 14356 6644 14368
rect 6696 14356 6702 14408
rect 11146 14396 11152 14408
rect 11107 14368 11152 14396
rect 11146 14356 11152 14368
rect 11204 14356 11210 14408
rect 14936 14396 14964 14427
rect 15286 14424 15292 14436
rect 15344 14424 15350 14476
rect 16206 14464 16212 14476
rect 16167 14436 16212 14464
rect 16206 14424 16212 14436
rect 16264 14424 16270 14476
rect 16942 14464 16948 14476
rect 16903 14436 16948 14464
rect 16942 14424 16948 14436
rect 17000 14424 17006 14476
rect 17144 14473 17172 14504
rect 18340 14504 18880 14532
rect 17129 14467 17187 14473
rect 17129 14433 17141 14467
rect 17175 14433 17187 14467
rect 17129 14427 17187 14433
rect 17954 14424 17960 14476
rect 18012 14464 18018 14476
rect 18340 14473 18368 14504
rect 18874 14492 18880 14504
rect 18932 14492 18938 14544
rect 18049 14467 18107 14473
rect 18049 14464 18061 14467
rect 18012 14436 18061 14464
rect 18012 14424 18018 14436
rect 18049 14433 18061 14436
rect 18095 14433 18107 14467
rect 18049 14427 18107 14433
rect 18325 14467 18383 14473
rect 18325 14433 18337 14467
rect 18371 14433 18383 14467
rect 18325 14427 18383 14433
rect 18417 14467 18475 14473
rect 18417 14433 18429 14467
rect 18463 14433 18475 14467
rect 18598 14464 18604 14476
rect 18559 14436 18604 14464
rect 18417 14427 18475 14433
rect 15470 14396 15476 14408
rect 14936 14368 15476 14396
rect 15470 14356 15476 14368
rect 15528 14396 15534 14408
rect 17037 14399 17095 14405
rect 17037 14396 17049 14399
rect 15528 14368 17049 14396
rect 15528 14356 15534 14368
rect 17037 14365 17049 14368
rect 17083 14365 17095 14399
rect 17037 14359 17095 14365
rect 17221 14399 17279 14405
rect 17221 14365 17233 14399
rect 17267 14396 17279 14399
rect 17402 14396 17408 14408
rect 17267 14368 17408 14396
rect 17267 14365 17279 14368
rect 17221 14359 17279 14365
rect 17402 14356 17408 14368
rect 17460 14356 17466 14408
rect 17494 14356 17500 14408
rect 17552 14396 17558 14408
rect 18233 14399 18291 14405
rect 18233 14396 18245 14399
rect 17552 14368 18245 14396
rect 17552 14356 17558 14368
rect 18233 14365 18245 14368
rect 18279 14365 18291 14399
rect 18432 14396 18460 14427
rect 18598 14424 18604 14436
rect 18656 14464 18662 14476
rect 19518 14464 19524 14476
rect 18656 14436 19524 14464
rect 18656 14424 18662 14436
rect 19518 14424 19524 14436
rect 19576 14424 19582 14476
rect 20162 14467 20220 14473
rect 20162 14433 20174 14467
rect 20208 14464 20220 14467
rect 20254 14464 20260 14476
rect 20208 14436 20260 14464
rect 20208 14433 20220 14436
rect 20162 14427 20220 14433
rect 20254 14424 20260 14436
rect 20312 14424 20318 14476
rect 20548 14473 20576 14572
rect 20533 14467 20591 14473
rect 20533 14433 20545 14467
rect 20579 14433 20591 14467
rect 20533 14427 20591 14433
rect 18782 14396 18788 14408
rect 18432 14368 18788 14396
rect 18233 14359 18291 14365
rect 18782 14356 18788 14368
rect 18840 14396 18846 14408
rect 20272 14396 20300 14424
rect 20625 14399 20683 14405
rect 20625 14396 20637 14399
rect 18840 14368 20637 14396
rect 18840 14356 18846 14368
rect 20625 14365 20637 14368
rect 20671 14365 20683 14399
rect 20625 14359 20683 14365
rect 16301 14331 16359 14337
rect 16301 14297 16313 14331
rect 16347 14328 16359 14331
rect 17310 14328 17316 14340
rect 16347 14300 17316 14328
rect 16347 14297 16359 14300
rect 16301 14291 16359 14297
rect 17310 14288 17316 14300
rect 17368 14288 17374 14340
rect 17954 14328 17960 14340
rect 17420 14300 17960 14328
rect 2314 14260 2320 14272
rect 2275 14232 2320 14260
rect 2314 14220 2320 14232
rect 2372 14220 2378 14272
rect 2961 14263 3019 14269
rect 2961 14229 2973 14263
rect 3007 14260 3019 14263
rect 3510 14260 3516 14272
rect 3007 14232 3516 14260
rect 3007 14229 3019 14232
rect 2961 14223 3019 14229
rect 3510 14220 3516 14232
rect 3568 14220 3574 14272
rect 12894 14260 12900 14272
rect 12855 14232 12900 14260
rect 12894 14220 12900 14232
rect 12952 14220 12958 14272
rect 14274 14220 14280 14272
rect 14332 14260 14338 14272
rect 17420 14269 17448 14300
rect 17954 14288 17960 14300
rect 18012 14288 18018 14340
rect 14737 14263 14795 14269
rect 14737 14260 14749 14263
rect 14332 14232 14749 14260
rect 14332 14220 14338 14232
rect 14737 14229 14749 14232
rect 14783 14229 14795 14263
rect 14737 14223 14795 14229
rect 17405 14263 17463 14269
rect 17405 14229 17417 14263
rect 17451 14229 17463 14263
rect 17405 14223 17463 14229
rect 17865 14263 17923 14269
rect 17865 14229 17877 14263
rect 17911 14260 17923 14263
rect 18046 14260 18052 14272
rect 17911 14232 18052 14260
rect 17911 14229 17923 14232
rect 17865 14223 17923 14229
rect 18046 14220 18052 14232
rect 18104 14220 18110 14272
rect 1104 14170 21804 14192
rect 1104 14118 4432 14170
rect 4484 14118 4496 14170
rect 4548 14118 4560 14170
rect 4612 14118 4624 14170
rect 4676 14118 11332 14170
rect 11384 14118 11396 14170
rect 11448 14118 11460 14170
rect 11512 14118 11524 14170
rect 11576 14118 18232 14170
rect 18284 14118 18296 14170
rect 18348 14118 18360 14170
rect 18412 14118 18424 14170
rect 18476 14118 21804 14170
rect 1104 14096 21804 14118
rect 1946 14056 1952 14068
rect 1907 14028 1952 14056
rect 1946 14016 1952 14028
rect 2004 14016 2010 14068
rect 4798 14056 4804 14068
rect 2516 14028 4804 14056
rect 2406 13920 2412 13932
rect 2367 13892 2412 13920
rect 2406 13880 2412 13892
rect 2464 13880 2470 13932
rect 2516 13929 2544 14028
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 8570 14056 8576 14068
rect 8531 14028 8576 14056
rect 8570 14016 8576 14028
rect 8628 14016 8634 14068
rect 15010 14016 15016 14068
rect 15068 14056 15074 14068
rect 15749 14059 15807 14065
rect 15749 14056 15761 14059
rect 15068 14028 15761 14056
rect 15068 14016 15074 14028
rect 15749 14025 15761 14028
rect 15795 14025 15807 14059
rect 17402 14056 17408 14068
rect 17363 14028 17408 14056
rect 15749 14019 15807 14025
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 17494 14016 17500 14068
rect 17552 14056 17558 14068
rect 19429 14059 19487 14065
rect 17552 14028 17597 14056
rect 17552 14016 17558 14028
rect 19429 14025 19441 14059
rect 19475 14056 19487 14059
rect 19610 14056 19616 14068
rect 19475 14028 19616 14056
rect 19475 14025 19487 14028
rect 19429 14019 19487 14025
rect 19610 14016 19616 14028
rect 19668 14016 19674 14068
rect 20622 14016 20628 14068
rect 20680 14056 20686 14068
rect 20717 14059 20775 14065
rect 20717 14056 20729 14059
rect 20680 14028 20729 14056
rect 20680 14016 20686 14028
rect 20717 14025 20729 14028
rect 20763 14025 20775 14059
rect 20717 14019 20775 14025
rect 3513 13991 3571 13997
rect 3513 13957 3525 13991
rect 3559 13988 3571 13991
rect 3973 13991 4031 13997
rect 3973 13988 3985 13991
rect 3559 13960 3985 13988
rect 3559 13957 3571 13960
rect 3513 13951 3571 13957
rect 3973 13957 3985 13960
rect 4019 13957 4031 13991
rect 3973 13951 4031 13957
rect 9493 13991 9551 13997
rect 9493 13957 9505 13991
rect 9539 13957 9551 13991
rect 9493 13951 9551 13957
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13889 2559 13923
rect 3142 13920 3148 13932
rect 3055 13892 3148 13920
rect 2501 13883 2559 13889
rect 2222 13812 2228 13864
rect 2280 13852 2286 13864
rect 2516 13852 2544 13883
rect 3142 13880 3148 13892
rect 3200 13920 3206 13932
rect 9508 13920 9536 13951
rect 16942 13948 16948 14000
rect 17000 13988 17006 14000
rect 17000 13960 18276 13988
rect 17000 13948 17006 13960
rect 3200 13892 9536 13920
rect 10137 13923 10195 13929
rect 3200 13880 3206 13892
rect 10137 13889 10149 13923
rect 10183 13920 10195 13923
rect 12250 13920 12256 13932
rect 10183 13892 12256 13920
rect 10183 13889 10195 13892
rect 10137 13883 10195 13889
rect 12250 13880 12256 13892
rect 12308 13880 12314 13932
rect 14274 13920 14280 13932
rect 14235 13892 14280 13920
rect 14274 13880 14280 13892
rect 14332 13880 14338 13932
rect 17310 13920 17316 13932
rect 17271 13892 17316 13920
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 2280 13824 2544 13852
rect 2280 13812 2286 13824
rect 2774 13812 2780 13864
rect 2832 13852 2838 13864
rect 4157 13855 4215 13861
rect 4157 13852 4169 13855
rect 2832 13824 4169 13852
rect 2832 13812 2838 13824
rect 4157 13821 4169 13824
rect 4203 13821 4215 13855
rect 4157 13815 4215 13821
rect 8665 13855 8723 13861
rect 8665 13821 8677 13855
rect 8711 13852 8723 13855
rect 8938 13852 8944 13864
rect 8711 13824 8944 13852
rect 8711 13821 8723 13824
rect 8665 13815 8723 13821
rect 8938 13812 8944 13824
rect 8996 13812 9002 13864
rect 9953 13855 10011 13861
rect 9953 13821 9965 13855
rect 9999 13852 10011 13855
rect 10318 13852 10324 13864
rect 9999 13824 10324 13852
rect 9999 13821 10011 13824
rect 9953 13815 10011 13821
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 11146 13812 11152 13864
rect 11204 13852 11210 13864
rect 11974 13852 11980 13864
rect 11204 13824 11980 13852
rect 11204 13812 11210 13824
rect 11974 13812 11980 13824
rect 12032 13852 12038 13864
rect 13998 13852 14004 13864
rect 12032 13824 14004 13852
rect 12032 13812 12038 13824
rect 13998 13812 14004 13824
rect 14056 13812 14062 13864
rect 17589 13855 17647 13861
rect 17589 13821 17601 13855
rect 17635 13852 17647 13855
rect 17862 13852 17868 13864
rect 17635 13824 17868 13852
rect 17635 13821 17647 13824
rect 17589 13815 17647 13821
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 18046 13852 18052 13864
rect 18007 13824 18052 13852
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 18248 13861 18276 13960
rect 19242 13880 19248 13932
rect 19300 13920 19306 13932
rect 19300 13892 19840 13920
rect 19300 13880 19306 13892
rect 18233 13855 18291 13861
rect 18233 13821 18245 13855
rect 18279 13821 18291 13855
rect 18233 13815 18291 13821
rect 19518 13812 19524 13864
rect 19576 13861 19582 13864
rect 19576 13855 19625 13861
rect 19576 13821 19579 13855
rect 19613 13821 19625 13855
rect 19702 13852 19708 13864
rect 19663 13824 19708 13852
rect 19576 13815 19625 13821
rect 19576 13812 19582 13815
rect 19702 13812 19708 13824
rect 19760 13812 19766 13864
rect 19812 13852 19840 13892
rect 19981 13855 20039 13861
rect 19981 13852 19993 13855
rect 19812 13824 19993 13852
rect 19981 13821 19993 13824
rect 20027 13821 20039 13855
rect 19981 13815 20039 13821
rect 20714 13812 20720 13864
rect 20772 13852 20778 13864
rect 20901 13855 20959 13861
rect 20901 13852 20913 13855
rect 20772 13824 20913 13852
rect 20772 13812 20778 13824
rect 20901 13821 20913 13824
rect 20947 13852 20959 13855
rect 20990 13852 20996 13864
rect 20947 13824 20996 13852
rect 20947 13821 20959 13824
rect 20901 13815 20959 13821
rect 20990 13812 20996 13824
rect 21048 13812 21054 13864
rect 2317 13787 2375 13793
rect 2317 13753 2329 13787
rect 2363 13784 2375 13787
rect 5626 13784 5632 13796
rect 2363 13756 5632 13784
rect 2363 13753 2375 13756
rect 2317 13747 2375 13753
rect 5626 13744 5632 13756
rect 5684 13744 5690 13796
rect 10686 13784 10692 13796
rect 9692 13756 10692 13784
rect 3510 13716 3516 13728
rect 3471 13688 3516 13716
rect 3510 13676 3516 13688
rect 3568 13676 3574 13728
rect 5442 13676 5448 13728
rect 5500 13716 5506 13728
rect 9692 13716 9720 13756
rect 10686 13744 10692 13756
rect 10744 13744 10750 13796
rect 15562 13784 15568 13796
rect 15502 13756 15568 13784
rect 15562 13744 15568 13756
rect 15620 13744 15626 13796
rect 19797 13787 19855 13793
rect 19797 13753 19809 13787
rect 19843 13784 19855 13787
rect 20254 13784 20260 13796
rect 19843 13756 20260 13784
rect 19843 13753 19855 13756
rect 19797 13747 19855 13753
rect 20254 13744 20260 13756
rect 20312 13744 20318 13796
rect 9858 13716 9864 13728
rect 5500 13688 9720 13716
rect 9819 13688 9864 13716
rect 5500 13676 5506 13688
rect 9858 13676 9864 13688
rect 9916 13676 9922 13728
rect 18417 13719 18475 13725
rect 18417 13685 18429 13719
rect 18463 13716 18475 13719
rect 18598 13716 18604 13728
rect 18463 13688 18604 13716
rect 18463 13685 18475 13688
rect 18417 13679 18475 13685
rect 18598 13676 18604 13688
rect 18656 13676 18662 13728
rect 1104 13626 21804 13648
rect 1104 13574 7882 13626
rect 7934 13574 7946 13626
rect 7998 13574 8010 13626
rect 8062 13574 8074 13626
rect 8126 13574 14782 13626
rect 14834 13574 14846 13626
rect 14898 13574 14910 13626
rect 14962 13574 14974 13626
rect 15026 13574 21804 13626
rect 1104 13552 21804 13574
rect 2314 13472 2320 13524
rect 2372 13512 2378 13524
rect 2409 13515 2467 13521
rect 2409 13512 2421 13515
rect 2372 13484 2421 13512
rect 2372 13472 2378 13484
rect 2409 13481 2421 13484
rect 2455 13481 2467 13515
rect 2774 13512 2780 13524
rect 2409 13475 2467 13481
rect 2746 13472 2780 13512
rect 2832 13512 2838 13524
rect 3145 13515 3203 13521
rect 3145 13512 3157 13515
rect 2832 13484 3157 13512
rect 2832 13472 2838 13484
rect 3145 13481 3157 13484
rect 3191 13481 3203 13515
rect 3145 13475 3203 13481
rect 4617 13515 4675 13521
rect 4617 13481 4629 13515
rect 4663 13512 4675 13515
rect 6733 13515 6791 13521
rect 6733 13512 6745 13515
rect 4663 13484 6745 13512
rect 4663 13481 4675 13484
rect 4617 13475 4675 13481
rect 6733 13481 6745 13484
rect 6779 13481 6791 13515
rect 6733 13475 6791 13481
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 7742 13512 7748 13524
rect 6972 13484 7748 13512
rect 6972 13472 6978 13484
rect 7742 13472 7748 13484
rect 7800 13512 7806 13524
rect 8297 13515 8355 13521
rect 8297 13512 8309 13515
rect 7800 13484 8309 13512
rect 7800 13472 7806 13484
rect 8297 13481 8309 13484
rect 8343 13481 8355 13515
rect 9858 13512 9864 13524
rect 9819 13484 9864 13512
rect 8297 13475 8355 13481
rect 9858 13472 9864 13484
rect 9916 13472 9922 13524
rect 15013 13515 15071 13521
rect 15013 13481 15025 13515
rect 15059 13512 15071 13515
rect 15102 13512 15108 13524
rect 15059 13484 15108 13512
rect 15059 13481 15071 13484
rect 15013 13475 15071 13481
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 15562 13512 15568 13524
rect 15523 13484 15568 13512
rect 15562 13472 15568 13484
rect 15620 13472 15626 13524
rect 1946 13336 1952 13388
rect 2004 13376 2010 13388
rect 2041 13379 2099 13385
rect 2041 13376 2053 13379
rect 2004 13348 2053 13376
rect 2004 13336 2010 13348
rect 2041 13345 2053 13348
rect 2087 13345 2099 13379
rect 2041 13339 2099 13345
rect 2409 13379 2467 13385
rect 2409 13345 2421 13379
rect 2455 13376 2467 13379
rect 2746 13376 2774 13472
rect 4246 13404 4252 13456
rect 4304 13444 4310 13456
rect 4709 13447 4767 13453
rect 4709 13444 4721 13447
rect 4304 13416 4721 13444
rect 4304 13404 4310 13416
rect 4709 13413 4721 13416
rect 4755 13413 4767 13447
rect 4709 13407 4767 13413
rect 7300 13416 8432 13444
rect 7300 13388 7328 13416
rect 3326 13376 3332 13388
rect 2455 13348 2774 13376
rect 3287 13348 3332 13376
rect 2455 13345 2467 13348
rect 2409 13339 2467 13345
rect 3326 13336 3332 13348
rect 3384 13336 3390 13388
rect 5813 13379 5871 13385
rect 5813 13345 5825 13379
rect 5859 13376 5871 13379
rect 6454 13376 6460 13388
rect 5859 13348 6460 13376
rect 5859 13345 5871 13348
rect 5813 13339 5871 13345
rect 6454 13336 6460 13348
rect 6512 13336 6518 13388
rect 6638 13336 6644 13388
rect 6696 13376 6702 13388
rect 6917 13379 6975 13385
rect 6917 13376 6929 13379
rect 6696 13348 6929 13376
rect 6696 13336 6702 13348
rect 6917 13345 6929 13348
rect 6963 13345 6975 13379
rect 6917 13339 6975 13345
rect 7101 13379 7159 13385
rect 7101 13345 7113 13379
rect 7147 13376 7159 13379
rect 7282 13376 7288 13388
rect 7147 13348 7288 13376
rect 7147 13345 7159 13348
rect 7101 13339 7159 13345
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 8404 13385 8432 13416
rect 14550 13404 14556 13456
rect 14608 13444 14614 13456
rect 16206 13444 16212 13456
rect 14608 13416 15148 13444
rect 16167 13416 16212 13444
rect 14608 13404 14614 13416
rect 7561 13379 7619 13385
rect 7561 13345 7573 13379
rect 7607 13345 7619 13379
rect 7561 13339 7619 13345
rect 8389 13379 8447 13385
rect 8389 13345 8401 13379
rect 8435 13345 8447 13379
rect 10042 13376 10048 13388
rect 8389 13339 8447 13345
rect 8496 13348 10048 13376
rect 4798 13308 4804 13320
rect 4759 13280 4804 13308
rect 4798 13268 4804 13280
rect 4856 13308 4862 13320
rect 5442 13308 5448 13320
rect 4856 13280 5448 13308
rect 4856 13268 4862 13280
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 5626 13308 5632 13320
rect 5587 13280 5632 13308
rect 5626 13268 5632 13280
rect 5684 13268 5690 13320
rect 5905 13311 5963 13317
rect 5905 13277 5917 13311
rect 5951 13277 5963 13311
rect 5905 13271 5963 13277
rect 5997 13311 6055 13317
rect 5997 13277 6009 13311
rect 6043 13277 6055 13311
rect 5997 13271 6055 13277
rect 6089 13311 6147 13317
rect 6089 13277 6101 13311
rect 6135 13308 6147 13311
rect 6656 13308 6684 13336
rect 6135 13280 6684 13308
rect 6135 13277 6147 13280
rect 6089 13271 6147 13277
rect 3602 13132 3608 13184
rect 3660 13172 3666 13184
rect 4249 13175 4307 13181
rect 4249 13172 4261 13175
rect 3660 13144 4261 13172
rect 3660 13132 3666 13144
rect 4249 13141 4261 13144
rect 4295 13141 4307 13175
rect 5920 13172 5948 13271
rect 6012 13240 6040 13271
rect 6822 13268 6828 13320
rect 6880 13308 6886 13320
rect 7576 13308 7604 13339
rect 8496 13308 8524 13348
rect 10042 13336 10048 13348
rect 10100 13336 10106 13388
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13376 10195 13379
rect 10502 13376 10508 13388
rect 10183 13348 10508 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 10502 13336 10508 13348
rect 10560 13336 10566 13388
rect 10597 13379 10655 13385
rect 10597 13345 10609 13379
rect 10643 13345 10655 13379
rect 10597 13339 10655 13345
rect 6880 13280 8524 13308
rect 6880 13268 6886 13280
rect 9490 13268 9496 13320
rect 9548 13308 9554 13320
rect 10612 13308 10640 13339
rect 11146 13336 11152 13388
rect 11204 13376 11210 13388
rect 15120 13385 15148 13416
rect 16206 13404 16212 13416
rect 16264 13404 16270 13456
rect 17310 13404 17316 13456
rect 17368 13404 17374 13456
rect 17954 13444 17960 13456
rect 17915 13416 17960 13444
rect 17954 13404 17960 13416
rect 18012 13404 18018 13456
rect 12253 13379 12311 13385
rect 12253 13376 12265 13379
rect 11204 13348 12265 13376
rect 11204 13336 11210 13348
rect 12253 13345 12265 13348
rect 12299 13345 12311 13379
rect 12253 13339 12311 13345
rect 14921 13379 14979 13385
rect 14921 13345 14933 13379
rect 14967 13345 14979 13379
rect 14921 13339 14979 13345
rect 15105 13379 15163 13385
rect 15105 13345 15117 13379
rect 15151 13345 15163 13379
rect 15746 13376 15752 13388
rect 15707 13348 15752 13376
rect 15105 13339 15163 13345
rect 9548 13280 10640 13308
rect 9548 13268 9554 13280
rect 10778 13268 10784 13320
rect 10836 13308 10842 13320
rect 11977 13311 12035 13317
rect 11977 13308 11989 13311
rect 10836 13280 11989 13308
rect 10836 13268 10842 13280
rect 11977 13277 11989 13280
rect 12023 13277 12035 13311
rect 12158 13308 12164 13320
rect 12119 13280 12164 13308
rect 11977 13271 12035 13277
rect 6012 13212 7052 13240
rect 6730 13172 6736 13184
rect 5920 13144 6736 13172
rect 4249 13135 4307 13141
rect 6730 13132 6736 13144
rect 6788 13132 6794 13184
rect 6914 13172 6920 13184
rect 6875 13144 6920 13172
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 7024 13172 7052 13212
rect 7098 13200 7104 13252
rect 7156 13240 7162 13252
rect 7653 13243 7711 13249
rect 7653 13240 7665 13243
rect 7156 13212 7665 13240
rect 7156 13200 7162 13212
rect 7653 13209 7665 13212
rect 7699 13240 7711 13243
rect 9398 13240 9404 13252
rect 7699 13212 9404 13240
rect 7699 13209 7711 13212
rect 7653 13203 7711 13209
rect 9398 13200 9404 13212
rect 9456 13200 9462 13252
rect 9582 13200 9588 13252
rect 9640 13240 9646 13252
rect 10229 13243 10287 13249
rect 10229 13240 10241 13243
rect 9640 13212 10241 13240
rect 9640 13200 9646 13212
rect 10229 13209 10241 13212
rect 10275 13209 10287 13243
rect 10229 13203 10287 13209
rect 10321 13243 10379 13249
rect 10321 13209 10333 13243
rect 10367 13240 10379 13243
rect 10594 13240 10600 13252
rect 10367 13212 10600 13240
rect 10367 13209 10379 13212
rect 10321 13203 10379 13209
rect 10594 13200 10600 13212
rect 10652 13200 10658 13252
rect 11992 13240 12020 13271
rect 12158 13268 12164 13280
rect 12216 13268 12222 13320
rect 14936 13308 14964 13339
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 16224 13308 16252 13404
rect 17954 13308 17960 13320
rect 14936 13280 16252 13308
rect 16776 13280 17960 13308
rect 12894 13240 12900 13252
rect 11992 13212 12900 13240
rect 12894 13200 12900 13212
rect 12952 13240 12958 13252
rect 13538 13240 13544 13252
rect 12952 13212 13544 13240
rect 12952 13200 12958 13212
rect 13538 13200 13544 13212
rect 13596 13200 13602 13252
rect 13998 13200 14004 13252
rect 14056 13240 14062 13252
rect 16776 13240 16804 13280
rect 17954 13268 17960 13280
rect 18012 13308 18018 13320
rect 18233 13311 18291 13317
rect 18233 13308 18245 13311
rect 18012 13280 18245 13308
rect 18012 13268 18018 13280
rect 18233 13277 18245 13280
rect 18279 13308 18291 13311
rect 19334 13308 19340 13320
rect 18279 13280 19340 13308
rect 18279 13277 18291 13280
rect 18233 13271 18291 13277
rect 19334 13268 19340 13280
rect 19392 13268 19398 13320
rect 14056 13212 16804 13240
rect 14056 13200 14062 13212
rect 7558 13172 7564 13184
rect 7024 13144 7564 13172
rect 7558 13132 7564 13144
rect 7616 13132 7622 13184
rect 10134 13132 10140 13184
rect 10192 13172 10198 13184
rect 10413 13175 10471 13181
rect 10413 13172 10425 13175
rect 10192 13144 10425 13172
rect 10192 13132 10198 13144
rect 10413 13141 10425 13144
rect 10459 13141 10471 13175
rect 12618 13172 12624 13184
rect 12579 13144 12624 13172
rect 10413 13135 10471 13141
rect 12618 13132 12624 13144
rect 12676 13132 12682 13184
rect 1104 13082 21804 13104
rect 1104 13030 4432 13082
rect 4484 13030 4496 13082
rect 4548 13030 4560 13082
rect 4612 13030 4624 13082
rect 4676 13030 11332 13082
rect 11384 13030 11396 13082
rect 11448 13030 11460 13082
rect 11512 13030 11524 13082
rect 11576 13030 18232 13082
rect 18284 13030 18296 13082
rect 18348 13030 18360 13082
rect 18412 13030 18424 13082
rect 18476 13030 21804 13082
rect 1104 13008 21804 13030
rect 1486 12968 1492 12980
rect 1447 12940 1492 12968
rect 1486 12928 1492 12940
rect 1544 12928 1550 12980
rect 3145 12971 3203 12977
rect 3145 12937 3157 12971
rect 3191 12968 3203 12971
rect 3326 12968 3332 12980
rect 3191 12940 3332 12968
rect 3191 12937 3203 12940
rect 3145 12931 3203 12937
rect 3326 12928 3332 12940
rect 3384 12968 3390 12980
rect 3973 12971 4031 12977
rect 3973 12968 3985 12971
rect 3384 12940 3985 12968
rect 3384 12928 3390 12940
rect 3973 12937 3985 12940
rect 4019 12937 4031 12971
rect 9398 12968 9404 12980
rect 9359 12940 9404 12968
rect 3973 12931 4031 12937
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 10686 12928 10692 12980
rect 10744 12968 10750 12980
rect 10744 12940 12480 12968
rect 10744 12928 10750 12940
rect 6638 12860 6644 12912
rect 6696 12900 6702 12912
rect 9769 12903 9827 12909
rect 6696 12872 9720 12900
rect 6696 12860 6702 12872
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 3602 12832 3608 12844
rect 2823 12804 3608 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 3602 12792 3608 12804
rect 3660 12792 3666 12844
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 9490 12832 9496 12844
rect 7156 12804 8524 12832
rect 9451 12804 9496 12832
rect 7156 12792 7162 12804
rect 3973 12767 4031 12773
rect 3973 12733 3985 12767
rect 4019 12764 4031 12767
rect 4338 12764 4344 12776
rect 4019 12736 4344 12764
rect 4019 12733 4031 12736
rect 3973 12727 4031 12733
rect 4338 12724 4344 12736
rect 4396 12724 4402 12776
rect 6822 12764 6828 12776
rect 6783 12736 6828 12764
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 7009 12767 7067 12773
rect 7009 12733 7021 12767
rect 7055 12764 7067 12767
rect 7558 12764 7564 12776
rect 7055 12736 7564 12764
rect 7055 12733 7067 12736
rect 7009 12727 7067 12733
rect 7558 12724 7564 12736
rect 7616 12724 7622 12776
rect 7650 12724 7656 12776
rect 7708 12764 7714 12776
rect 8205 12767 8263 12773
rect 8205 12764 8217 12767
rect 7708 12736 8217 12764
rect 7708 12724 7714 12736
rect 8205 12733 8217 12736
rect 8251 12733 8263 12767
rect 8205 12727 8263 12733
rect 1581 12699 1639 12705
rect 1581 12665 1593 12699
rect 1627 12696 1639 12699
rect 2406 12696 2412 12708
rect 1627 12668 2412 12696
rect 1627 12665 1639 12668
rect 1581 12659 1639 12665
rect 2406 12656 2412 12668
rect 2464 12656 2470 12708
rect 3142 12696 3148 12708
rect 3103 12668 3148 12696
rect 3142 12656 3148 12668
rect 3200 12656 3206 12708
rect 8386 12696 8392 12708
rect 8347 12668 8392 12696
rect 8386 12656 8392 12668
rect 8444 12656 8450 12708
rect 8496 12696 8524 12804
rect 9490 12792 9496 12804
rect 9548 12792 9554 12844
rect 9692 12832 9720 12872
rect 9769 12869 9781 12903
rect 9815 12900 9827 12903
rect 11146 12900 11152 12912
rect 9815 12872 11152 12900
rect 9815 12869 9827 12872
rect 9769 12863 9827 12869
rect 11146 12860 11152 12872
rect 11204 12860 11210 12912
rect 10778 12832 10784 12844
rect 9692 12804 10784 12832
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 12250 12832 12256 12844
rect 12211 12804 12256 12832
rect 12250 12792 12256 12804
rect 12308 12792 12314 12844
rect 12452 12841 12480 12940
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12801 12495 12835
rect 12437 12795 12495 12801
rect 17954 12792 17960 12844
rect 18012 12832 18018 12844
rect 18233 12835 18291 12841
rect 18233 12832 18245 12835
rect 18012 12804 18245 12832
rect 18012 12792 18018 12804
rect 18233 12801 18245 12804
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 18509 12835 18567 12841
rect 18509 12801 18521 12835
rect 18555 12832 18567 12835
rect 18598 12832 18604 12844
rect 18555 12804 18604 12832
rect 18555 12801 18567 12804
rect 18509 12795 18567 12801
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 20254 12832 20260 12844
rect 20215 12804 20260 12832
rect 20254 12792 20260 12804
rect 20312 12792 20318 12844
rect 8573 12767 8631 12773
rect 8573 12733 8585 12767
rect 8619 12764 8631 12767
rect 9398 12764 9404 12776
rect 8619 12736 9404 12764
rect 8619 12733 8631 12736
rect 8573 12727 8631 12733
rect 9398 12724 9404 12736
rect 9456 12724 9462 12776
rect 10594 12724 10600 12776
rect 10652 12764 10658 12776
rect 10965 12767 11023 12773
rect 10965 12764 10977 12767
rect 10652 12736 10977 12764
rect 10652 12724 10658 12736
rect 10965 12733 10977 12736
rect 11011 12733 11023 12767
rect 11146 12764 11152 12776
rect 11107 12736 11152 12764
rect 10965 12727 11023 12733
rect 11146 12724 11152 12736
rect 11204 12724 11210 12776
rect 13538 12764 13544 12776
rect 13499 12736 13544 12764
rect 13538 12724 13544 12736
rect 13596 12724 13602 12776
rect 21082 12764 21088 12776
rect 21043 12736 21088 12764
rect 21082 12724 21088 12736
rect 21140 12724 21146 12776
rect 9582 12696 9588 12708
rect 8496 12668 9588 12696
rect 9582 12656 9588 12668
rect 9640 12656 9646 12708
rect 12158 12656 12164 12708
rect 12216 12696 12222 12708
rect 13357 12699 13415 12705
rect 13357 12696 13369 12699
rect 12216 12668 13369 12696
rect 12216 12656 12222 12668
rect 13357 12665 13369 12668
rect 13403 12665 13415 12699
rect 19978 12696 19984 12708
rect 19734 12668 19984 12696
rect 13357 12659 13415 12665
rect 19978 12656 19984 12668
rect 20036 12656 20042 12708
rect 7101 12631 7159 12637
rect 7101 12597 7113 12631
rect 7147 12628 7159 12631
rect 7282 12628 7288 12640
rect 7147 12600 7288 12628
rect 7147 12597 7159 12600
rect 7101 12591 7159 12597
rect 7282 12588 7288 12600
rect 7340 12628 7346 12640
rect 10962 12628 10968 12640
rect 7340 12600 10968 12628
rect 7340 12588 7346 12600
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 11057 12631 11115 12637
rect 11057 12597 11069 12631
rect 11103 12628 11115 12631
rect 12342 12628 12348 12640
rect 11103 12600 12348 12628
rect 11103 12597 11115 12600
rect 11057 12591 11115 12597
rect 12342 12588 12348 12600
rect 12400 12588 12406 12640
rect 12526 12588 12532 12640
rect 12584 12628 12590 12640
rect 12894 12628 12900 12640
rect 12584 12600 12629 12628
rect 12855 12600 12900 12628
rect 12584 12588 12590 12600
rect 12894 12588 12900 12600
rect 12952 12588 12958 12640
rect 13725 12631 13783 12637
rect 13725 12597 13737 12631
rect 13771 12628 13783 12631
rect 15102 12628 15108 12640
rect 13771 12600 15108 12628
rect 13771 12597 13783 12600
rect 13725 12591 13783 12597
rect 15102 12588 15108 12600
rect 15160 12588 15166 12640
rect 20898 12628 20904 12640
rect 20859 12600 20904 12628
rect 20898 12588 20904 12600
rect 20956 12588 20962 12640
rect 1104 12538 21804 12560
rect 1104 12486 7882 12538
rect 7934 12486 7946 12538
rect 7998 12486 8010 12538
rect 8062 12486 8074 12538
rect 8126 12486 14782 12538
rect 14834 12486 14846 12538
rect 14898 12486 14910 12538
rect 14962 12486 14974 12538
rect 15026 12486 21804 12538
rect 1104 12464 21804 12486
rect 4338 12424 4344 12436
rect 4299 12396 4344 12424
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 11885 12427 11943 12433
rect 11885 12393 11897 12427
rect 11931 12424 11943 12427
rect 12158 12424 12164 12436
rect 11931 12396 12164 12424
rect 11931 12393 11943 12396
rect 11885 12387 11943 12393
rect 12158 12384 12164 12396
rect 12216 12384 12222 12436
rect 12250 12384 12256 12436
rect 12308 12384 12314 12436
rect 12345 12427 12403 12433
rect 12345 12393 12357 12427
rect 12391 12424 12403 12427
rect 12526 12424 12532 12436
rect 12391 12396 12532 12424
rect 12391 12393 12403 12396
rect 12345 12387 12403 12393
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 15102 12424 15108 12436
rect 15063 12396 15108 12424
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 15197 12427 15255 12433
rect 15197 12393 15209 12427
rect 15243 12424 15255 12427
rect 15838 12424 15844 12436
rect 15243 12396 15844 12424
rect 15243 12393 15255 12396
rect 15197 12387 15255 12393
rect 15838 12384 15844 12396
rect 15896 12384 15902 12436
rect 17310 12424 17316 12436
rect 17271 12396 17316 12424
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 19978 12424 19984 12436
rect 19939 12396 19984 12424
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 6086 12356 6092 12368
rect 6047 12328 6092 12356
rect 6086 12316 6092 12328
rect 6144 12316 6150 12368
rect 6454 12356 6460 12368
rect 6367 12328 6460 12356
rect 6454 12316 6460 12328
rect 6512 12356 6518 12368
rect 11701 12359 11759 12365
rect 11701 12356 11713 12359
rect 6512 12328 11713 12356
rect 6512 12316 6518 12328
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 4249 12291 4307 12297
rect 4249 12288 4261 12291
rect 4212 12260 4261 12288
rect 4212 12248 4218 12260
rect 4249 12257 4261 12260
rect 4295 12257 4307 12291
rect 4249 12251 4307 12257
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12288 6331 12291
rect 7098 12288 7104 12300
rect 6319 12260 7104 12288
rect 6319 12257 6331 12260
rect 6273 12251 6331 12257
rect 7098 12248 7104 12260
rect 7156 12248 7162 12300
rect 7208 12297 7236 12328
rect 10428 12300 10456 12328
rect 11701 12325 11713 12328
rect 11747 12325 11759 12359
rect 12268 12356 12296 12384
rect 11701 12319 11759 12325
rect 12084 12328 12296 12356
rect 7193 12291 7251 12297
rect 7193 12257 7205 12291
rect 7239 12257 7251 12291
rect 7193 12251 7251 12257
rect 7742 12248 7748 12300
rect 7800 12288 7806 12300
rect 7929 12291 7987 12297
rect 7929 12288 7941 12291
rect 7800 12260 7941 12288
rect 7800 12248 7806 12260
rect 7929 12257 7941 12260
rect 7975 12257 7987 12291
rect 7929 12251 7987 12257
rect 8205 12291 8263 12297
rect 8205 12257 8217 12291
rect 8251 12257 8263 12291
rect 8205 12251 8263 12257
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 7837 12223 7895 12229
rect 7837 12220 7849 12223
rect 7524 12192 7849 12220
rect 7524 12180 7530 12192
rect 7837 12189 7849 12192
rect 7883 12189 7895 12223
rect 8220 12220 8248 12251
rect 9490 12248 9496 12300
rect 9548 12288 9554 12300
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 9548 12260 10057 12288
rect 9548 12248 9554 12260
rect 10045 12257 10057 12260
rect 10091 12257 10103 12291
rect 10226 12288 10232 12300
rect 10187 12260 10232 12288
rect 10045 12251 10103 12257
rect 10226 12248 10232 12260
rect 10284 12248 10290 12300
rect 10410 12288 10416 12300
rect 10323 12260 10416 12288
rect 10410 12248 10416 12260
rect 10468 12248 10474 12300
rect 10505 12291 10563 12297
rect 10505 12257 10517 12291
rect 10551 12288 10563 12291
rect 10594 12288 10600 12300
rect 10551 12260 10600 12288
rect 10551 12257 10563 12260
rect 10505 12251 10563 12257
rect 10594 12248 10600 12260
rect 10652 12248 10658 12300
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12288 11483 12291
rect 11517 12291 11575 12297
rect 11517 12288 11529 12291
rect 11471 12260 11529 12288
rect 11471 12257 11483 12260
rect 11425 12251 11483 12257
rect 11517 12257 11529 12260
rect 11563 12257 11575 12291
rect 11517 12251 11575 12257
rect 9858 12220 9864 12232
rect 8220 12192 9864 12220
rect 7837 12183 7895 12189
rect 9858 12180 9864 12192
rect 9916 12220 9922 12232
rect 10321 12223 10379 12229
rect 10321 12220 10333 12223
rect 9916 12192 10333 12220
rect 9916 12180 9922 12192
rect 10321 12189 10333 12192
rect 10367 12220 10379 12223
rect 10686 12220 10692 12232
rect 10367 12192 10692 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 12084 12220 12112 12328
rect 12158 12248 12164 12300
rect 12216 12288 12222 12300
rect 12529 12291 12587 12297
rect 12529 12288 12541 12291
rect 12216 12260 12541 12288
rect 12216 12248 12222 12260
rect 12529 12257 12541 12260
rect 12575 12257 12587 12291
rect 12529 12251 12587 12257
rect 12618 12248 12624 12300
rect 12676 12288 12682 12300
rect 12676 12260 12721 12288
rect 12676 12248 12682 12260
rect 15746 12248 15752 12300
rect 15804 12288 15810 12300
rect 17497 12291 17555 12297
rect 17497 12288 17509 12291
rect 15804 12260 17509 12288
rect 15804 12248 15810 12260
rect 17497 12257 17509 12260
rect 17543 12288 17555 12291
rect 20165 12291 20223 12297
rect 20165 12288 20177 12291
rect 17543 12260 20177 12288
rect 17543 12257 17555 12260
rect 17497 12251 17555 12257
rect 20165 12257 20177 12260
rect 20211 12288 20223 12291
rect 20622 12288 20628 12300
rect 20211 12260 20628 12288
rect 20211 12257 20223 12260
rect 20165 12251 20223 12257
rect 20622 12248 20628 12260
rect 20680 12248 20686 12300
rect 20806 12248 20812 12300
rect 20864 12288 20870 12300
rect 20901 12291 20959 12297
rect 20901 12288 20913 12291
rect 20864 12260 20913 12288
rect 20864 12248 20870 12260
rect 20901 12257 20913 12260
rect 20947 12257 20959 12291
rect 20901 12251 20959 12257
rect 12342 12220 12348 12232
rect 12084 12192 12348 12220
rect 12342 12180 12348 12192
rect 12400 12220 12406 12232
rect 15289 12223 15347 12229
rect 15289 12220 15301 12223
rect 12400 12192 15301 12220
rect 12400 12180 12406 12192
rect 15289 12189 15301 12192
rect 15335 12220 15347 12223
rect 15562 12220 15568 12232
rect 15335 12192 15568 12220
rect 15335 12189 15347 12192
rect 15289 12183 15347 12189
rect 15562 12180 15568 12192
rect 15620 12180 15626 12232
rect 10781 12155 10839 12161
rect 10781 12121 10793 12155
rect 10827 12152 10839 12155
rect 15838 12152 15844 12164
rect 10827 12124 15844 12152
rect 10827 12121 10839 12124
rect 10781 12115 10839 12121
rect 15838 12112 15844 12124
rect 15896 12112 15902 12164
rect 7285 12087 7343 12093
rect 7285 12053 7297 12087
rect 7331 12084 7343 12087
rect 7374 12084 7380 12096
rect 7331 12056 7380 12084
rect 7331 12053 7343 12056
rect 7285 12047 7343 12053
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 10502 12044 10508 12096
rect 10560 12084 10566 12096
rect 10962 12084 10968 12096
rect 10560 12056 10968 12084
rect 10560 12044 10566 12056
rect 10962 12044 10968 12056
rect 11020 12084 11026 12096
rect 11425 12087 11483 12093
rect 11425 12084 11437 12087
rect 11020 12056 11437 12084
rect 11020 12044 11026 12056
rect 11425 12053 11437 12056
rect 11471 12053 11483 12087
rect 11425 12047 11483 12053
rect 14090 12044 14096 12096
rect 14148 12084 14154 12096
rect 14737 12087 14795 12093
rect 14737 12084 14749 12087
rect 14148 12056 14749 12084
rect 14148 12044 14154 12056
rect 14737 12053 14749 12056
rect 14783 12053 14795 12087
rect 20714 12084 20720 12096
rect 20675 12056 20720 12084
rect 14737 12047 14795 12053
rect 20714 12044 20720 12056
rect 20772 12044 20778 12096
rect 1104 11994 21804 12016
rect 1104 11942 4432 11994
rect 4484 11942 4496 11994
rect 4548 11942 4560 11994
rect 4612 11942 4624 11994
rect 4676 11942 11332 11994
rect 11384 11942 11396 11994
rect 11448 11942 11460 11994
rect 11512 11942 11524 11994
rect 11576 11942 18232 11994
rect 18284 11942 18296 11994
rect 18348 11942 18360 11994
rect 18412 11942 18424 11994
rect 18476 11942 21804 11994
rect 1104 11920 21804 11942
rect 5813 11883 5871 11889
rect 5813 11849 5825 11883
rect 5859 11880 5871 11883
rect 7282 11880 7288 11892
rect 5859 11852 7288 11880
rect 5859 11849 5871 11852
rect 5813 11843 5871 11849
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 2222 11812 2228 11824
rect 1964 11784 2228 11812
rect 1964 11753 1992 11784
rect 2222 11772 2228 11784
rect 2280 11772 2286 11824
rect 3697 11815 3755 11821
rect 3697 11781 3709 11815
rect 3743 11812 3755 11815
rect 4154 11812 4160 11824
rect 3743 11784 4160 11812
rect 3743 11781 3755 11784
rect 3697 11775 3755 11781
rect 4154 11772 4160 11784
rect 4212 11772 4218 11824
rect 13262 11812 13268 11824
rect 13223 11784 13268 11812
rect 13262 11772 13268 11784
rect 13320 11772 13326 11824
rect 1949 11747 2007 11753
rect 1949 11713 1961 11747
rect 1995 11713 2007 11747
rect 1949 11707 2007 11713
rect 2038 11704 2044 11756
rect 2096 11744 2102 11756
rect 2133 11747 2191 11753
rect 2133 11744 2145 11747
rect 2096 11716 2145 11744
rect 2096 11704 2102 11716
rect 2133 11713 2145 11716
rect 2179 11713 2191 11747
rect 2133 11707 2191 11713
rect 3142 11704 3148 11756
rect 3200 11744 3206 11756
rect 3513 11747 3571 11753
rect 3513 11744 3525 11747
rect 3200 11716 3525 11744
rect 3200 11704 3206 11716
rect 3513 11713 3525 11716
rect 3559 11744 3571 11747
rect 3786 11744 3792 11756
rect 3559 11716 3792 11744
rect 3559 11713 3571 11716
rect 3513 11707 3571 11713
rect 3786 11704 3792 11716
rect 3844 11744 3850 11756
rect 6825 11747 6883 11753
rect 3844 11716 4568 11744
rect 3844 11704 3850 11716
rect 3881 11679 3939 11685
rect 3881 11645 3893 11679
rect 3927 11676 3939 11679
rect 4338 11676 4344 11688
rect 3927 11648 4344 11676
rect 3927 11645 3939 11648
rect 3881 11639 3939 11645
rect 4338 11636 4344 11648
rect 4396 11636 4402 11688
rect 4540 11685 4568 11716
rect 6825 11713 6837 11747
rect 6871 11744 6883 11747
rect 7006 11744 7012 11756
rect 6871 11716 7012 11744
rect 6871 11713 6883 11716
rect 6825 11707 6883 11713
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 8849 11747 8907 11753
rect 8849 11713 8861 11747
rect 8895 11744 8907 11747
rect 9858 11744 9864 11756
rect 8895 11716 9864 11744
rect 8895 11713 8907 11716
rect 8849 11707 8907 11713
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 10410 11704 10416 11756
rect 10468 11744 10474 11756
rect 10597 11747 10655 11753
rect 10597 11744 10609 11747
rect 10468 11716 10609 11744
rect 10468 11704 10474 11716
rect 10597 11713 10609 11716
rect 10643 11713 10655 11747
rect 12894 11744 12900 11756
rect 12855 11716 12900 11744
rect 10597 11707 10655 11713
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 15562 11744 15568 11756
rect 13464 11716 14044 11744
rect 15523 11716 15568 11744
rect 4525 11679 4583 11685
rect 4525 11645 4537 11679
rect 4571 11645 4583 11679
rect 4525 11639 4583 11645
rect 5629 11679 5687 11685
rect 5629 11645 5641 11679
rect 5675 11645 5687 11679
rect 5629 11639 5687 11645
rect 5905 11679 5963 11685
rect 5905 11645 5917 11679
rect 5951 11676 5963 11679
rect 7098 11676 7104 11688
rect 5951 11648 7104 11676
rect 5951 11645 5963 11648
rect 5905 11639 5963 11645
rect 2225 11611 2283 11617
rect 2225 11577 2237 11611
rect 2271 11608 2283 11611
rect 5445 11611 5503 11617
rect 5445 11608 5457 11611
rect 2271 11580 5457 11608
rect 2271 11577 2283 11580
rect 2225 11571 2283 11577
rect 5445 11577 5457 11580
rect 5491 11577 5503 11611
rect 5644 11608 5672 11639
rect 7098 11636 7104 11648
rect 7156 11636 7162 11688
rect 8478 11636 8484 11688
rect 8536 11676 8542 11688
rect 8573 11679 8631 11685
rect 8573 11676 8585 11679
rect 8536 11648 8585 11676
rect 8536 11636 8542 11648
rect 8573 11645 8585 11648
rect 8619 11645 8631 11679
rect 8573 11639 8631 11645
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 6638 11608 6644 11620
rect 5644 11580 6644 11608
rect 5445 11571 5503 11577
rect 6638 11568 6644 11580
rect 6696 11608 6702 11620
rect 7009 11611 7067 11617
rect 7009 11608 7021 11611
rect 6696 11580 7021 11608
rect 6696 11568 6702 11580
rect 7009 11577 7021 11580
rect 7055 11577 7067 11611
rect 7009 11571 7067 11577
rect 7193 11611 7251 11617
rect 7193 11577 7205 11611
rect 7239 11608 7251 11611
rect 7558 11608 7564 11620
rect 7239 11580 7564 11608
rect 7239 11577 7251 11580
rect 7193 11571 7251 11577
rect 2590 11540 2596 11552
rect 2551 11512 2596 11540
rect 2590 11500 2596 11512
rect 2648 11500 2654 11552
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 4341 11543 4399 11549
rect 4341 11540 4353 11543
rect 4304 11512 4353 11540
rect 4304 11500 4310 11512
rect 4341 11509 4353 11512
rect 4387 11509 4399 11543
rect 7024 11540 7052 11571
rect 7558 11568 7564 11580
rect 7616 11608 7622 11620
rect 8680 11608 8708 11639
rect 8754 11636 8760 11688
rect 8812 11676 8818 11688
rect 8812 11648 8857 11676
rect 8812 11636 8818 11648
rect 10686 11636 10692 11688
rect 10744 11676 10750 11688
rect 10873 11679 10931 11685
rect 10744 11648 10789 11676
rect 10744 11636 10750 11648
rect 10873 11645 10885 11679
rect 10919 11645 10931 11679
rect 10873 11639 10931 11645
rect 11057 11679 11115 11685
rect 11057 11645 11069 11679
rect 11103 11676 11115 11679
rect 13464 11676 13492 11716
rect 13906 11676 13912 11688
rect 11103 11648 13492 11676
rect 13556 11648 13912 11676
rect 11103 11645 11115 11648
rect 11057 11639 11115 11645
rect 9674 11608 9680 11620
rect 7616 11580 9680 11608
rect 7616 11568 7622 11580
rect 9674 11568 9680 11580
rect 9732 11568 9738 11620
rect 10778 11568 10784 11620
rect 10836 11608 10842 11620
rect 10888 11608 10916 11639
rect 10836 11580 10916 11608
rect 13265 11611 13323 11617
rect 10836 11568 10842 11580
rect 13265 11577 13277 11611
rect 13311 11577 13323 11611
rect 13265 11571 13323 11577
rect 7742 11540 7748 11552
rect 7024 11512 7748 11540
rect 4341 11503 4399 11509
rect 7742 11500 7748 11512
rect 7800 11500 7806 11552
rect 9033 11543 9091 11549
rect 9033 11509 9045 11543
rect 9079 11540 9091 11543
rect 9122 11540 9128 11552
rect 9079 11512 9128 11540
rect 9079 11509 9091 11512
rect 9033 11503 9091 11509
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 13280 11540 13308 11571
rect 13556 11540 13584 11648
rect 13906 11636 13912 11648
rect 13964 11636 13970 11688
rect 14016 11608 14044 11716
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 15654 11704 15660 11756
rect 15712 11744 15718 11756
rect 20806 11744 20812 11756
rect 15712 11716 20812 11744
rect 15712 11704 15718 11716
rect 20806 11704 20812 11716
rect 20864 11704 20870 11756
rect 15749 11679 15807 11685
rect 15749 11645 15761 11679
rect 15795 11676 15807 11679
rect 20714 11676 20720 11688
rect 15795 11648 20720 11676
rect 15795 11645 15807 11648
rect 15749 11639 15807 11645
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 20898 11676 20904 11688
rect 20859 11648 20904 11676
rect 20898 11636 20904 11648
rect 20956 11636 20962 11688
rect 15841 11611 15899 11617
rect 15841 11608 15853 11611
rect 14016 11580 15853 11608
rect 15841 11577 15853 11580
rect 15887 11577 15899 11611
rect 15841 11571 15899 11577
rect 13722 11540 13728 11552
rect 13280 11512 13584 11540
rect 13683 11512 13728 11540
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 16209 11543 16267 11549
rect 16209 11509 16221 11543
rect 16255 11540 16267 11543
rect 16390 11540 16396 11552
rect 16255 11512 16396 11540
rect 16255 11509 16267 11512
rect 16209 11503 16267 11509
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 20714 11540 20720 11552
rect 20675 11512 20720 11540
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 1104 11450 21804 11472
rect 1104 11398 7882 11450
rect 7934 11398 7946 11450
rect 7998 11398 8010 11450
rect 8062 11398 8074 11450
rect 8126 11398 14782 11450
rect 14834 11398 14846 11450
rect 14898 11398 14910 11450
rect 14962 11398 14974 11450
rect 15026 11398 21804 11450
rect 1104 11376 21804 11398
rect 4154 11296 4160 11348
rect 4212 11336 4218 11348
rect 4249 11339 4307 11345
rect 4249 11336 4261 11339
rect 4212 11308 4261 11336
rect 4212 11296 4218 11308
rect 4249 11305 4261 11308
rect 4295 11305 4307 11339
rect 4249 11299 4307 11305
rect 5537 11339 5595 11345
rect 5537 11305 5549 11339
rect 5583 11336 5595 11339
rect 6365 11339 6423 11345
rect 6365 11336 6377 11339
rect 5583 11308 6377 11336
rect 5583 11305 5595 11308
rect 5537 11299 5595 11305
rect 6365 11305 6377 11308
rect 6411 11305 6423 11339
rect 6365 11299 6423 11305
rect 6454 11296 6460 11348
rect 6512 11336 6518 11348
rect 11241 11339 11299 11345
rect 11241 11336 11253 11339
rect 6512 11308 11253 11336
rect 6512 11296 6518 11308
rect 11241 11305 11253 11308
rect 11287 11305 11299 11339
rect 11241 11299 11299 11305
rect 11609 11339 11667 11345
rect 11609 11305 11621 11339
rect 11655 11336 11667 11339
rect 12158 11336 12164 11348
rect 11655 11308 12164 11336
rect 11655 11305 11667 11308
rect 11609 11299 11667 11305
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 13262 11336 13268 11348
rect 13223 11308 13268 11336
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 15105 11339 15163 11345
rect 15105 11305 15117 11339
rect 15151 11336 15163 11339
rect 15933 11339 15991 11345
rect 15933 11336 15945 11339
rect 15151 11308 15945 11336
rect 15151 11305 15163 11308
rect 15105 11299 15163 11305
rect 15933 11305 15945 11308
rect 15979 11336 15991 11339
rect 16761 11339 16819 11345
rect 16761 11336 16773 11339
rect 15979 11308 16773 11336
rect 15979 11305 15991 11308
rect 15933 11299 15991 11305
rect 16761 11305 16773 11308
rect 16807 11305 16819 11339
rect 16761 11299 16819 11305
rect 5629 11271 5687 11277
rect 5629 11237 5641 11271
rect 5675 11268 5687 11271
rect 10321 11271 10379 11277
rect 5675 11240 10272 11268
rect 5675 11237 5687 11240
rect 5629 11231 5687 11237
rect 2225 11203 2283 11209
rect 2225 11169 2237 11203
rect 2271 11200 2283 11203
rect 2314 11200 2320 11212
rect 2271 11172 2320 11200
rect 2271 11169 2283 11172
rect 2225 11163 2283 11169
rect 2314 11160 2320 11172
rect 2372 11160 2378 11212
rect 4246 11200 4252 11212
rect 4207 11172 4252 11200
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 4338 11160 4344 11212
rect 4396 11200 4402 11212
rect 4617 11203 4675 11209
rect 4617 11200 4629 11203
rect 4396 11172 4629 11200
rect 4396 11160 4402 11172
rect 4617 11169 4629 11172
rect 4663 11200 4675 11203
rect 6454 11200 6460 11212
rect 4663 11172 6460 11200
rect 4663 11169 4675 11172
rect 4617 11163 4675 11169
rect 6454 11160 6460 11172
rect 6512 11160 6518 11212
rect 6549 11203 6607 11209
rect 6549 11169 6561 11203
rect 6595 11200 6607 11203
rect 6914 11200 6920 11212
rect 6595 11172 6920 11200
rect 6595 11169 6607 11172
rect 6549 11163 6607 11169
rect 6914 11160 6920 11172
rect 6972 11200 6978 11212
rect 7745 11203 7803 11209
rect 7745 11200 7757 11203
rect 6972 11172 7757 11200
rect 6972 11160 6978 11172
rect 7745 11169 7757 11172
rect 7791 11169 7803 11203
rect 7745 11163 7803 11169
rect 7834 11160 7840 11212
rect 7892 11200 7898 11212
rect 8389 11203 8447 11209
rect 7892 11172 7937 11200
rect 7892 11160 7898 11172
rect 8389 11169 8401 11203
rect 8435 11169 8447 11203
rect 8389 11163 8447 11169
rect 5442 11092 5448 11144
rect 5500 11132 5506 11144
rect 5721 11135 5779 11141
rect 5721 11132 5733 11135
rect 5500 11104 5733 11132
rect 5500 11092 5506 11104
rect 5721 11101 5733 11104
rect 5767 11101 5779 11135
rect 5721 11095 5779 11101
rect 6086 11092 6092 11144
rect 6144 11132 6150 11144
rect 6638 11132 6644 11144
rect 6144 11104 6644 11132
rect 6144 11092 6150 11104
rect 6638 11092 6644 11104
rect 6696 11092 6702 11144
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11132 6883 11135
rect 7006 11132 7012 11144
rect 6871 11104 7012 11132
rect 6871 11101 6883 11104
rect 6825 11095 6883 11101
rect 4154 11024 4160 11076
rect 4212 11064 4218 11076
rect 5169 11067 5227 11073
rect 5169 11064 5181 11067
rect 4212 11036 5181 11064
rect 4212 11024 4218 11036
rect 5169 11033 5181 11036
rect 5215 11033 5227 11067
rect 6748 11064 6776 11095
rect 7006 11092 7012 11104
rect 7064 11092 7070 11144
rect 7190 11092 7196 11144
rect 7248 11132 7254 11144
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 7248 11104 7389 11132
rect 7248 11092 7254 11104
rect 7377 11101 7389 11104
rect 7423 11101 7435 11135
rect 7558 11132 7564 11144
rect 7519 11104 7564 11132
rect 7377 11095 7435 11101
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 7650 11092 7656 11144
rect 7708 11132 7714 11144
rect 7708 11104 7753 11132
rect 7708 11092 7714 11104
rect 7024 11064 7052 11092
rect 8404 11064 8432 11163
rect 8754 11160 8760 11212
rect 8812 11200 8818 11212
rect 9306 11200 9312 11212
rect 8812 11172 9312 11200
rect 8812 11160 8818 11172
rect 9306 11160 9312 11172
rect 9364 11200 9370 11212
rect 9585 11203 9643 11209
rect 9585 11200 9597 11203
rect 9364 11172 9597 11200
rect 9364 11160 9370 11172
rect 9585 11169 9597 11172
rect 9631 11169 9643 11203
rect 9585 11163 9643 11169
rect 9674 11160 9680 11212
rect 9732 11200 9738 11212
rect 9858 11200 9864 11212
rect 9732 11172 9777 11200
rect 9819 11172 9864 11200
rect 9732 11160 9738 11172
rect 9858 11160 9864 11172
rect 9916 11160 9922 11212
rect 10244 11200 10272 11240
rect 10321 11237 10333 11271
rect 10367 11268 10379 11271
rect 10502 11268 10508 11280
rect 10367 11240 10508 11268
rect 10367 11237 10379 11240
rect 10321 11231 10379 11237
rect 10502 11228 10508 11240
rect 10560 11268 10566 11280
rect 10686 11268 10692 11280
rect 10560 11240 10692 11268
rect 10560 11228 10566 11240
rect 10686 11228 10692 11240
rect 10744 11228 10750 11280
rect 20714 11268 20720 11280
rect 10796 11240 20720 11268
rect 10796 11200 10824 11240
rect 20714 11228 20720 11240
rect 20772 11228 20778 11280
rect 10244 11172 10824 11200
rect 11701 11203 11759 11209
rect 11701 11169 11713 11203
rect 11747 11200 11759 11203
rect 12894 11200 12900 11212
rect 11747 11172 12756 11200
rect 12855 11172 12900 11200
rect 11747 11169 11759 11172
rect 11701 11163 11759 11169
rect 11885 11135 11943 11141
rect 11885 11101 11897 11135
rect 11931 11132 11943 11135
rect 12342 11132 12348 11144
rect 11931 11104 12348 11132
rect 11931 11101 11943 11104
rect 11885 11095 11943 11101
rect 12342 11092 12348 11104
rect 12400 11132 12406 11144
rect 12728 11132 12756 11172
rect 12894 11160 12900 11172
rect 12952 11160 12958 11212
rect 13265 11203 13323 11209
rect 13265 11169 13277 11203
rect 13311 11200 13323 11203
rect 13722 11200 13728 11212
rect 13311 11172 13728 11200
rect 13311 11169 13323 11172
rect 13265 11163 13323 11169
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 15565 11203 15623 11209
rect 15565 11169 15577 11203
rect 15611 11200 15623 11203
rect 16390 11200 16396 11212
rect 15611 11172 16396 11200
rect 15611 11169 15623 11172
rect 15565 11163 15623 11169
rect 16390 11160 16396 11172
rect 16448 11160 16454 11212
rect 16758 11200 16764 11212
rect 16671 11172 16764 11200
rect 16758 11160 16764 11172
rect 16816 11200 16822 11212
rect 17405 11203 17463 11209
rect 17405 11200 17417 11203
rect 16816 11172 17417 11200
rect 16816 11160 16822 11172
rect 17405 11169 17417 11172
rect 17451 11169 17463 11203
rect 17405 11163 17463 11169
rect 15654 11132 15660 11144
rect 12400 11092 12434 11132
rect 12728 11104 15660 11132
rect 15654 11092 15660 11104
rect 15712 11092 15718 11144
rect 6748 11036 6960 11064
rect 7024 11036 8432 11064
rect 12406 11064 12434 11092
rect 13170 11064 13176 11076
rect 12406 11036 13176 11064
rect 5169 11027 5227 11033
rect 2409 10999 2467 11005
rect 2409 10965 2421 10999
rect 2455 10996 2467 10999
rect 2682 10996 2688 11008
rect 2455 10968 2688 10996
rect 2455 10965 2467 10968
rect 2409 10959 2467 10965
rect 2682 10956 2688 10968
rect 2740 10956 2746 11008
rect 6932 10996 6960 11036
rect 13170 11024 13176 11036
rect 13228 11024 13234 11076
rect 15933 11067 15991 11073
rect 15933 11033 15945 11067
rect 15979 11064 15991 11067
rect 17221 11067 17279 11073
rect 17221 11064 17233 11067
rect 15979 11036 17233 11064
rect 15979 11033 15991 11036
rect 15933 11027 15991 11033
rect 17221 11033 17233 11036
rect 17267 11033 17279 11067
rect 17221 11027 17279 11033
rect 7098 10996 7104 11008
rect 6932 10968 7104 10996
rect 7098 10956 7104 10968
rect 7156 10996 7162 11008
rect 7650 10996 7656 11008
rect 7156 10968 7656 10996
rect 7156 10956 7162 10968
rect 7650 10956 7656 10968
rect 7708 10956 7714 11008
rect 8478 10996 8484 11008
rect 8439 10968 8484 10996
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 15010 10996 15016 11008
rect 14971 10968 15016 10996
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 1104 10906 21804 10928
rect 1104 10854 4432 10906
rect 4484 10854 4496 10906
rect 4548 10854 4560 10906
rect 4612 10854 4624 10906
rect 4676 10854 11332 10906
rect 11384 10854 11396 10906
rect 11448 10854 11460 10906
rect 11512 10854 11524 10906
rect 11576 10854 18232 10906
rect 18284 10854 18296 10906
rect 18348 10854 18360 10906
rect 18412 10854 18424 10906
rect 18476 10854 21804 10906
rect 1104 10832 21804 10854
rect 3786 10792 3792 10804
rect 3747 10764 3792 10792
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7466 10792 7472 10804
rect 6972 10764 7472 10792
rect 6972 10752 6978 10764
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 8205 10795 8263 10801
rect 8205 10761 8217 10795
rect 8251 10792 8263 10795
rect 8386 10792 8392 10804
rect 8251 10764 8392 10792
rect 8251 10761 8263 10764
rect 8205 10755 8263 10761
rect 8386 10752 8392 10764
rect 8444 10752 8450 10804
rect 8478 10752 8484 10804
rect 8536 10792 8542 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8536 10764 8953 10792
rect 8536 10752 8542 10764
rect 8941 10761 8953 10764
rect 8987 10792 8999 10795
rect 9677 10795 9735 10801
rect 9677 10792 9689 10795
rect 8987 10764 9689 10792
rect 8987 10761 8999 10764
rect 8941 10755 8999 10761
rect 9677 10761 9689 10764
rect 9723 10761 9735 10795
rect 9677 10755 9735 10761
rect 10410 10752 10416 10804
rect 10468 10792 10474 10804
rect 10505 10795 10563 10801
rect 10505 10792 10517 10795
rect 10468 10764 10517 10792
rect 10468 10752 10474 10764
rect 10505 10761 10517 10764
rect 10551 10761 10563 10795
rect 10505 10755 10563 10761
rect 13906 10752 13912 10804
rect 13964 10792 13970 10804
rect 14461 10795 14519 10801
rect 14461 10792 14473 10795
rect 13964 10764 14473 10792
rect 13964 10752 13970 10764
rect 14461 10761 14473 10764
rect 14507 10761 14519 10795
rect 14461 10755 14519 10761
rect 20717 10795 20775 10801
rect 20717 10761 20729 10795
rect 20763 10792 20775 10795
rect 20806 10792 20812 10804
rect 20763 10764 20812 10792
rect 20763 10761 20775 10764
rect 20717 10755 20775 10761
rect 20806 10752 20812 10764
rect 20864 10752 20870 10804
rect 7374 10684 7380 10736
rect 7432 10724 7438 10736
rect 9033 10727 9091 10733
rect 7432 10696 8892 10724
rect 7432 10684 7438 10696
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10656 1915 10659
rect 2590 10656 2596 10668
rect 1903 10628 2596 10656
rect 1903 10625 1915 10628
rect 1857 10619 1915 10625
rect 2590 10616 2596 10628
rect 2648 10656 2654 10668
rect 3053 10659 3111 10665
rect 3053 10656 3065 10659
rect 2648 10628 3065 10656
rect 2648 10616 2654 10628
rect 3053 10625 3065 10628
rect 3099 10625 3111 10659
rect 3053 10619 3111 10625
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10656 8447 10659
rect 8478 10656 8484 10668
rect 8435 10628 8484 10656
rect 8435 10625 8447 10628
rect 8389 10619 8447 10625
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10588 2283 10591
rect 2314 10588 2320 10600
rect 2271 10560 2320 10588
rect 2271 10557 2283 10560
rect 2225 10551 2283 10557
rect 2314 10548 2320 10560
rect 2372 10548 2378 10600
rect 2682 10588 2688 10600
rect 2643 10560 2688 10588
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 3973 10591 4031 10597
rect 3973 10557 3985 10591
rect 4019 10588 4031 10591
rect 4062 10588 4068 10600
rect 4019 10560 4068 10588
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 8113 10591 8171 10597
rect 8113 10557 8125 10591
rect 8159 10588 8171 10591
rect 8754 10588 8760 10600
rect 8159 10560 8760 10588
rect 8159 10557 8171 10560
rect 8113 10551 8171 10557
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 8864 10597 8892 10696
rect 9033 10693 9045 10727
rect 9079 10724 9091 10727
rect 9079 10696 10824 10724
rect 9079 10693 9091 10696
rect 9033 10687 9091 10693
rect 9122 10656 9128 10668
rect 9083 10628 9128 10656
rect 9122 10616 9128 10628
rect 9180 10656 9186 10668
rect 9861 10659 9919 10665
rect 9861 10656 9873 10659
rect 9180 10628 9873 10656
rect 9180 10616 9186 10628
rect 9861 10625 9873 10628
rect 9907 10625 9919 10659
rect 10796 10656 10824 10696
rect 10870 10684 10876 10736
rect 10928 10724 10934 10736
rect 10928 10696 13492 10724
rect 10928 10684 10934 10696
rect 13170 10656 13176 10668
rect 10796 10628 12572 10656
rect 13131 10628 13176 10656
rect 9861 10619 9919 10625
rect 8849 10591 8907 10597
rect 8849 10557 8861 10591
rect 8895 10557 8907 10591
rect 8849 10551 8907 10557
rect 9585 10591 9643 10597
rect 9585 10557 9597 10591
rect 9631 10557 9643 10591
rect 11698 10588 11704 10600
rect 9585 10551 9643 10557
rect 9876 10560 11704 10588
rect 8478 10480 8484 10532
rect 8536 10520 8542 10532
rect 9600 10520 9628 10551
rect 9876 10529 9904 10560
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 10502 10529 10508 10532
rect 8536 10492 9628 10520
rect 9861 10523 9919 10529
rect 8536 10480 8542 10492
rect 9861 10489 9873 10523
rect 9907 10489 9919 10523
rect 9861 10483 9919 10489
rect 10484 10523 10508 10529
rect 10484 10489 10496 10523
rect 10484 10483 10508 10489
rect 10502 10480 10508 10483
rect 10560 10480 10566 10532
rect 10689 10523 10747 10529
rect 10689 10489 10701 10523
rect 10735 10520 10747 10523
rect 10962 10520 10968 10532
rect 10735 10492 10968 10520
rect 10735 10489 10747 10492
rect 10689 10483 10747 10489
rect 10962 10480 10968 10492
rect 11020 10480 11026 10532
rect 12544 10520 12572 10628
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 13354 10656 13360 10668
rect 13315 10628 13360 10656
rect 13354 10616 13360 10628
rect 13412 10616 13418 10668
rect 12621 10591 12679 10597
rect 12621 10557 12633 10591
rect 12667 10588 12679 10591
rect 13262 10588 13268 10600
rect 12667 10560 13268 10588
rect 12667 10557 12679 10560
rect 12621 10551 12679 10557
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 13464 10597 13492 10696
rect 15010 10684 15016 10736
rect 15068 10724 15074 10736
rect 15105 10727 15163 10733
rect 15105 10724 15117 10727
rect 15068 10696 15117 10724
rect 15068 10684 15074 10696
rect 15105 10693 15117 10696
rect 15151 10693 15163 10727
rect 15105 10687 15163 10693
rect 16117 10727 16175 10733
rect 16117 10693 16129 10727
rect 16163 10693 16175 10727
rect 16117 10687 16175 10693
rect 13449 10591 13507 10597
rect 13449 10557 13461 10591
rect 13495 10557 13507 10591
rect 13449 10551 13507 10557
rect 14645 10591 14703 10597
rect 14645 10557 14657 10591
rect 14691 10588 14703 10591
rect 15470 10588 15476 10600
rect 14691 10560 15148 10588
rect 15431 10560 15476 10588
rect 14691 10557 14703 10560
rect 14645 10551 14703 10557
rect 12544 10492 14688 10520
rect 14660 10464 14688 10492
rect 2225 10455 2283 10461
rect 2225 10421 2237 10455
rect 2271 10452 2283 10455
rect 2685 10455 2743 10461
rect 2685 10452 2697 10455
rect 2271 10424 2697 10452
rect 2271 10421 2283 10424
rect 2225 10415 2283 10421
rect 2685 10421 2697 10424
rect 2731 10452 2743 10455
rect 2958 10452 2964 10464
rect 2731 10424 2964 10452
rect 2731 10421 2743 10424
rect 2685 10415 2743 10421
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 8389 10455 8447 10461
rect 8389 10421 8401 10455
rect 8435 10452 8447 10455
rect 8662 10452 8668 10464
rect 8435 10424 8668 10452
rect 8435 10421 8447 10424
rect 8389 10415 8447 10421
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 10321 10455 10379 10461
rect 10321 10421 10333 10455
rect 10367 10452 10379 10455
rect 10594 10452 10600 10464
rect 10367 10424 10600 10452
rect 10367 10421 10379 10424
rect 10321 10415 10379 10421
rect 10594 10412 10600 10424
rect 10652 10412 10658 10464
rect 12526 10452 12532 10464
rect 12487 10424 12532 10452
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 13814 10452 13820 10464
rect 13775 10424 13820 10452
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 14642 10412 14648 10464
rect 14700 10412 14706 10464
rect 15120 10461 15148 10560
rect 15470 10548 15476 10560
rect 15528 10588 15534 10600
rect 15933 10591 15991 10597
rect 15933 10588 15945 10591
rect 15528 10560 15945 10588
rect 15528 10548 15534 10560
rect 15933 10557 15945 10560
rect 15979 10557 15991 10591
rect 15933 10551 15991 10557
rect 15105 10455 15163 10461
rect 15105 10421 15117 10455
rect 15151 10452 15163 10455
rect 16132 10452 16160 10687
rect 20898 10588 20904 10600
rect 20859 10560 20904 10588
rect 20898 10548 20904 10560
rect 20956 10548 20962 10600
rect 16301 10523 16359 10529
rect 16301 10489 16313 10523
rect 16347 10520 16359 10523
rect 16758 10520 16764 10532
rect 16347 10492 16764 10520
rect 16347 10489 16359 10492
rect 16301 10483 16359 10489
rect 16758 10480 16764 10492
rect 16816 10480 16822 10532
rect 15151 10424 16160 10452
rect 15151 10421 15163 10424
rect 15105 10415 15163 10421
rect 1104 10362 21804 10384
rect 1104 10310 7882 10362
rect 7934 10310 7946 10362
rect 7998 10310 8010 10362
rect 8062 10310 8074 10362
rect 8126 10310 14782 10362
rect 14834 10310 14846 10362
rect 14898 10310 14910 10362
rect 14962 10310 14974 10362
rect 15026 10310 21804 10362
rect 1104 10288 21804 10310
rect 1486 10248 1492 10260
rect 1447 10220 1492 10248
rect 1486 10208 1492 10220
rect 1544 10208 1550 10260
rect 2314 10248 2320 10260
rect 2275 10220 2320 10248
rect 2314 10208 2320 10220
rect 2372 10208 2378 10260
rect 2958 10248 2964 10260
rect 2919 10220 2964 10248
rect 2958 10208 2964 10220
rect 3016 10208 3022 10260
rect 5902 10208 5908 10260
rect 5960 10248 5966 10260
rect 5997 10251 6055 10257
rect 5997 10248 6009 10251
rect 5960 10220 6009 10248
rect 5960 10208 5966 10220
rect 5997 10217 6009 10220
rect 6043 10217 6055 10251
rect 5997 10211 6055 10217
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7101 10251 7159 10257
rect 7101 10248 7113 10251
rect 7064 10220 7113 10248
rect 7064 10208 7070 10220
rect 7101 10217 7113 10220
rect 7147 10217 7159 10251
rect 7101 10211 7159 10217
rect 7469 10251 7527 10257
rect 7469 10217 7481 10251
rect 7515 10248 7527 10251
rect 15470 10248 15476 10260
rect 7515 10220 15476 10248
rect 7515 10217 7527 10220
rect 7469 10211 7527 10217
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10112 1639 10115
rect 1762 10112 1768 10124
rect 1627 10084 1768 10112
rect 1627 10081 1639 10084
rect 1581 10075 1639 10081
rect 1762 10072 1768 10084
rect 1820 10072 1826 10124
rect 2501 10115 2559 10121
rect 2501 10081 2513 10115
rect 2547 10112 2559 10115
rect 2682 10112 2688 10124
rect 2547 10084 2688 10112
rect 2547 10081 2559 10084
rect 2501 10075 2559 10081
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 5905 10115 5963 10121
rect 5905 10081 5917 10115
rect 5951 10112 5963 10115
rect 6914 10112 6920 10124
rect 5951 10084 6920 10112
rect 5951 10081 5963 10084
rect 5905 10075 5963 10081
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 7116 10112 7144 10211
rect 15470 10208 15476 10220
rect 15528 10208 15534 10260
rect 15933 10251 15991 10257
rect 15933 10217 15945 10251
rect 15979 10248 15991 10251
rect 16758 10248 16764 10260
rect 15979 10220 16764 10248
rect 15979 10217 15991 10220
rect 15933 10211 15991 10217
rect 16758 10208 16764 10220
rect 16816 10208 16822 10260
rect 20898 10248 20904 10260
rect 20859 10220 20904 10248
rect 20898 10208 20904 10220
rect 20956 10208 20962 10260
rect 8846 10180 8852 10192
rect 8404 10152 8852 10180
rect 8404 10121 8432 10152
rect 8846 10140 8852 10152
rect 8904 10180 8910 10192
rect 10870 10180 10876 10192
rect 8904 10152 10876 10180
rect 8904 10140 8910 10152
rect 10870 10140 10876 10152
rect 10928 10140 10934 10192
rect 12989 10183 13047 10189
rect 12989 10149 13001 10183
rect 13035 10180 13047 10183
rect 13906 10180 13912 10192
rect 13035 10152 13912 10180
rect 13035 10149 13047 10152
rect 12989 10143 13047 10149
rect 13906 10140 13912 10152
rect 13964 10140 13970 10192
rect 8113 10115 8171 10121
rect 8113 10112 8125 10115
rect 7116 10084 8125 10112
rect 8113 10081 8125 10084
rect 8159 10081 8171 10115
rect 8113 10075 8171 10081
rect 8389 10115 8447 10121
rect 8389 10081 8401 10115
rect 8435 10081 8447 10115
rect 8389 10075 8447 10081
rect 9398 10072 9404 10124
rect 9456 10112 9462 10124
rect 9493 10115 9551 10121
rect 9493 10112 9505 10115
rect 9456 10084 9505 10112
rect 9456 10072 9462 10084
rect 9493 10081 9505 10084
rect 9539 10081 9551 10115
rect 10502 10112 10508 10124
rect 10463 10084 10508 10112
rect 9493 10075 9551 10081
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 10686 10112 10692 10124
rect 10647 10084 10692 10112
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 15746 10112 15752 10124
rect 15707 10084 15752 10112
rect 15746 10072 15752 10084
rect 15804 10072 15810 10124
rect 21082 10112 21088 10124
rect 21043 10084 21088 10112
rect 21082 10072 21088 10084
rect 21140 10072 21146 10124
rect 5442 10004 5448 10056
rect 5500 10044 5506 10056
rect 6089 10047 6147 10053
rect 6089 10044 6101 10047
rect 5500 10016 6101 10044
rect 5500 10004 5506 10016
rect 6089 10013 6101 10016
rect 6135 10044 6147 10047
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6135 10016 6837 10044
rect 6135 10013 6147 10016
rect 6089 10007 6147 10013
rect 3050 9908 3056 9920
rect 3011 9880 3056 9908
rect 3050 9868 3056 9880
rect 3108 9868 3114 9920
rect 5534 9908 5540 9920
rect 5495 9880 5540 9908
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 6564 9908 6592 10016
rect 6825 10013 6837 10016
rect 6871 10013 6883 10047
rect 7006 10044 7012 10056
rect 6967 10016 7012 10044
rect 6825 10007 6883 10013
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10013 8263 10047
rect 8205 10007 8263 10013
rect 8297 10047 8355 10053
rect 8297 10013 8309 10047
rect 8343 10044 8355 10047
rect 9582 10044 9588 10056
rect 8343 10016 9588 10044
rect 8343 10013 8355 10016
rect 8297 10007 8355 10013
rect 6638 9936 6644 9988
rect 6696 9976 6702 9988
rect 7650 9976 7656 9988
rect 6696 9948 7656 9976
rect 6696 9936 6702 9948
rect 7650 9936 7656 9948
rect 7708 9976 7714 9988
rect 8220 9976 8248 10007
rect 9582 10004 9588 10016
rect 9640 10044 9646 10056
rect 10413 10047 10471 10053
rect 10413 10044 10425 10047
rect 9640 10016 10425 10044
rect 9640 10004 9646 10016
rect 10413 10013 10425 10016
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 12621 10047 12679 10053
rect 12621 10013 12633 10047
rect 12667 10044 12679 10047
rect 12710 10044 12716 10056
rect 12667 10016 12716 10044
rect 12667 10013 12679 10016
rect 12621 10007 12679 10013
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 7708 9948 8248 9976
rect 10873 9979 10931 9985
rect 7708 9936 7714 9948
rect 10873 9945 10885 9979
rect 10919 9976 10931 9979
rect 12802 9976 12808 9988
rect 10919 9948 12808 9976
rect 10919 9945 10931 9948
rect 10873 9939 10931 9945
rect 12802 9936 12808 9948
rect 12860 9936 12866 9988
rect 7098 9908 7104 9920
rect 6564 9880 7104 9908
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 7558 9868 7564 9920
rect 7616 9908 7622 9920
rect 7929 9911 7987 9917
rect 7929 9908 7941 9911
rect 7616 9880 7941 9908
rect 7616 9868 7622 9880
rect 7929 9877 7941 9880
rect 7975 9877 7987 9911
rect 9582 9908 9588 9920
rect 9543 9880 9588 9908
rect 7929 9871 7987 9877
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 12894 9908 12900 9920
rect 12855 9880 12900 9908
rect 12894 9868 12900 9880
rect 12952 9868 12958 9920
rect 1104 9818 21804 9840
rect 1104 9766 4432 9818
rect 4484 9766 4496 9818
rect 4548 9766 4560 9818
rect 4612 9766 4624 9818
rect 4676 9766 11332 9818
rect 11384 9766 11396 9818
rect 11448 9766 11460 9818
rect 11512 9766 11524 9818
rect 11576 9766 18232 9818
rect 18284 9766 18296 9818
rect 18348 9766 18360 9818
rect 18412 9766 18424 9818
rect 18476 9766 21804 9818
rect 1104 9744 21804 9766
rect 6914 9664 6920 9716
rect 6972 9704 6978 9716
rect 8846 9704 8852 9716
rect 6972 9676 8708 9704
rect 8807 9676 8852 9704
rect 6972 9664 6978 9676
rect 8680 9636 8708 9676
rect 8846 9664 8852 9676
rect 8904 9664 8910 9716
rect 10045 9707 10103 9713
rect 8956 9676 9536 9704
rect 8956 9636 8984 9676
rect 8680 9608 8984 9636
rect 2685 9571 2743 9577
rect 2685 9537 2697 9571
rect 2731 9568 2743 9571
rect 3050 9568 3056 9580
rect 2731 9540 3056 9568
rect 2731 9537 2743 9540
rect 2685 9531 2743 9537
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 4154 9568 4160 9580
rect 4115 9540 4160 9568
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 5534 9568 5540 9580
rect 5495 9540 5540 9568
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 2038 9460 2044 9512
rect 2096 9500 2102 9512
rect 2133 9503 2191 9509
rect 2133 9500 2145 9503
rect 2096 9472 2145 9500
rect 2096 9460 2102 9472
rect 2133 9469 2145 9472
rect 2179 9469 2191 9503
rect 2133 9463 2191 9469
rect 5169 9503 5227 9509
rect 5169 9469 5181 9503
rect 5215 9500 5227 9503
rect 5718 9500 5724 9512
rect 5215 9472 5724 9500
rect 5215 9469 5227 9472
rect 5169 9463 5227 9469
rect 5718 9460 5724 9472
rect 5776 9460 5782 9512
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9469 7527 9503
rect 7650 9500 7656 9512
rect 7611 9472 7656 9500
rect 7469 9463 7527 9469
rect 2593 9435 2651 9441
rect 2593 9401 2605 9435
rect 2639 9432 2651 9435
rect 2866 9432 2872 9444
rect 2639 9404 2872 9432
rect 2639 9401 2651 9404
rect 2593 9395 2651 9401
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 4617 9435 4675 9441
rect 4617 9432 4629 9435
rect 4120 9404 4629 9432
rect 4120 9392 4126 9404
rect 4617 9401 4629 9404
rect 4663 9401 4675 9435
rect 4617 9395 4675 9401
rect 4709 9435 4767 9441
rect 4709 9401 4721 9435
rect 4755 9432 4767 9435
rect 4890 9432 4896 9444
rect 4755 9404 4896 9432
rect 4755 9401 4767 9404
rect 4709 9395 4767 9401
rect 4890 9392 4896 9404
rect 4948 9392 4954 9444
rect 7484 9432 7512 9463
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 7745 9503 7803 9509
rect 7745 9469 7757 9503
rect 7791 9500 7803 9503
rect 8941 9503 8999 9509
rect 7791 9472 8892 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 8662 9432 8668 9444
rect 7484 9404 8668 9432
rect 8662 9392 8668 9404
rect 8720 9392 8726 9444
rect 8864 9432 8892 9472
rect 8941 9469 8953 9503
rect 8987 9500 8999 9503
rect 9122 9500 9128 9512
rect 8987 9472 9128 9500
rect 8987 9469 8999 9472
rect 8941 9463 8999 9469
rect 9122 9460 9128 9472
rect 9180 9460 9186 9512
rect 9508 9500 9536 9676
rect 10045 9673 10057 9707
rect 10091 9704 10103 9707
rect 10502 9704 10508 9716
rect 10091 9676 10508 9704
rect 10091 9673 10103 9676
rect 10045 9667 10103 9673
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 15473 9707 15531 9713
rect 15473 9673 15485 9707
rect 15519 9704 15531 9707
rect 15746 9704 15752 9716
rect 15519 9676 15752 9704
rect 15519 9673 15531 9676
rect 15473 9667 15531 9673
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 12526 9596 12532 9648
rect 12584 9636 12590 9648
rect 12897 9639 12955 9645
rect 12897 9636 12909 9639
rect 12584 9608 12909 9636
rect 12584 9596 12590 9608
rect 12897 9605 12909 9608
rect 12943 9605 12955 9639
rect 12897 9599 12955 9605
rect 9582 9528 9588 9580
rect 9640 9568 9646 9580
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 9640 9540 10149 9568
rect 9640 9528 9646 9540
rect 10137 9537 10149 9540
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 13814 9528 13820 9580
rect 13872 9568 13878 9580
rect 15102 9568 15108 9580
rect 13872 9540 15108 9568
rect 13872 9528 13878 9540
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 9861 9503 9919 9509
rect 9861 9500 9873 9503
rect 9508 9472 9873 9500
rect 9861 9469 9873 9472
rect 9907 9500 9919 9503
rect 10686 9500 10692 9512
rect 9907 9472 10692 9500
rect 9907 9469 9919 9472
rect 9861 9463 9919 9469
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 10962 9460 10968 9512
rect 11020 9500 11026 9512
rect 12253 9503 12311 9509
rect 12253 9500 12265 9503
rect 11020 9472 12265 9500
rect 11020 9460 11026 9472
rect 12253 9469 12265 9472
rect 12299 9469 12311 9503
rect 12253 9463 12311 9469
rect 12710 9460 12716 9512
rect 12768 9500 12774 9512
rect 13265 9503 13323 9509
rect 13265 9500 13277 9503
rect 12768 9472 13277 9500
rect 12768 9460 12774 9472
rect 13265 9469 13277 9472
rect 13311 9469 13323 9503
rect 13265 9463 13323 9469
rect 9766 9432 9772 9444
rect 8864 9404 9772 9432
rect 9766 9392 9772 9404
rect 9824 9432 9830 9444
rect 10410 9432 10416 9444
rect 9824 9404 10416 9432
rect 9824 9392 9830 9404
rect 10410 9392 10416 9404
rect 10468 9432 10474 9444
rect 12069 9435 12127 9441
rect 12069 9432 12081 9435
rect 10468 9404 12081 9432
rect 10468 9392 10474 9404
rect 12069 9401 12081 9404
rect 12115 9401 12127 9435
rect 12069 9395 12127 9401
rect 15194 9392 15200 9444
rect 15252 9432 15258 9444
rect 15473 9435 15531 9441
rect 15473 9432 15485 9435
rect 15252 9404 15485 9432
rect 15252 9392 15258 9404
rect 15473 9401 15485 9404
rect 15519 9401 15531 9435
rect 15473 9395 15531 9401
rect 5169 9367 5227 9373
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 5258 9364 5264 9376
rect 5215 9336 5264 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 7282 9364 7288 9376
rect 7243 9336 7288 9364
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 9674 9364 9680 9376
rect 9635 9336 9680 9364
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 12434 9364 12440 9376
rect 12395 9336 12440 9364
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 12894 9364 12900 9376
rect 12855 9336 12900 9364
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 1104 9274 21804 9296
rect 1104 9222 7882 9274
rect 7934 9222 7946 9274
rect 7998 9222 8010 9274
rect 8062 9222 8074 9274
rect 8126 9222 14782 9274
rect 14834 9222 14846 9274
rect 14898 9222 14910 9274
rect 14962 9222 14974 9274
rect 15026 9222 21804 9274
rect 1104 9200 21804 9222
rect 2038 9160 2044 9172
rect 1999 9132 2044 9160
rect 2038 9120 2044 9132
rect 2096 9120 2102 9172
rect 2409 9163 2467 9169
rect 2409 9129 2421 9163
rect 2455 9160 2467 9163
rect 7282 9160 7288 9172
rect 2455 9132 7288 9160
rect 2455 9129 2467 9132
rect 2409 9123 2467 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 9953 9163 10011 9169
rect 9953 9129 9965 9163
rect 9999 9160 10011 9163
rect 10318 9160 10324 9172
rect 9999 9132 10324 9160
rect 9999 9129 10011 9132
rect 9953 9123 10011 9129
rect 10318 9120 10324 9132
rect 10376 9120 10382 9172
rect 12434 9120 12440 9172
rect 12492 9160 12498 9172
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 12492 9132 13093 9160
rect 12492 9120 12498 9132
rect 13081 9129 13093 9132
rect 13127 9129 13139 9163
rect 13081 9123 13139 9129
rect 15657 9163 15715 9169
rect 15657 9129 15669 9163
rect 15703 9160 15715 9163
rect 15746 9160 15752 9172
rect 15703 9132 15752 9160
rect 15703 9129 15715 9132
rect 15657 9123 15715 9129
rect 15746 9120 15752 9132
rect 15804 9120 15810 9172
rect 5718 9092 5724 9104
rect 4816 9064 5724 9092
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 8984 1458 9036
rect 4154 8984 4160 9036
rect 4212 9024 4218 9036
rect 4816 9033 4844 9064
rect 5718 9052 5724 9064
rect 5776 9092 5782 9104
rect 7193 9095 7251 9101
rect 7193 9092 7205 9095
rect 5776 9064 6132 9092
rect 5776 9052 5782 9064
rect 6104 9036 6132 9064
rect 6380 9064 7205 9092
rect 4249 9027 4307 9033
rect 4249 9024 4261 9027
rect 4212 8996 4261 9024
rect 4212 8984 4218 8996
rect 4249 8993 4261 8996
rect 4295 8993 4307 9027
rect 4249 8987 4307 8993
rect 4801 9027 4859 9033
rect 4801 8993 4813 9027
rect 4847 8993 4859 9027
rect 4801 8987 4859 8993
rect 4908 8996 5396 9024
rect 1670 8916 1676 8968
rect 1728 8956 1734 8968
rect 2501 8959 2559 8965
rect 2501 8956 2513 8959
rect 1728 8928 2513 8956
rect 1728 8916 1734 8928
rect 2501 8925 2513 8928
rect 2547 8925 2559 8959
rect 2501 8919 2559 8925
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8925 2743 8959
rect 2685 8919 2743 8925
rect 2700 8888 2728 8919
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 4617 8959 4675 8965
rect 4617 8956 4629 8959
rect 4120 8928 4629 8956
rect 4120 8916 4126 8928
rect 4617 8925 4629 8928
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 2700 8860 2774 8888
rect 1486 8780 1492 8832
rect 1544 8820 1550 8832
rect 1581 8823 1639 8829
rect 1581 8820 1593 8823
rect 1544 8792 1593 8820
rect 1544 8780 1550 8792
rect 1581 8789 1593 8792
rect 1627 8789 1639 8823
rect 2746 8820 2774 8860
rect 3694 8848 3700 8900
rect 3752 8888 3758 8900
rect 4908 8888 4936 8996
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8925 5319 8959
rect 5368 8956 5396 8996
rect 5534 8984 5540 9036
rect 5592 9024 5598 9036
rect 5629 9027 5687 9033
rect 5629 9024 5641 9027
rect 5592 8996 5641 9024
rect 5592 8984 5598 8996
rect 5629 8993 5641 8996
rect 5675 8993 5687 9027
rect 5629 8987 5687 8993
rect 6086 8984 6092 9036
rect 6144 9024 6150 9036
rect 6273 9027 6331 9033
rect 6273 9024 6285 9027
rect 6144 8996 6285 9024
rect 6144 8984 6150 8996
rect 6273 8993 6285 8996
rect 6319 8993 6331 9027
rect 6273 8987 6331 8993
rect 6380 8956 6408 9064
rect 7193 9061 7205 9064
rect 7239 9061 7251 9095
rect 7193 9055 7251 9061
rect 7377 9095 7435 9101
rect 7377 9061 7389 9095
rect 7423 9092 7435 9095
rect 7558 9092 7564 9104
rect 7423 9064 7564 9092
rect 7423 9061 7435 9064
rect 7377 9055 7435 9061
rect 7558 9052 7564 9064
rect 7616 9052 7622 9104
rect 9766 9052 9772 9104
rect 9824 9092 9830 9104
rect 9824 9064 10456 9092
rect 9824 9052 9830 9064
rect 7098 9024 7104 9036
rect 7059 8996 7104 9024
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 9858 9024 9864 9036
rect 9819 8996 9864 9024
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 5368 8928 6408 8956
rect 10137 8959 10195 8965
rect 5261 8919 5319 8925
rect 10137 8925 10149 8959
rect 10183 8956 10195 8959
rect 10226 8956 10232 8968
rect 10183 8928 10232 8956
rect 10183 8925 10195 8928
rect 10137 8919 10195 8925
rect 3752 8860 4936 8888
rect 5276 8888 5304 8919
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 10428 8956 10456 9064
rect 10962 9052 10968 9104
rect 11020 9092 11026 9104
rect 11020 9064 11100 9092
rect 11020 9052 11026 9064
rect 11072 9033 11100 9064
rect 11057 9027 11115 9033
rect 11057 8993 11069 9027
rect 11103 8993 11115 9027
rect 11057 8987 11115 8993
rect 12069 9027 12127 9033
rect 12069 8993 12081 9027
rect 12115 9024 12127 9027
rect 12894 9024 12900 9036
rect 12115 8996 12900 9024
rect 12115 8993 12127 8996
rect 12069 8987 12127 8993
rect 12894 8984 12900 8996
rect 12952 8984 12958 9036
rect 13173 9027 13231 9033
rect 13173 8993 13185 9027
rect 13219 9024 13231 9027
rect 16114 9024 16120 9036
rect 13219 8996 15424 9024
rect 16075 8996 16120 9024
rect 13219 8993 13231 8996
rect 13173 8987 13231 8993
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 10428 8928 10977 8956
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 13262 8956 13268 8968
rect 13223 8928 13268 8956
rect 10965 8919 11023 8925
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 15102 8916 15108 8968
rect 15160 8956 15166 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 15160 8928 15301 8956
rect 15160 8916 15166 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 15396 8956 15424 8996
rect 16114 8984 16120 8996
rect 16172 8984 16178 9036
rect 20901 9027 20959 9033
rect 20901 8993 20913 9027
rect 20947 9024 20959 9027
rect 21358 9024 21364 9036
rect 20947 8996 21364 9024
rect 20947 8993 20959 8996
rect 20901 8987 20959 8993
rect 21358 8984 21364 8996
rect 21416 8984 21422 9036
rect 20622 8956 20628 8968
rect 15396 8928 20628 8956
rect 15289 8919 15347 8925
rect 20622 8916 20628 8928
rect 20680 8916 20686 8968
rect 6089 8891 6147 8897
rect 6089 8888 6101 8891
rect 5276 8860 6101 8888
rect 3752 8848 3758 8860
rect 6089 8857 6101 8860
rect 6135 8857 6147 8891
rect 6089 8851 6147 8857
rect 9582 8848 9588 8900
rect 9640 8888 9646 8900
rect 12710 8888 12716 8900
rect 9640 8860 10916 8888
rect 12671 8860 12716 8888
rect 9640 8848 9646 8860
rect 5074 8820 5080 8832
rect 2746 8792 5080 8820
rect 1581 8783 1639 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 5258 8820 5264 8832
rect 5219 8792 5264 8820
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 7650 8820 7656 8832
rect 7611 8792 7656 8820
rect 7650 8780 7656 8792
rect 7708 8780 7714 8832
rect 9490 8820 9496 8832
rect 9451 8792 9496 8820
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 10686 8820 10692 8832
rect 10647 8792 10692 8820
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 10888 8829 10916 8860
rect 12710 8848 12716 8860
rect 12768 8848 12774 8900
rect 15657 8891 15715 8897
rect 15657 8857 15669 8891
rect 15703 8888 15715 8891
rect 16209 8891 16267 8897
rect 16209 8888 16221 8891
rect 15703 8860 16221 8888
rect 15703 8857 15715 8860
rect 15657 8851 15715 8857
rect 16209 8857 16221 8860
rect 16255 8857 16267 8891
rect 16209 8851 16267 8857
rect 10873 8823 10931 8829
rect 10873 8789 10885 8823
rect 10919 8789 10931 8823
rect 11882 8820 11888 8832
rect 11843 8792 11888 8820
rect 10873 8783 10931 8789
rect 11882 8780 11888 8792
rect 11940 8780 11946 8832
rect 20714 8820 20720 8832
rect 20675 8792 20720 8820
rect 20714 8780 20720 8792
rect 20772 8780 20778 8832
rect 1104 8730 21804 8752
rect 1104 8678 4432 8730
rect 4484 8678 4496 8730
rect 4548 8678 4560 8730
rect 4612 8678 4624 8730
rect 4676 8678 11332 8730
rect 11384 8678 11396 8730
rect 11448 8678 11460 8730
rect 11512 8678 11524 8730
rect 11576 8678 18232 8730
rect 18284 8678 18296 8730
rect 18348 8678 18360 8730
rect 18412 8678 18424 8730
rect 18476 8678 21804 8730
rect 1104 8656 21804 8678
rect 1670 8616 1676 8628
rect 1631 8588 1676 8616
rect 1670 8576 1676 8588
rect 1728 8576 1734 8628
rect 4890 8616 4896 8628
rect 4851 8588 4896 8616
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 5442 8616 5448 8628
rect 5132 8588 5448 8616
rect 5132 8576 5138 8588
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 9493 8619 9551 8625
rect 9493 8585 9505 8619
rect 9539 8616 9551 8619
rect 9582 8616 9588 8628
rect 9539 8588 9588 8616
rect 9539 8585 9551 8588
rect 9493 8579 9551 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 9858 8616 9864 8628
rect 9819 8588 9864 8616
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 13096 8588 16574 8616
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8480 9459 8483
rect 9766 8480 9772 8492
rect 9447 8452 9772 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 13096 8489 13124 8588
rect 14921 8551 14979 8557
rect 14921 8517 14933 8551
rect 14967 8517 14979 8551
rect 14921 8511 14979 8517
rect 15749 8551 15807 8557
rect 15749 8517 15761 8551
rect 15795 8548 15807 8551
rect 16209 8551 16267 8557
rect 16209 8548 16221 8551
rect 15795 8520 16221 8548
rect 15795 8517 15807 8520
rect 15749 8511 15807 8517
rect 16209 8517 16221 8520
rect 16255 8517 16267 8551
rect 16209 8511 16267 8517
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8449 13139 8483
rect 13262 8480 13268 8492
rect 13223 8452 13268 8480
rect 13081 8443 13139 8449
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 14936 8480 14964 8511
rect 16114 8480 16120 8492
rect 14936 8452 16120 8480
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 16546 8480 16574 8588
rect 20622 8576 20628 8628
rect 20680 8616 20686 8628
rect 20717 8619 20775 8625
rect 20717 8616 20729 8619
rect 20680 8588 20729 8616
rect 20680 8576 20686 8588
rect 20717 8585 20729 8588
rect 20763 8585 20775 8619
rect 20717 8579 20775 8585
rect 20714 8480 20720 8492
rect 16546 8452 20720 8480
rect 20714 8440 20720 8452
rect 20772 8440 20778 8492
rect 1486 8412 1492 8424
rect 1447 8384 1492 8412
rect 1486 8372 1492 8384
rect 1544 8372 1550 8424
rect 2038 8372 2044 8424
rect 2096 8412 2102 8424
rect 2133 8415 2191 8421
rect 2133 8412 2145 8415
rect 2096 8384 2145 8412
rect 2096 8372 2102 8384
rect 2133 8381 2145 8384
rect 2179 8381 2191 8415
rect 2682 8412 2688 8424
rect 2643 8384 2688 8412
rect 2133 8375 2191 8381
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 3386 8415 3444 8421
rect 3386 8381 3398 8415
rect 3432 8412 3444 8415
rect 4062 8412 4068 8424
rect 3432 8384 4068 8412
rect 3432 8381 3444 8384
rect 3386 8375 3444 8381
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 4985 8415 5043 8421
rect 4985 8381 4997 8415
rect 5031 8412 5043 8415
rect 5258 8412 5264 8424
rect 5031 8384 5264 8412
rect 5031 8381 5043 8384
rect 4985 8375 5043 8381
rect 5258 8372 5264 8384
rect 5316 8372 5322 8424
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 10870 8412 10876 8424
rect 9723 8384 10876 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 12894 8372 12900 8424
rect 12952 8412 12958 8424
rect 13280 8412 13308 8440
rect 12952 8384 13308 8412
rect 14553 8415 14611 8421
rect 12952 8372 12958 8384
rect 14553 8381 14565 8415
rect 14599 8412 14611 8415
rect 15381 8415 15439 8421
rect 15381 8412 15393 8415
rect 14599 8384 15393 8412
rect 14599 8381 14611 8384
rect 14553 8375 14611 8381
rect 15381 8381 15393 8384
rect 15427 8412 15439 8415
rect 15470 8412 15476 8424
rect 15427 8384 15476 8412
rect 15427 8381 15439 8384
rect 15381 8375 15439 8381
rect 15470 8372 15476 8384
rect 15528 8372 15534 8424
rect 16393 8415 16451 8421
rect 16393 8412 16405 8415
rect 15672 8384 16405 8412
rect 2593 8347 2651 8353
rect 2593 8313 2605 8347
rect 2639 8344 2651 8347
rect 2866 8344 2872 8356
rect 2639 8316 2872 8344
rect 2639 8313 2651 8316
rect 2593 8307 2651 8313
rect 2866 8304 2872 8316
rect 2924 8304 2930 8356
rect 14921 8347 14979 8353
rect 14921 8313 14933 8347
rect 14967 8344 14979 8347
rect 15102 8344 15108 8356
rect 14967 8316 15108 8344
rect 14967 8313 14979 8316
rect 14921 8307 14979 8313
rect 15102 8304 15108 8316
rect 15160 8344 15166 8356
rect 15672 8344 15700 8384
rect 16393 8381 16405 8384
rect 16439 8381 16451 8415
rect 20898 8412 20904 8424
rect 20859 8384 20904 8412
rect 16393 8375 16451 8381
rect 20898 8372 20904 8384
rect 20956 8372 20962 8424
rect 16114 8344 16120 8356
rect 15160 8316 15700 8344
rect 15764 8316 16120 8344
rect 15160 8304 15166 8316
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 3283 8279 3341 8285
rect 3283 8276 3295 8279
rect 3016 8248 3295 8276
rect 3016 8236 3022 8248
rect 3283 8245 3295 8248
rect 3329 8245 3341 8279
rect 10962 8276 10968 8288
rect 10923 8248 10968 8276
rect 3283 8239 3341 8245
rect 10962 8236 10968 8248
rect 11020 8236 11026 8288
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 12618 8276 12624 8288
rect 11112 8248 11157 8276
rect 12579 8248 12624 8276
rect 11112 8236 11118 8248
rect 12618 8236 12624 8248
rect 12676 8236 12682 8288
rect 12986 8276 12992 8288
rect 12947 8248 12992 8276
rect 12986 8236 12992 8248
rect 13044 8236 13050 8288
rect 15764 8285 15792 8316
rect 16114 8304 16120 8316
rect 16172 8304 16178 8356
rect 15749 8279 15807 8285
rect 15749 8245 15761 8279
rect 15795 8245 15807 8279
rect 15749 8239 15807 8245
rect 1104 8186 21804 8208
rect 1104 8134 7882 8186
rect 7934 8134 7946 8186
rect 7998 8134 8010 8186
rect 8062 8134 8074 8186
rect 8126 8134 14782 8186
rect 14834 8134 14846 8186
rect 14898 8134 14910 8186
rect 14962 8134 14974 8186
rect 15026 8134 21804 8186
rect 1104 8112 21804 8134
rect 6086 8072 6092 8084
rect 6047 8044 6092 8072
rect 6086 8032 6092 8044
rect 6144 8032 6150 8084
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 9861 8075 9919 8081
rect 9861 8072 9873 8075
rect 9732 8044 9873 8072
rect 9732 8032 9738 8044
rect 9861 8041 9873 8044
rect 9907 8041 9919 8075
rect 9861 8035 9919 8041
rect 10870 8032 10876 8084
rect 10928 8072 10934 8084
rect 12986 8072 12992 8084
rect 10928 8044 12434 8072
rect 12947 8044 12992 8072
rect 10928 8032 10934 8044
rect 11146 8004 11152 8016
rect 6288 7976 11152 8004
rect 6288 7945 6316 7976
rect 11146 7964 11152 7976
rect 11204 8004 11210 8016
rect 11241 8007 11299 8013
rect 11241 8004 11253 8007
rect 11204 7976 11253 8004
rect 11204 7964 11210 7976
rect 11241 7973 11253 7976
rect 11287 7973 11299 8007
rect 11241 7967 11299 7973
rect 6273 7939 6331 7945
rect 6273 7905 6285 7939
rect 6319 7905 6331 7939
rect 6273 7899 6331 7905
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7653 7939 7711 7945
rect 7653 7936 7665 7939
rect 7156 7908 7665 7936
rect 7156 7896 7162 7908
rect 7653 7905 7665 7908
rect 7699 7905 7711 7939
rect 7653 7899 7711 7905
rect 8205 7939 8263 7945
rect 8205 7905 8217 7939
rect 8251 7936 8263 7939
rect 10226 7936 10232 7948
rect 8251 7908 10232 7936
rect 8251 7905 8263 7908
rect 8205 7899 8263 7905
rect 9600 7877 9628 7908
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7936 10839 7939
rect 10870 7936 10876 7948
rect 10827 7908 10876 7936
rect 10827 7905 10839 7908
rect 10781 7899 10839 7905
rect 10870 7896 10876 7908
rect 10928 7896 10934 7948
rect 11333 7939 11391 7945
rect 11333 7905 11345 7939
rect 11379 7936 11391 7939
rect 11882 7936 11888 7948
rect 11379 7908 11888 7936
rect 11379 7905 11391 7908
rect 11333 7899 11391 7905
rect 11882 7896 11888 7908
rect 11940 7936 11946 7948
rect 11977 7939 12035 7945
rect 11977 7936 11989 7939
rect 11940 7908 11989 7936
rect 11940 7896 11946 7908
rect 11977 7905 11989 7908
rect 12023 7905 12035 7939
rect 12406 7936 12434 8044
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 15013 8075 15071 8081
rect 15013 8041 15025 8075
rect 15059 8072 15071 8075
rect 15102 8072 15108 8084
rect 15059 8044 15108 8072
rect 15059 8041 15071 8044
rect 15013 8035 15071 8041
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 15470 8072 15476 8084
rect 15431 8044 15476 8072
rect 15470 8032 15476 8044
rect 15528 8032 15534 8084
rect 15838 8072 15844 8084
rect 15799 8044 15844 8072
rect 15838 8032 15844 8044
rect 15896 8032 15902 8084
rect 20898 8072 20904 8084
rect 20859 8044 20904 8072
rect 20898 8032 20904 8044
rect 20956 8032 20962 8084
rect 12805 7939 12863 7945
rect 12805 7936 12817 7939
rect 12406 7908 12817 7936
rect 11977 7899 12035 7905
rect 12805 7905 12817 7908
rect 12851 7905 12863 7939
rect 12805 7899 12863 7905
rect 13722 7896 13728 7948
rect 13780 7936 13786 7948
rect 14829 7939 14887 7945
rect 14829 7936 14841 7939
rect 13780 7908 14841 7936
rect 13780 7896 13786 7908
rect 14829 7905 14841 7908
rect 14875 7905 14887 7939
rect 14829 7899 14887 7905
rect 15933 7939 15991 7945
rect 15933 7905 15945 7939
rect 15979 7936 15991 7939
rect 17954 7936 17960 7948
rect 15979 7908 17960 7936
rect 15979 7905 15991 7908
rect 15933 7899 15991 7905
rect 17954 7896 17960 7908
rect 18012 7896 18018 7948
rect 21082 7936 21088 7948
rect 21043 7908 21088 7936
rect 21082 7896 21088 7908
rect 21140 7896 21146 7948
rect 9585 7871 9643 7877
rect 9585 7837 9597 7871
rect 9631 7837 9643 7871
rect 9766 7868 9772 7880
rect 9727 7840 9772 7868
rect 9585 7831 9643 7837
rect 9766 7828 9772 7840
rect 9824 7828 9830 7880
rect 12894 7828 12900 7880
rect 12952 7868 12958 7880
rect 16025 7871 16083 7877
rect 16025 7868 16037 7871
rect 12952 7840 16037 7868
rect 12952 7828 12958 7840
rect 16025 7837 16037 7840
rect 16071 7837 16083 7871
rect 16025 7831 16083 7837
rect 10229 7735 10287 7741
rect 10229 7701 10241 7735
rect 10275 7732 10287 7735
rect 10318 7732 10324 7744
rect 10275 7704 10324 7732
rect 10275 7701 10287 7704
rect 10229 7695 10287 7701
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 11790 7732 11796 7744
rect 11751 7704 11796 7732
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 1104 7642 21804 7664
rect 1104 7590 4432 7642
rect 4484 7590 4496 7642
rect 4548 7590 4560 7642
rect 4612 7590 4624 7642
rect 4676 7590 11332 7642
rect 11384 7590 11396 7642
rect 11448 7590 11460 7642
rect 11512 7590 11524 7642
rect 11576 7590 18232 7642
rect 18284 7590 18296 7642
rect 18348 7590 18360 7642
rect 18412 7590 18424 7642
rect 18476 7590 21804 7642
rect 1104 7568 21804 7590
rect 11790 7528 11796 7540
rect 10244 7500 11796 7528
rect 10244 7469 10272 7500
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 13081 7531 13139 7537
rect 13081 7497 13093 7531
rect 13127 7528 13139 7531
rect 13722 7528 13728 7540
rect 13127 7500 13728 7528
rect 13127 7497 13139 7500
rect 13081 7491 13139 7497
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 10229 7463 10287 7469
rect 10229 7429 10241 7463
rect 10275 7429 10287 7463
rect 11054 7460 11060 7472
rect 11015 7432 11060 7460
rect 10229 7423 10287 7429
rect 11054 7420 11060 7432
rect 11112 7420 11118 7472
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 10318 7392 10324 7404
rect 9907 7364 10324 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 10318 7352 10324 7364
rect 10376 7392 10382 7404
rect 10376 7364 11008 7392
rect 10376 7352 10382 7364
rect 2958 7324 2964 7336
rect 2919 7296 2964 7324
rect 2958 7284 2964 7296
rect 3016 7284 3022 7336
rect 4706 7284 4712 7336
rect 4764 7324 4770 7336
rect 5169 7327 5227 7333
rect 5169 7324 5181 7327
rect 4764 7296 5181 7324
rect 4764 7284 4770 7296
rect 5169 7293 5181 7296
rect 5215 7324 5227 7327
rect 5442 7324 5448 7336
rect 5215 7296 5448 7324
rect 5215 7293 5227 7296
rect 5169 7287 5227 7293
rect 5442 7284 5448 7296
rect 5500 7284 5506 7336
rect 5718 7324 5724 7336
rect 5679 7296 5724 7324
rect 5718 7284 5724 7296
rect 5776 7284 5782 7336
rect 10689 7327 10747 7333
rect 10689 7293 10701 7327
rect 10735 7324 10747 7327
rect 10870 7324 10876 7336
rect 10735 7296 10876 7324
rect 10735 7293 10747 7296
rect 10689 7287 10747 7293
rect 10870 7284 10876 7296
rect 10928 7284 10934 7336
rect 10980 7324 11008 7364
rect 11882 7352 11888 7404
rect 11940 7392 11946 7404
rect 12069 7395 12127 7401
rect 12069 7392 12081 7395
rect 11940 7364 12081 7392
rect 11940 7352 11946 7364
rect 12069 7361 12081 7364
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 13265 7395 13323 7401
rect 13265 7361 13277 7395
rect 13311 7392 13323 7395
rect 14090 7392 14096 7404
rect 13311 7364 14096 7392
rect 13311 7361 13323 7364
rect 13265 7355 13323 7361
rect 14090 7352 14096 7364
rect 14148 7352 14154 7404
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 10980 7296 12449 7324
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 13722 7324 13728 7336
rect 13683 7296 13728 7324
rect 12437 7287 12495 7293
rect 13722 7284 13728 7296
rect 13780 7284 13786 7336
rect 17681 7327 17739 7333
rect 17681 7293 17693 7327
rect 17727 7324 17739 7327
rect 17770 7324 17776 7336
rect 17727 7296 17776 7324
rect 17727 7293 17739 7296
rect 17681 7287 17739 7293
rect 17770 7284 17776 7296
rect 17828 7284 17834 7336
rect 10962 7256 10968 7268
rect 10244 7228 10968 7256
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 2869 7191 2927 7197
rect 2869 7188 2881 7191
rect 2832 7160 2881 7188
rect 2832 7148 2838 7160
rect 2869 7157 2881 7160
rect 2915 7157 2927 7191
rect 4798 7188 4804 7200
rect 4759 7160 4804 7188
rect 2869 7151 2927 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 10244 7197 10272 7228
rect 10962 7216 10968 7228
rect 11020 7256 11026 7268
rect 12897 7259 12955 7265
rect 11020 7228 12112 7256
rect 11020 7216 11026 7228
rect 10229 7191 10287 7197
rect 10229 7157 10241 7191
rect 10275 7157 10287 7191
rect 10229 7151 10287 7157
rect 11057 7191 11115 7197
rect 11057 7157 11069 7191
rect 11103 7188 11115 7191
rect 11146 7188 11152 7200
rect 11103 7160 11152 7188
rect 11103 7157 11115 7160
rect 11057 7151 11115 7157
rect 11146 7148 11152 7160
rect 11204 7148 11210 7200
rect 12084 7197 12112 7228
rect 12897 7225 12909 7259
rect 12943 7256 12955 7259
rect 12986 7256 12992 7268
rect 12943 7228 12992 7256
rect 12943 7225 12955 7228
rect 12897 7219 12955 7225
rect 12986 7216 12992 7228
rect 13044 7216 13050 7268
rect 17494 7256 17500 7268
rect 17455 7228 17500 7256
rect 17494 7216 17500 7228
rect 17552 7216 17558 7268
rect 12069 7191 12127 7197
rect 12069 7157 12081 7191
rect 12115 7157 12127 7191
rect 12069 7151 12127 7157
rect 1104 7098 21804 7120
rect 1104 7046 7882 7098
rect 7934 7046 7946 7098
rect 7998 7046 8010 7098
rect 8062 7046 8074 7098
rect 8126 7046 14782 7098
rect 14834 7046 14846 7098
rect 14898 7046 14910 7098
rect 14962 7046 14974 7098
rect 15026 7046 21804 7098
rect 1104 7024 21804 7046
rect 4985 6987 5043 6993
rect 4985 6953 4997 6987
rect 5031 6984 5043 6987
rect 7190 6984 7196 6996
rect 5031 6956 7196 6984
rect 5031 6953 5043 6956
rect 4985 6947 5043 6953
rect 7190 6944 7196 6956
rect 7248 6944 7254 6996
rect 10870 6984 10876 6996
rect 10831 6956 10876 6984
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 11241 6987 11299 6993
rect 11241 6953 11253 6987
rect 11287 6984 11299 6987
rect 11698 6984 11704 6996
rect 11287 6956 11704 6984
rect 11287 6953 11299 6956
rect 11241 6947 11299 6953
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 13170 6984 13176 6996
rect 13131 6956 13176 6984
rect 13170 6944 13176 6956
rect 13228 6944 13234 6996
rect 12894 6916 12900 6928
rect 11256 6888 12900 6916
rect 1949 6851 2007 6857
rect 1949 6817 1961 6851
rect 1995 6848 2007 6851
rect 2498 6848 2504 6860
rect 1995 6820 2504 6848
rect 1995 6817 2007 6820
rect 1949 6811 2007 6817
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 2590 6808 2596 6860
rect 2648 6848 2654 6860
rect 6825 6851 6883 6857
rect 2648 6820 2693 6848
rect 2648 6808 2654 6820
rect 6825 6817 6837 6851
rect 6871 6848 6883 6851
rect 6914 6848 6920 6860
rect 6871 6820 6920 6848
rect 6871 6817 6883 6820
rect 6825 6811 6883 6817
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 4706 6780 4712 6792
rect 4667 6752 4712 6780
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 4890 6780 4896 6792
rect 4851 6752 4896 6780
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 11256 6780 11284 6888
rect 12894 6876 12900 6888
rect 12952 6876 12958 6928
rect 12986 6876 12992 6928
rect 13044 6916 13050 6928
rect 13044 6888 13860 6916
rect 13044 6876 13050 6888
rect 13832 6857 13860 6888
rect 11333 6851 11391 6857
rect 11333 6817 11345 6851
rect 11379 6848 11391 6851
rect 13817 6851 13875 6857
rect 11379 6820 13768 6848
rect 11379 6817 11391 6820
rect 11333 6811 11391 6817
rect 11425 6783 11483 6789
rect 11425 6780 11437 6783
rect 10284 6752 11437 6780
rect 10284 6740 10290 6752
rect 11425 6749 11437 6752
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 12805 6783 12863 6789
rect 12805 6749 12817 6783
rect 12851 6749 12863 6783
rect 13740 6780 13768 6820
rect 13817 6817 13829 6851
rect 13863 6848 13875 6851
rect 13863 6820 13897 6848
rect 13863 6817 13875 6820
rect 13817 6811 13875 6817
rect 19702 6808 19708 6860
rect 19760 6848 19766 6860
rect 20717 6851 20775 6857
rect 20717 6848 20729 6851
rect 19760 6820 20729 6848
rect 19760 6808 19766 6820
rect 20717 6817 20729 6820
rect 20763 6817 20775 6851
rect 20717 6811 20775 6817
rect 20622 6780 20628 6792
rect 13740 6752 20628 6780
rect 12805 6743 12863 6749
rect 1762 6712 1768 6724
rect 1723 6684 1768 6712
rect 1762 6672 1768 6684
rect 1820 6672 1826 6724
rect 2406 6712 2412 6724
rect 2367 6684 2412 6712
rect 2406 6672 2412 6684
rect 2464 6672 2470 6724
rect 5353 6715 5411 6721
rect 5353 6681 5365 6715
rect 5399 6712 5411 6715
rect 12710 6712 12716 6724
rect 5399 6684 12716 6712
rect 5399 6681 5411 6684
rect 5353 6675 5411 6681
rect 12710 6672 12716 6684
rect 12768 6712 12774 6724
rect 12820 6712 12848 6743
rect 20622 6740 20628 6752
rect 20680 6740 20686 6792
rect 12768 6684 12848 6712
rect 13173 6715 13231 6721
rect 12768 6672 12774 6684
rect 13173 6681 13185 6715
rect 13219 6712 13231 6715
rect 13633 6715 13691 6721
rect 13633 6712 13645 6715
rect 13219 6684 13645 6712
rect 13219 6681 13231 6684
rect 13173 6675 13231 6681
rect 13633 6681 13645 6684
rect 13679 6681 13691 6715
rect 13633 6675 13691 6681
rect 20901 6715 20959 6721
rect 20901 6681 20913 6715
rect 20947 6712 20959 6715
rect 21174 6712 21180 6724
rect 20947 6684 21180 6712
rect 20947 6681 20959 6684
rect 20901 6675 20959 6681
rect 21174 6672 21180 6684
rect 21232 6672 21238 6724
rect 6825 6647 6883 6653
rect 6825 6613 6837 6647
rect 6871 6644 6883 6647
rect 11974 6644 11980 6656
rect 6871 6616 11980 6644
rect 6871 6613 6883 6616
rect 6825 6607 6883 6613
rect 11974 6604 11980 6616
rect 12032 6644 12038 6656
rect 12250 6644 12256 6656
rect 12032 6616 12256 6644
rect 12032 6604 12038 6616
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 1104 6554 21804 6576
rect 1104 6502 4432 6554
rect 4484 6502 4496 6554
rect 4548 6502 4560 6554
rect 4612 6502 4624 6554
rect 4676 6502 11332 6554
rect 11384 6502 11396 6554
rect 11448 6502 11460 6554
rect 11512 6502 11524 6554
rect 11576 6502 18232 6554
rect 18284 6502 18296 6554
rect 18348 6502 18360 6554
rect 18412 6502 18424 6554
rect 18476 6502 21804 6554
rect 1104 6480 21804 6502
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 13170 6440 13176 6452
rect 2556 6412 12434 6440
rect 13131 6412 13176 6440
rect 2556 6400 2562 6412
rect 9585 6375 9643 6381
rect 9585 6372 9597 6375
rect 8220 6344 9597 6372
rect 2409 6307 2467 6313
rect 2409 6273 2421 6307
rect 2455 6304 2467 6307
rect 2774 6304 2780 6316
rect 2455 6276 2780 6304
rect 2455 6273 2467 6276
rect 2409 6267 2467 6273
rect 2774 6264 2780 6276
rect 2832 6264 2838 6316
rect 8220 6313 8248 6344
rect 9585 6341 9597 6344
rect 9631 6341 9643 6375
rect 12406 6372 12434 6412
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 13722 6440 13728 6452
rect 13683 6412 13728 6440
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 19702 6440 19708 6452
rect 19663 6412 19708 6440
rect 19702 6400 19708 6412
rect 19760 6400 19766 6452
rect 20622 6400 20628 6452
rect 20680 6440 20686 6452
rect 20717 6443 20775 6449
rect 20717 6440 20729 6443
rect 20680 6412 20729 6440
rect 20680 6400 20686 6412
rect 20717 6409 20729 6412
rect 20763 6409 20775 6443
rect 20717 6403 20775 6409
rect 14277 6375 14335 6381
rect 14277 6372 14289 6375
rect 12406 6344 14289 6372
rect 9585 6335 9643 6341
rect 14277 6341 14289 6344
rect 14323 6341 14335 6375
rect 14277 6335 14335 6341
rect 8205 6307 8263 6313
rect 8205 6304 8217 6307
rect 7668 6276 8217 6304
rect 4430 6236 4436 6248
rect 4391 6208 4436 6236
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 7668 6245 7696 6276
rect 8205 6273 8217 6276
rect 8251 6273 8263 6307
rect 10226 6304 10232 6316
rect 10187 6276 10232 6304
rect 8205 6267 8263 6273
rect 10226 6264 10232 6276
rect 10284 6264 10290 6316
rect 12710 6264 12716 6316
rect 12768 6304 12774 6316
rect 12805 6307 12863 6313
rect 12805 6304 12817 6307
rect 12768 6276 12817 6304
rect 12768 6264 12774 6276
rect 12805 6273 12817 6276
rect 12851 6273 12863 6307
rect 14737 6307 14795 6313
rect 14737 6304 14749 6307
rect 12805 6267 12863 6273
rect 12912 6276 14749 6304
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6205 7711 6239
rect 7653 6199 7711 6205
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6236 9183 6239
rect 10410 6236 10416 6248
rect 9171 6208 10416 6236
rect 9171 6205 9183 6208
rect 9125 6199 9183 6205
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 12161 6239 12219 6245
rect 12161 6205 12173 6239
rect 12207 6205 12219 6239
rect 12161 6199 12219 6205
rect 2590 6128 2596 6180
rect 2648 6168 2654 6180
rect 2685 6171 2743 6177
rect 2685 6168 2697 6171
rect 2648 6140 2697 6168
rect 2648 6128 2654 6140
rect 2685 6137 2697 6140
rect 2731 6137 2743 6171
rect 4062 6168 4068 6180
rect 3910 6140 4068 6168
rect 2685 6131 2743 6137
rect 2700 6100 2728 6131
rect 4062 6128 4068 6140
rect 4120 6128 4126 6180
rect 5718 6128 5724 6180
rect 5776 6168 5782 6180
rect 7469 6171 7527 6177
rect 7469 6168 7481 6171
rect 5776 6140 7481 6168
rect 5776 6128 5782 6140
rect 7469 6137 7481 6140
rect 7515 6137 7527 6171
rect 7469 6131 7527 6137
rect 8202 6128 8208 6180
rect 8260 6168 8266 6180
rect 8849 6171 8907 6177
rect 8849 6168 8861 6171
rect 8260 6140 8861 6168
rect 8260 6128 8266 6140
rect 8849 6137 8861 6140
rect 8895 6168 8907 6171
rect 12176 6168 12204 6199
rect 12250 6196 12256 6248
rect 12308 6236 12314 6248
rect 12912 6236 12940 6276
rect 14737 6273 14749 6276
rect 14783 6273 14795 6307
rect 14737 6267 14795 6273
rect 14921 6307 14979 6313
rect 14921 6273 14933 6307
rect 14967 6304 14979 6307
rect 15473 6307 15531 6313
rect 15473 6304 15485 6307
rect 14967 6276 15485 6304
rect 14967 6273 14979 6276
rect 14921 6267 14979 6273
rect 15473 6273 15485 6276
rect 15519 6273 15531 6307
rect 15473 6267 15531 6273
rect 15657 6307 15715 6313
rect 15657 6273 15669 6307
rect 15703 6304 15715 6307
rect 16206 6304 16212 6316
rect 15703 6276 16212 6304
rect 15703 6273 15715 6276
rect 15657 6267 15715 6273
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 17957 6307 18015 6313
rect 17957 6273 17969 6307
rect 18003 6304 18015 6307
rect 18046 6304 18052 6316
rect 18003 6276 18052 6304
rect 18003 6273 18015 6276
rect 17957 6267 18015 6273
rect 18046 6264 18052 6276
rect 18104 6304 18110 6316
rect 19702 6304 19708 6316
rect 18104 6276 19708 6304
rect 18104 6264 18110 6276
rect 19702 6264 19708 6276
rect 19760 6264 19766 6316
rect 12308 6208 12940 6236
rect 12308 6196 12314 6208
rect 13262 6196 13268 6248
rect 13320 6236 13326 6248
rect 13633 6239 13691 6245
rect 13633 6236 13645 6239
rect 13320 6208 13645 6236
rect 13320 6196 13326 6208
rect 13633 6205 13645 6208
rect 13679 6205 13691 6239
rect 13633 6199 13691 6205
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6205 15899 6239
rect 16114 6236 16120 6248
rect 16075 6208 16120 6236
rect 15841 6199 15899 6205
rect 12986 6168 12992 6180
rect 8895 6140 12204 6168
rect 12360 6140 12992 6168
rect 8895 6137 8907 6140
rect 8849 6131 8907 6137
rect 4430 6100 4436 6112
rect 2700 6072 4436 6100
rect 4430 6060 4436 6072
rect 4488 6060 4494 6112
rect 7282 6100 7288 6112
rect 7243 6072 7288 6100
rect 7282 6060 7288 6072
rect 7340 6060 7346 6112
rect 8662 6060 8668 6112
rect 8720 6100 8726 6112
rect 9953 6103 10011 6109
rect 9953 6100 9965 6103
rect 8720 6072 9965 6100
rect 8720 6060 8726 6072
rect 9953 6069 9965 6072
rect 9999 6069 10011 6103
rect 9953 6063 10011 6069
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 12360 6109 12388 6140
rect 12986 6128 12992 6140
rect 13044 6168 13050 6180
rect 13173 6171 13231 6177
rect 13173 6168 13185 6171
rect 13044 6140 13185 6168
rect 13044 6128 13050 6140
rect 13173 6137 13185 6140
rect 13219 6137 13231 6171
rect 15856 6168 15884 6199
rect 16114 6196 16120 6208
rect 16172 6196 16178 6248
rect 16482 6196 16488 6248
rect 16540 6236 16546 6248
rect 17681 6239 17739 6245
rect 17681 6236 17693 6239
rect 16540 6208 17693 6236
rect 16540 6196 16546 6208
rect 17681 6205 17693 6208
rect 17727 6205 17739 6239
rect 17681 6199 17739 6205
rect 20901 6239 20959 6245
rect 20901 6205 20913 6239
rect 20947 6236 20959 6239
rect 20990 6236 20996 6248
rect 20947 6208 20996 6236
rect 20947 6205 20959 6208
rect 20901 6199 20959 6205
rect 20990 6196 20996 6208
rect 21048 6196 21054 6248
rect 16574 6168 16580 6180
rect 15856 6140 16580 6168
rect 13173 6131 13231 6137
rect 16574 6128 16580 6140
rect 16632 6168 16638 6180
rect 17494 6168 17500 6180
rect 16632 6140 17500 6168
rect 16632 6128 16638 6140
rect 17494 6128 17500 6140
rect 17552 6128 17558 6180
rect 18598 6128 18604 6180
rect 18656 6128 18662 6180
rect 12345 6103 12403 6109
rect 10100 6072 10145 6100
rect 10100 6060 10106 6072
rect 12345 6069 12357 6103
rect 12391 6069 12403 6103
rect 14642 6100 14648 6112
rect 14603 6072 14648 6100
rect 12345 6063 12403 6069
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 1104 6010 21804 6032
rect 1104 5958 7882 6010
rect 7934 5958 7946 6010
rect 7998 5958 8010 6010
rect 8062 5958 8074 6010
rect 8126 5958 14782 6010
rect 14834 5958 14846 6010
rect 14898 5958 14910 6010
rect 14962 5958 14974 6010
rect 15026 5958 21804 6010
rect 1104 5936 21804 5958
rect 9674 5856 9680 5908
rect 9732 5896 9738 5908
rect 9861 5899 9919 5905
rect 9861 5896 9873 5899
rect 9732 5868 9873 5896
rect 9732 5856 9738 5868
rect 9861 5865 9873 5868
rect 9907 5865 9919 5899
rect 10410 5896 10416 5908
rect 10371 5868 10416 5896
rect 9861 5859 9919 5865
rect 6549 5831 6607 5837
rect 6549 5797 6561 5831
rect 6595 5828 6607 5831
rect 7098 5828 7104 5840
rect 6595 5800 7104 5828
rect 6595 5797 6607 5800
rect 6549 5791 6607 5797
rect 7098 5788 7104 5800
rect 7156 5828 7162 5840
rect 8202 5828 8208 5840
rect 7156 5800 8208 5828
rect 7156 5788 7162 5800
rect 8202 5788 8208 5800
rect 8260 5828 8266 5840
rect 8297 5831 8355 5837
rect 8297 5828 8309 5831
rect 8260 5800 8309 5828
rect 8260 5788 8266 5800
rect 8297 5797 8309 5800
rect 8343 5797 8355 5831
rect 8297 5791 8355 5797
rect 1578 5760 1584 5772
rect 1539 5732 1584 5760
rect 1578 5720 1584 5732
rect 1636 5720 1642 5772
rect 5718 5720 5724 5772
rect 5776 5760 5782 5772
rect 5905 5763 5963 5769
rect 5905 5760 5917 5763
rect 5776 5732 5917 5760
rect 5776 5720 5782 5732
rect 5905 5729 5917 5732
rect 5951 5729 5963 5763
rect 6638 5760 6644 5772
rect 6599 5732 6644 5760
rect 5905 5723 5963 5729
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 7282 5720 7288 5772
rect 7340 5760 7346 5772
rect 7653 5763 7711 5769
rect 7653 5760 7665 5763
rect 7340 5732 7665 5760
rect 7340 5720 7346 5732
rect 7653 5729 7665 5732
rect 7699 5729 7711 5763
rect 7653 5723 7711 5729
rect 8573 5763 8631 5769
rect 8573 5729 8585 5763
rect 8619 5760 8631 5763
rect 8662 5760 8668 5772
rect 8619 5732 8668 5760
rect 8619 5729 8631 5732
rect 8573 5723 8631 5729
rect 8662 5720 8668 5732
rect 8720 5720 8726 5772
rect 9490 5760 9496 5772
rect 9451 5732 9496 5760
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 9876 5760 9904 5859
rect 10410 5856 10416 5868
rect 10468 5856 10474 5908
rect 14642 5856 14648 5908
rect 14700 5896 14706 5908
rect 14829 5899 14887 5905
rect 14829 5896 14841 5899
rect 14700 5868 14841 5896
rect 14700 5856 14706 5868
rect 14829 5865 14841 5868
rect 14875 5865 14887 5899
rect 14829 5859 14887 5865
rect 15197 5899 15255 5905
rect 15197 5865 15209 5899
rect 15243 5896 15255 5899
rect 16117 5899 16175 5905
rect 16117 5896 16129 5899
rect 15243 5868 16129 5896
rect 15243 5865 15255 5868
rect 15197 5859 15255 5865
rect 16117 5865 16129 5868
rect 16163 5865 16175 5899
rect 16117 5859 16175 5865
rect 16485 5899 16543 5905
rect 16485 5865 16497 5899
rect 16531 5896 16543 5899
rect 17313 5899 17371 5905
rect 17313 5896 17325 5899
rect 16531 5868 17325 5896
rect 16531 5865 16543 5868
rect 16485 5859 16543 5865
rect 17313 5865 17325 5868
rect 17359 5865 17371 5899
rect 17313 5859 17371 5865
rect 17773 5899 17831 5905
rect 17773 5865 17785 5899
rect 17819 5896 17831 5899
rect 18046 5896 18052 5908
rect 17819 5868 18052 5896
rect 17819 5865 17831 5868
rect 17773 5859 17831 5865
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 20717 5899 20775 5905
rect 20717 5865 20729 5899
rect 20763 5865 20775 5899
rect 20717 5859 20775 5865
rect 10042 5788 10048 5840
rect 10100 5828 10106 5840
rect 20732 5828 20760 5859
rect 10100 5800 20760 5828
rect 10100 5788 10106 5800
rect 10321 5763 10379 5769
rect 10321 5760 10333 5763
rect 9876 5732 10333 5760
rect 10321 5729 10333 5732
rect 10367 5729 10379 5763
rect 10321 5723 10379 5729
rect 11885 5763 11943 5769
rect 11885 5729 11897 5763
rect 11931 5760 11943 5763
rect 12618 5760 12624 5772
rect 11931 5732 12624 5760
rect 11931 5729 11943 5732
rect 11885 5723 11943 5729
rect 12618 5720 12624 5732
rect 12676 5720 12682 5772
rect 17681 5763 17739 5769
rect 17681 5729 17693 5763
rect 17727 5760 17739 5763
rect 18046 5760 18052 5772
rect 17727 5732 18052 5760
rect 17727 5729 17739 5732
rect 17681 5723 17739 5729
rect 18046 5720 18052 5732
rect 18104 5720 18110 5772
rect 20898 5760 20904 5772
rect 20859 5732 20904 5760
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 4430 5652 4436 5704
rect 4488 5692 4494 5704
rect 12253 5695 12311 5701
rect 4488 5664 9996 5692
rect 4488 5652 4494 5664
rect 9858 5624 9864 5636
rect 9819 5596 9864 5624
rect 9858 5584 9864 5596
rect 9916 5584 9922 5636
rect 9968 5624 9996 5664
rect 12253 5661 12265 5695
rect 12299 5692 12311 5695
rect 12526 5692 12532 5704
rect 12299 5664 12532 5692
rect 12299 5661 12311 5664
rect 12253 5655 12311 5661
rect 12526 5652 12532 5664
rect 12584 5652 12590 5704
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 15473 5695 15531 5701
rect 15473 5661 15485 5695
rect 15519 5692 15531 5695
rect 15654 5692 15660 5704
rect 15519 5664 15660 5692
rect 15519 5661 15531 5664
rect 15473 5655 15531 5661
rect 15304 5624 15332 5655
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 15746 5652 15752 5704
rect 15804 5692 15810 5704
rect 16482 5692 16488 5704
rect 15804 5664 16488 5692
rect 15804 5652 15810 5664
rect 16482 5652 16488 5664
rect 16540 5692 16546 5704
rect 16577 5695 16635 5701
rect 16577 5692 16589 5695
rect 16540 5664 16589 5692
rect 16540 5652 16546 5664
rect 16577 5661 16589 5664
rect 16623 5661 16635 5695
rect 16577 5655 16635 5661
rect 16669 5695 16727 5701
rect 16669 5661 16681 5695
rect 16715 5661 16727 5695
rect 17862 5692 17868 5704
rect 17823 5664 17868 5692
rect 16669 5655 16727 5661
rect 9968 5596 15332 5624
rect 16390 5584 16396 5636
rect 16448 5624 16454 5636
rect 16684 5624 16712 5655
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 16448 5596 16712 5624
rect 16448 5584 16454 5596
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 12250 5556 12256 5568
rect 12211 5528 12256 5556
rect 12250 5516 12256 5528
rect 12308 5516 12314 5568
rect 1104 5466 21804 5488
rect 1104 5414 4432 5466
rect 4484 5414 4496 5466
rect 4548 5414 4560 5466
rect 4612 5414 4624 5466
rect 4676 5414 11332 5466
rect 11384 5414 11396 5466
rect 11448 5414 11460 5466
rect 11512 5414 11524 5466
rect 11576 5414 18232 5466
rect 18284 5414 18296 5466
rect 18348 5414 18360 5466
rect 18412 5414 18424 5466
rect 18476 5414 21804 5466
rect 1104 5392 21804 5414
rect 1578 5312 1584 5364
rect 1636 5352 1642 5364
rect 1765 5355 1823 5361
rect 1765 5352 1777 5355
rect 1636 5324 1777 5352
rect 1636 5312 1642 5324
rect 1765 5321 1777 5324
rect 1811 5321 1823 5355
rect 1765 5315 1823 5321
rect 5629 5355 5687 5361
rect 5629 5321 5641 5355
rect 5675 5352 5687 5355
rect 5718 5352 5724 5364
rect 5675 5324 5724 5352
rect 5675 5321 5687 5324
rect 5629 5315 5687 5321
rect 5718 5312 5724 5324
rect 5776 5312 5782 5364
rect 6914 5352 6920 5364
rect 6875 5324 6920 5352
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 8941 5355 8999 5361
rect 8941 5321 8953 5355
rect 8987 5352 8999 5355
rect 9674 5352 9680 5364
rect 8987 5324 9680 5352
rect 8987 5321 8999 5324
rect 8941 5315 8999 5321
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 9769 5355 9827 5361
rect 9769 5321 9781 5355
rect 9815 5352 9827 5355
rect 9858 5352 9864 5364
rect 9815 5324 9864 5352
rect 9815 5321 9827 5324
rect 9769 5315 9827 5321
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 15746 5352 15752 5364
rect 9968 5324 15752 5352
rect 9968 5284 9996 5324
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 18046 5312 18052 5364
rect 18104 5352 18110 5364
rect 18141 5355 18199 5361
rect 18141 5352 18153 5355
rect 18104 5324 18153 5352
rect 18104 5312 18110 5324
rect 18141 5321 18153 5324
rect 18187 5321 18199 5355
rect 18141 5315 18199 5321
rect 4540 5256 9996 5284
rect 12437 5287 12495 5293
rect 2777 5219 2835 5225
rect 2777 5216 2789 5219
rect 1964 5188 2789 5216
rect 1964 5157 1992 5188
rect 2777 5185 2789 5188
rect 2823 5216 2835 5219
rect 4540 5216 4568 5256
rect 12437 5253 12449 5287
rect 12483 5284 12495 5287
rect 12897 5287 12955 5293
rect 12897 5284 12909 5287
rect 12483 5256 12909 5284
rect 12483 5253 12495 5256
rect 12437 5247 12495 5253
rect 12897 5253 12909 5256
rect 12943 5253 12955 5287
rect 12897 5247 12955 5253
rect 2823 5188 4568 5216
rect 2823 5185 2835 5188
rect 2777 5179 2835 5185
rect 1949 5151 2007 5157
rect 1949 5117 1961 5151
rect 1995 5117 2007 5151
rect 2498 5148 2504 5160
rect 2459 5120 2504 5148
rect 1949 5111 2007 5117
rect 2498 5108 2504 5120
rect 2556 5108 2562 5160
rect 4540 5157 4568 5188
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5216 9183 5219
rect 9490 5216 9496 5228
rect 9171 5188 9496 5216
rect 9171 5185 9183 5188
rect 9125 5179 9183 5185
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 12069 5219 12127 5225
rect 12069 5185 12081 5219
rect 12115 5216 12127 5219
rect 12618 5216 12624 5228
rect 12115 5188 12624 5216
rect 12115 5185 12127 5188
rect 12069 5179 12127 5185
rect 12618 5176 12624 5188
rect 12676 5176 12682 5228
rect 15654 5216 15660 5228
rect 15615 5188 15660 5216
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 18156 5216 18184 5315
rect 19702 5312 19708 5364
rect 19760 5352 19766 5364
rect 20898 5352 20904 5364
rect 19760 5324 20208 5352
rect 20859 5324 20904 5352
rect 19760 5312 19766 5324
rect 19242 5216 19248 5228
rect 18156 5188 19248 5216
rect 19242 5176 19248 5188
rect 19300 5216 19306 5228
rect 20180 5225 20208 5324
rect 20898 5312 20904 5324
rect 20956 5312 20962 5364
rect 19889 5219 19947 5225
rect 19889 5216 19901 5219
rect 19300 5188 19901 5216
rect 19300 5176 19306 5188
rect 19889 5185 19901 5188
rect 19935 5185 19947 5219
rect 19889 5179 19947 5185
rect 20165 5219 20223 5225
rect 20165 5185 20177 5219
rect 20211 5185 20223 5219
rect 20165 5179 20223 5185
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5117 4583 5151
rect 4525 5111 4583 5117
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5117 5779 5151
rect 7098 5148 7104 5160
rect 7059 5120 7104 5148
rect 5721 5111 5779 5117
rect 4062 5080 4068 5092
rect 4002 5052 4068 5080
rect 4062 5040 4068 5052
rect 4120 5040 4126 5092
rect 5736 5080 5764 5111
rect 7098 5108 7104 5120
rect 7156 5108 7162 5160
rect 9585 5151 9643 5157
rect 9585 5148 9597 5151
rect 8772 5120 9597 5148
rect 4264 5052 5764 5080
rect 5905 5083 5963 5089
rect 2682 4972 2688 5024
rect 2740 5012 2746 5024
rect 4264 5012 4292 5052
rect 5905 5049 5917 5083
rect 5951 5080 5963 5083
rect 5994 5080 6000 5092
rect 5951 5052 6000 5080
rect 5951 5049 5963 5052
rect 5905 5043 5963 5049
rect 5994 5040 6000 5052
rect 6052 5040 6058 5092
rect 8662 5040 8668 5092
rect 8720 5080 8726 5092
rect 8772 5089 8800 5120
rect 9585 5117 9597 5120
rect 9631 5117 9643 5151
rect 9585 5111 9643 5117
rect 12526 5108 12532 5160
rect 12584 5148 12590 5160
rect 13081 5151 13139 5157
rect 13081 5148 13093 5151
rect 12584 5120 13093 5148
rect 12584 5108 12590 5120
rect 13081 5117 13093 5120
rect 13127 5117 13139 5151
rect 15838 5148 15844 5160
rect 15799 5120 15844 5148
rect 13081 5111 13139 5117
rect 15838 5108 15844 5120
rect 15896 5108 15902 5160
rect 16025 5151 16083 5157
rect 16025 5117 16037 5151
rect 16071 5117 16083 5151
rect 16025 5111 16083 5117
rect 8757 5083 8815 5089
rect 8757 5080 8769 5083
rect 8720 5052 8769 5080
rect 8720 5040 8726 5052
rect 8757 5049 8769 5052
rect 8803 5049 8815 5083
rect 16040 5080 16068 5111
rect 16114 5108 16120 5160
rect 16172 5148 16178 5160
rect 16209 5151 16267 5157
rect 16209 5148 16221 5151
rect 16172 5120 16221 5148
rect 16172 5108 16178 5120
rect 16209 5117 16221 5120
rect 16255 5148 16267 5151
rect 16666 5148 16672 5160
rect 16255 5120 16672 5148
rect 16255 5117 16267 5120
rect 16209 5111 16267 5117
rect 16666 5108 16672 5120
rect 16724 5108 16730 5160
rect 17497 5151 17555 5157
rect 17497 5117 17509 5151
rect 17543 5117 17555 5151
rect 21082 5148 21088 5160
rect 21043 5120 21088 5148
rect 17497 5111 17555 5117
rect 16574 5080 16580 5092
rect 16040 5052 16580 5080
rect 8757 5043 8815 5049
rect 16574 5040 16580 5052
rect 16632 5080 16638 5092
rect 17512 5080 17540 5111
rect 21082 5108 21088 5120
rect 21140 5108 21146 5160
rect 16632 5052 17540 5080
rect 16632 5040 16638 5052
rect 18138 5040 18144 5092
rect 18196 5080 18202 5092
rect 18598 5080 18604 5092
rect 18196 5052 18604 5080
rect 18196 5040 18202 5052
rect 18598 5040 18604 5052
rect 18656 5080 18662 5092
rect 18656 5052 18722 5080
rect 18656 5040 18662 5052
rect 2740 4984 4292 5012
rect 2740 4972 2746 4984
rect 12250 4972 12256 5024
rect 12308 5012 12314 5024
rect 12437 5015 12495 5021
rect 12437 5012 12449 5015
rect 12308 4984 12449 5012
rect 12308 4972 12314 4984
rect 12437 4981 12449 4984
rect 12483 4981 12495 5015
rect 17402 5012 17408 5024
rect 17363 4984 17408 5012
rect 12437 4975 12495 4981
rect 17402 4972 17408 4984
rect 17460 4972 17466 5024
rect 1104 4922 21804 4944
rect 1104 4870 7882 4922
rect 7934 4870 7946 4922
rect 7998 4870 8010 4922
rect 8062 4870 8074 4922
rect 8126 4870 14782 4922
rect 14834 4870 14846 4922
rect 14898 4870 14910 4922
rect 14962 4870 14974 4922
rect 15026 4870 21804 4922
rect 1104 4848 21804 4870
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 5813 4811 5871 4817
rect 5813 4808 5825 4811
rect 4120 4780 5825 4808
rect 4120 4768 4126 4780
rect 5813 4777 5825 4780
rect 5859 4777 5871 4811
rect 6638 4808 6644 4820
rect 6599 4780 6644 4808
rect 5813 4771 5871 4777
rect 5828 4740 5856 4771
rect 6638 4768 6644 4780
rect 6696 4768 6702 4820
rect 10505 4811 10563 4817
rect 10505 4777 10517 4811
rect 10551 4808 10563 4811
rect 10686 4808 10692 4820
rect 10551 4780 10692 4808
rect 10551 4777 10563 4780
rect 10505 4771 10563 4777
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 11146 4768 11152 4820
rect 11204 4808 11210 4820
rect 11701 4811 11759 4817
rect 11701 4808 11713 4811
rect 11204 4780 11713 4808
rect 11204 4768 11210 4780
rect 11701 4777 11713 4780
rect 11747 4808 11759 4811
rect 12529 4811 12587 4817
rect 12529 4808 12541 4811
rect 11747 4780 12541 4808
rect 11747 4777 11759 4780
rect 11701 4771 11759 4777
rect 12529 4777 12541 4780
rect 12575 4777 12587 4811
rect 16390 4808 16396 4820
rect 16351 4780 16396 4808
rect 12529 4771 12587 4777
rect 16390 4768 16396 4780
rect 16448 4768 16454 4820
rect 17773 4743 17831 4749
rect 5828 4712 16344 4740
rect 5905 4675 5963 4681
rect 5905 4641 5917 4675
rect 5951 4672 5963 4675
rect 5994 4672 6000 4684
rect 5951 4644 6000 4672
rect 5951 4641 5963 4644
rect 5905 4635 5963 4641
rect 5994 4632 6000 4644
rect 6052 4632 6058 4684
rect 12526 4672 12532 4684
rect 12487 4644 12532 4672
rect 12526 4632 12532 4644
rect 12584 4632 12590 4684
rect 13262 4672 13268 4684
rect 13223 4644 13268 4672
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 10226 4604 10232 4616
rect 10139 4576 10232 4604
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 10410 4604 10416 4616
rect 10371 4576 10416 4604
rect 10410 4564 10416 4576
rect 10468 4564 10474 4616
rect 11333 4607 11391 4613
rect 11333 4573 11345 4607
rect 11379 4604 11391 4607
rect 12161 4607 12219 4613
rect 12161 4604 12173 4607
rect 11379 4576 12173 4604
rect 11379 4573 11391 4576
rect 11333 4567 11391 4573
rect 12161 4573 12173 4576
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 10244 4536 10272 4564
rect 10778 4536 10784 4548
rect 10244 4508 10784 4536
rect 10778 4496 10784 4508
rect 10836 4496 10842 4548
rect 10873 4539 10931 4545
rect 10873 4505 10885 4539
rect 10919 4536 10931 4539
rect 11348 4536 11376 4567
rect 11698 4536 11704 4548
rect 10919 4508 11376 4536
rect 11659 4508 11704 4536
rect 10919 4505 10931 4508
rect 10873 4499 10931 4505
rect 11698 4496 11704 4508
rect 11756 4496 11762 4548
rect 12544 4536 12572 4632
rect 16206 4604 16212 4616
rect 16167 4576 16212 4604
rect 16206 4564 16212 4576
rect 16264 4564 16270 4616
rect 16316 4604 16344 4712
rect 16408 4712 17448 4740
rect 16408 4681 16436 4712
rect 17420 4684 17448 4712
rect 17773 4709 17785 4743
rect 17819 4740 17831 4743
rect 17862 4740 17868 4752
rect 17819 4712 17868 4740
rect 17819 4709 17831 4712
rect 17773 4703 17831 4709
rect 17862 4700 17868 4712
rect 17920 4700 17926 4752
rect 16393 4675 16451 4681
rect 16393 4641 16405 4675
rect 16439 4641 16451 4675
rect 16666 4672 16672 4684
rect 16579 4644 16672 4672
rect 16393 4635 16451 4641
rect 16666 4632 16672 4644
rect 16724 4672 16730 4684
rect 17218 4672 17224 4684
rect 16724 4644 17224 4672
rect 16724 4632 16730 4644
rect 17218 4632 17224 4644
rect 17276 4632 17282 4684
rect 17402 4672 17408 4684
rect 17363 4644 17408 4672
rect 17402 4632 17408 4644
rect 17460 4632 17466 4684
rect 18138 4672 18144 4684
rect 17512 4644 18144 4672
rect 17512 4604 17540 4644
rect 18138 4632 18144 4644
rect 18196 4632 18202 4684
rect 16316 4576 17540 4604
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4573 17647 4607
rect 17589 4567 17647 4573
rect 13081 4539 13139 4545
rect 13081 4536 13093 4539
rect 12544 4508 13093 4536
rect 13081 4505 13093 4508
rect 13127 4505 13139 4539
rect 13081 4499 13139 4505
rect 15838 4496 15844 4548
rect 15896 4536 15902 4548
rect 17604 4536 17632 4567
rect 15896 4508 17632 4536
rect 15896 4496 15902 4508
rect 1104 4378 21804 4400
rect 1104 4326 4432 4378
rect 4484 4326 4496 4378
rect 4548 4326 4560 4378
rect 4612 4326 4624 4378
rect 4676 4326 11332 4378
rect 11384 4326 11396 4378
rect 11448 4326 11460 4378
rect 11512 4326 11524 4378
rect 11576 4326 18232 4378
rect 18284 4326 18296 4378
rect 18348 4326 18360 4378
rect 18412 4326 18424 4378
rect 18476 4326 21804 4378
rect 1104 4304 21804 4326
rect 11698 4224 11704 4276
rect 11756 4264 11762 4276
rect 12161 4267 12219 4273
rect 12161 4264 12173 4267
rect 11756 4236 12173 4264
rect 11756 4224 11762 4236
rect 12161 4233 12173 4236
rect 12207 4233 12219 4267
rect 13262 4264 13268 4276
rect 13223 4236 13268 4264
rect 12161 4227 12219 4233
rect 13262 4224 13268 4236
rect 13320 4224 13326 4276
rect 15838 4224 15844 4276
rect 15896 4264 15902 4276
rect 16301 4267 16359 4273
rect 16301 4264 16313 4267
rect 15896 4236 16313 4264
rect 15896 4224 15902 4236
rect 16301 4233 16313 4236
rect 16347 4233 16359 4267
rect 16301 4227 16359 4233
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4128 3571 4131
rect 13265 4131 13323 4137
rect 13265 4128 13277 4131
rect 3559 4100 13277 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 13265 4097 13277 4100
rect 13311 4128 13323 4131
rect 14090 4128 14096 4140
rect 13311 4100 14096 4128
rect 13311 4097 13323 4100
rect 13265 4091 13323 4097
rect 14090 4088 14096 4100
rect 14148 4088 14154 4140
rect 2041 4063 2099 4069
rect 2041 4029 2053 4063
rect 2087 4060 2099 4063
rect 2774 4060 2780 4072
rect 2087 4032 2780 4060
rect 2087 4029 2099 4032
rect 2041 4023 2099 4029
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 2866 4020 2872 4072
rect 2924 4060 2930 4072
rect 3329 4063 3387 4069
rect 3329 4060 3341 4063
rect 2924 4032 3341 4060
rect 2924 4020 2930 4032
rect 3329 4029 3341 4032
rect 3375 4029 3387 4063
rect 3329 4023 3387 4029
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 8021 4063 8079 4069
rect 8021 4060 8033 4063
rect 7708 4032 8033 4060
rect 7708 4020 7714 4032
rect 8021 4029 8033 4032
rect 8067 4029 8079 4063
rect 8021 4023 8079 4029
rect 10781 4063 10839 4069
rect 10781 4029 10793 4063
rect 10827 4060 10839 4063
rect 11146 4060 11152 4072
rect 10827 4032 11152 4060
rect 10827 4029 10839 4032
rect 10781 4023 10839 4029
rect 11146 4020 11152 4032
rect 11204 4020 11210 4072
rect 12250 4060 12256 4072
rect 12211 4032 12256 4060
rect 12250 4020 12256 4032
rect 12308 4020 12314 4072
rect 13630 4060 13636 4072
rect 13591 4032 13636 4060
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 15470 4020 15476 4072
rect 15528 4060 15534 4072
rect 16206 4060 16212 4072
rect 15528 4032 16212 4060
rect 15528 4020 15534 4032
rect 16206 4020 16212 4032
rect 16264 4020 16270 4072
rect 19242 4020 19248 4072
rect 19300 4060 19306 4072
rect 20257 4063 20315 4069
rect 20257 4060 20269 4063
rect 19300 4032 20269 4060
rect 19300 4020 19306 4032
rect 20257 4029 20269 4032
rect 20303 4029 20315 4063
rect 20257 4023 20315 4029
rect 8662 3992 8668 4004
rect 8623 3964 8668 3992
rect 8662 3952 8668 3964
rect 8720 3952 8726 4004
rect 8941 3995 8999 4001
rect 8941 3961 8953 3995
rect 8987 3961 8999 3995
rect 8941 3955 8999 3961
rect 1854 3924 1860 3936
rect 1815 3896 1860 3924
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 8956 3924 8984 3955
rect 13906 3952 13912 4004
rect 13964 3992 13970 4004
rect 14093 3995 14151 4001
rect 14093 3992 14105 3995
rect 13964 3964 14105 3992
rect 13964 3952 13970 3964
rect 14093 3961 14105 3964
rect 14139 3961 14151 3995
rect 14093 3955 14151 3961
rect 10502 3924 10508 3936
rect 8956 3896 10508 3924
rect 10502 3884 10508 3896
rect 10560 3924 10566 3936
rect 10689 3927 10747 3933
rect 10689 3924 10701 3927
rect 10560 3896 10701 3924
rect 10560 3884 10566 3896
rect 10689 3893 10701 3896
rect 10735 3893 10747 3927
rect 14182 3924 14188 3936
rect 14143 3896 14188 3924
rect 10689 3887 10747 3893
rect 14182 3884 14188 3896
rect 14240 3884 14246 3936
rect 20441 3927 20499 3933
rect 20441 3893 20453 3927
rect 20487 3924 20499 3927
rect 20898 3924 20904 3936
rect 20487 3896 20904 3924
rect 20487 3893 20499 3896
rect 20441 3887 20499 3893
rect 20898 3884 20904 3896
rect 20956 3884 20962 3936
rect 1104 3834 21804 3856
rect 1104 3782 7882 3834
rect 7934 3782 7946 3834
rect 7998 3782 8010 3834
rect 8062 3782 8074 3834
rect 8126 3782 14782 3834
rect 14834 3782 14846 3834
rect 14898 3782 14910 3834
rect 14962 3782 14974 3834
rect 15026 3782 21804 3834
rect 1104 3760 21804 3782
rect 13262 3680 13268 3732
rect 13320 3720 13326 3732
rect 13357 3723 13415 3729
rect 13357 3720 13369 3723
rect 13320 3692 13369 3720
rect 13320 3680 13326 3692
rect 13357 3689 13369 3692
rect 13403 3689 13415 3723
rect 15102 3720 15108 3732
rect 15063 3692 15108 3720
rect 13357 3683 13415 3689
rect 15102 3680 15108 3692
rect 15160 3680 15166 3732
rect 20901 3723 20959 3729
rect 20901 3689 20913 3723
rect 20947 3720 20959 3723
rect 20990 3720 20996 3732
rect 20947 3692 20996 3720
rect 20947 3689 20959 3692
rect 20901 3683 20959 3689
rect 20990 3680 20996 3692
rect 21048 3680 21054 3732
rect 5994 3652 6000 3664
rect 5955 3624 6000 3652
rect 5994 3612 6000 3624
rect 6052 3612 6058 3664
rect 8297 3655 8355 3661
rect 8297 3621 8309 3655
rect 8343 3652 8355 3655
rect 8662 3652 8668 3664
rect 8343 3624 8668 3652
rect 8343 3621 8355 3624
rect 8297 3615 8355 3621
rect 8662 3612 8668 3624
rect 8720 3612 8726 3664
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 6181 3587 6239 3593
rect 6181 3553 6193 3587
rect 6227 3584 6239 3587
rect 6914 3584 6920 3596
rect 6227 3556 6920 3584
rect 6227 3553 6239 3556
rect 6181 3547 6239 3553
rect 6914 3544 6920 3556
rect 6972 3544 6978 3596
rect 7650 3584 7656 3596
rect 7611 3556 7656 3584
rect 7650 3544 7656 3556
rect 7708 3544 7714 3596
rect 8570 3584 8576 3596
rect 8531 3556 8576 3584
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 9493 3587 9551 3593
rect 9493 3553 9505 3587
rect 9539 3584 9551 3587
rect 10502 3584 10508 3596
rect 9539 3556 10508 3584
rect 9539 3553 9551 3556
rect 9493 3547 9551 3553
rect 10502 3544 10508 3556
rect 10560 3544 10566 3596
rect 11425 3587 11483 3593
rect 11425 3553 11437 3587
rect 11471 3584 11483 3587
rect 11471 3556 12020 3584
rect 11471 3553 11483 3556
rect 11425 3547 11483 3553
rect 9858 3516 9864 3528
rect 9819 3488 9864 3516
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 11992 3457 12020 3556
rect 12066 3544 12072 3596
rect 12124 3584 12130 3596
rect 12161 3587 12219 3593
rect 12161 3584 12173 3587
rect 12124 3556 12173 3584
rect 12124 3544 12130 3556
rect 12161 3553 12173 3556
rect 12207 3553 12219 3587
rect 12161 3547 12219 3553
rect 13357 3587 13415 3593
rect 13357 3553 13369 3587
rect 13403 3584 13415 3587
rect 14182 3584 14188 3596
rect 13403 3556 14188 3584
rect 13403 3553 13415 3556
rect 13357 3547 13415 3553
rect 14182 3544 14188 3556
rect 14240 3544 14246 3596
rect 15197 3587 15255 3593
rect 15197 3553 15209 3587
rect 15243 3584 15255 3587
rect 20714 3584 20720 3596
rect 15243 3556 20720 3584
rect 15243 3553 15255 3556
rect 15197 3547 15255 3553
rect 20714 3544 20720 3556
rect 20772 3544 20778 3596
rect 21085 3587 21143 3593
rect 21085 3553 21097 3587
rect 21131 3584 21143 3587
rect 22094 3584 22100 3596
rect 21131 3556 22100 3584
rect 21131 3553 21143 3556
rect 21085 3547 21143 3553
rect 22094 3544 22100 3556
rect 22152 3544 22158 3596
rect 13630 3476 13636 3528
rect 13688 3516 13694 3528
rect 13725 3519 13783 3525
rect 13725 3516 13737 3519
rect 13688 3488 13737 3516
rect 13688 3476 13694 3488
rect 13725 3485 13737 3488
rect 13771 3485 13783 3519
rect 15378 3516 15384 3528
rect 15339 3488 15384 3516
rect 13725 3479 13783 3485
rect 11977 3451 12035 3457
rect 11977 3417 11989 3451
rect 12023 3417 12035 3451
rect 13740 3448 13768 3479
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 14737 3451 14795 3457
rect 14737 3448 14749 3451
rect 13740 3420 14749 3448
rect 11977 3411 12035 3417
rect 14737 3417 14749 3420
rect 14783 3417 14795 3451
rect 14737 3411 14795 3417
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3380 1639 3383
rect 2498 3380 2504 3392
rect 1627 3352 2504 3380
rect 1627 3349 1639 3352
rect 1581 3343 1639 3349
rect 2498 3340 2504 3352
rect 2556 3340 2562 3392
rect 9306 3340 9312 3392
rect 9364 3380 9370 3392
rect 9493 3383 9551 3389
rect 9493 3380 9505 3383
rect 9364 3352 9505 3380
rect 9364 3340 9370 3352
rect 9493 3349 9505 3352
rect 9539 3349 9551 3383
rect 9493 3343 9551 3349
rect 9582 3340 9588 3392
rect 9640 3380 9646 3392
rect 10321 3383 10379 3389
rect 10321 3380 10333 3383
rect 9640 3352 10333 3380
rect 9640 3340 9646 3352
rect 10321 3349 10333 3352
rect 10367 3349 10379 3383
rect 10321 3343 10379 3349
rect 10686 3340 10692 3392
rect 10744 3380 10750 3392
rect 11241 3383 11299 3389
rect 11241 3380 11253 3383
rect 10744 3352 11253 3380
rect 10744 3340 10750 3352
rect 11241 3349 11253 3352
rect 11287 3349 11299 3383
rect 11241 3343 11299 3349
rect 1104 3290 21804 3312
rect 1104 3238 4432 3290
rect 4484 3238 4496 3290
rect 4548 3238 4560 3290
rect 4612 3238 4624 3290
rect 4676 3238 11332 3290
rect 11384 3238 11396 3290
rect 11448 3238 11460 3290
rect 11512 3238 11524 3290
rect 11576 3238 18232 3290
rect 18284 3238 18296 3290
rect 18348 3238 18360 3290
rect 18412 3238 18424 3290
rect 18476 3238 21804 3290
rect 1104 3216 21804 3238
rect 1946 3136 1952 3188
rect 2004 3176 2010 3188
rect 2041 3179 2099 3185
rect 2041 3176 2053 3179
rect 2004 3148 2053 3176
rect 2004 3136 2010 3148
rect 2041 3145 2053 3148
rect 2087 3145 2099 3179
rect 2041 3139 2099 3145
rect 4617 3179 4675 3185
rect 4617 3145 4629 3179
rect 4663 3176 4675 3179
rect 4890 3176 4896 3188
rect 4663 3148 4896 3176
rect 4663 3145 4675 3148
rect 4617 3139 4675 3145
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 7006 3176 7012 3188
rect 6967 3148 7012 3176
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 8570 3136 8576 3188
rect 8628 3176 8634 3188
rect 8757 3179 8815 3185
rect 8757 3176 8769 3179
rect 8628 3148 8769 3176
rect 8628 3136 8634 3148
rect 8757 3145 8769 3148
rect 8803 3145 8815 3179
rect 9306 3176 9312 3188
rect 8757 3139 8815 3145
rect 8864 3148 9312 3176
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 2314 2972 2320 2984
rect 1903 2944 2320 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 2314 2932 2320 2944
rect 2372 2932 2378 2984
rect 2498 2972 2504 2984
rect 2459 2944 2504 2972
rect 2498 2932 2504 2944
rect 2556 2932 2562 2984
rect 4430 2972 4436 2984
rect 4391 2944 4436 2972
rect 4430 2932 4436 2944
rect 4488 2932 4494 2984
rect 6822 2972 6828 2984
rect 6783 2944 6828 2972
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 8864 2981 8892 3148
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 15378 3176 15384 3188
rect 12728 3148 15384 3176
rect 9858 3108 9864 3120
rect 9692 3080 9864 3108
rect 9309 3043 9367 3049
rect 9309 3009 9321 3043
rect 9355 3040 9367 3043
rect 9582 3040 9588 3052
rect 9355 3012 9588 3040
rect 9355 3009 9367 3012
rect 9309 3003 9367 3009
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 9692 3049 9720 3080
rect 9858 3068 9864 3080
rect 9916 3108 9922 3120
rect 10229 3111 10287 3117
rect 10229 3108 10241 3111
rect 9916 3080 10241 3108
rect 9916 3068 9922 3080
rect 10229 3077 10241 3080
rect 10275 3077 10287 3111
rect 10229 3071 10287 3077
rect 9677 3043 9735 3049
rect 9677 3009 9689 3043
rect 9723 3009 9735 3043
rect 10686 3040 10692 3052
rect 10647 3012 10692 3040
rect 9677 3003 9735 3009
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 10778 3000 10784 3052
rect 10836 3040 10842 3052
rect 12728 3049 12756 3148
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 17954 3136 17960 3188
rect 18012 3176 18018 3188
rect 18049 3179 18107 3185
rect 18049 3176 18061 3179
rect 18012 3148 18061 3176
rect 18012 3136 18018 3148
rect 18049 3145 18061 3148
rect 18095 3145 18107 3179
rect 20714 3176 20720 3188
rect 20675 3148 20720 3176
rect 18049 3139 18107 3145
rect 20714 3136 20720 3148
rect 20772 3136 20778 3188
rect 13906 3108 13912 3120
rect 13867 3080 13912 3108
rect 13906 3068 13912 3080
rect 13964 3068 13970 3120
rect 14553 3111 14611 3117
rect 14553 3077 14565 3111
rect 14599 3077 14611 3111
rect 14553 3071 14611 3077
rect 10873 3043 10931 3049
rect 10873 3040 10885 3043
rect 10836 3012 10885 3040
rect 10836 3000 10842 3012
rect 10873 3009 10885 3012
rect 10919 3040 10931 3043
rect 12713 3043 12771 3049
rect 12713 3040 12725 3043
rect 10919 3012 12725 3040
rect 10919 3009 10931 3012
rect 10873 3003 10931 3009
rect 12713 3009 12725 3012
rect 12759 3009 12771 3043
rect 12713 3003 12771 3009
rect 12805 3043 12863 3049
rect 12805 3009 12817 3043
rect 12851 3040 12863 3043
rect 14568 3040 14596 3071
rect 17218 3068 17224 3120
rect 17276 3108 17282 3120
rect 17313 3111 17371 3117
rect 17313 3108 17325 3111
rect 17276 3080 17325 3108
rect 17276 3068 17282 3080
rect 17313 3077 17325 3080
rect 17359 3077 17371 3111
rect 17313 3071 17371 3077
rect 20257 3111 20315 3117
rect 20257 3077 20269 3111
rect 20303 3077 20315 3111
rect 20257 3071 20315 3077
rect 15378 3040 15384 3052
rect 12851 3012 14596 3040
rect 15339 3012 15384 3040
rect 12851 3009 12863 3012
rect 12805 3003 12863 3009
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 8849 2975 8907 2981
rect 8849 2941 8861 2975
rect 8895 2941 8907 2975
rect 10594 2972 10600 2984
rect 10555 2944 10600 2972
rect 8849 2935 8907 2941
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 13725 2975 13783 2981
rect 13725 2972 13737 2975
rect 13280 2944 13737 2972
rect 9766 2904 9772 2916
rect 2700 2876 9772 2904
rect 2700 2845 2728 2876
rect 9766 2864 9772 2876
rect 9824 2864 9830 2916
rect 12802 2864 12808 2916
rect 12860 2904 12866 2916
rect 12897 2907 12955 2913
rect 12897 2904 12909 2907
rect 12860 2876 12909 2904
rect 12860 2864 12866 2876
rect 12897 2873 12909 2876
rect 12943 2873 12955 2907
rect 12897 2867 12955 2873
rect 13280 2848 13308 2944
rect 13725 2941 13737 2944
rect 13771 2941 13783 2975
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 13725 2935 13783 2941
rect 13832 2944 14749 2972
rect 13354 2864 13360 2916
rect 13412 2904 13418 2916
rect 13832 2904 13860 2944
rect 14737 2941 14749 2944
rect 14783 2941 14795 2975
rect 16114 2972 16120 2984
rect 16075 2944 16120 2972
rect 14737 2935 14795 2941
rect 16114 2932 16120 2944
rect 16172 2932 16178 2984
rect 18230 2972 18236 2984
rect 18191 2944 18236 2972
rect 18230 2932 18236 2944
rect 18288 2932 18294 2984
rect 20070 2972 20076 2984
rect 20031 2944 20076 2972
rect 20070 2932 20076 2944
rect 20128 2932 20134 2984
rect 20272 2972 20300 3071
rect 20901 2975 20959 2981
rect 20901 2972 20913 2975
rect 20272 2944 20913 2972
rect 20901 2941 20913 2944
rect 20947 2941 20959 2975
rect 20901 2935 20959 2941
rect 14090 2904 14096 2916
rect 13412 2876 13860 2904
rect 14051 2876 14096 2904
rect 13412 2864 13418 2876
rect 14090 2864 14096 2876
rect 14148 2864 14154 2916
rect 17494 2904 17500 2916
rect 17455 2876 17500 2904
rect 17494 2864 17500 2876
rect 17552 2864 17558 2916
rect 2685 2839 2743 2845
rect 2685 2805 2697 2839
rect 2731 2805 2743 2839
rect 13262 2836 13268 2848
rect 13223 2808 13268 2836
rect 2685 2799 2743 2805
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 1104 2746 21804 2768
rect 1104 2694 7882 2746
rect 7934 2694 7946 2746
rect 7998 2694 8010 2746
rect 8062 2694 8074 2746
rect 8126 2694 14782 2746
rect 14834 2694 14846 2746
rect 14898 2694 14910 2746
rect 14962 2694 14974 2746
rect 15026 2694 21804 2746
rect 1104 2672 21804 2694
rect 2314 2592 2320 2644
rect 2372 2632 2378 2644
rect 2593 2635 2651 2641
rect 2593 2632 2605 2635
rect 2372 2604 2605 2632
rect 2372 2592 2378 2604
rect 2593 2601 2605 2604
rect 2639 2601 2651 2635
rect 4430 2632 4436 2644
rect 4391 2604 4436 2632
rect 2593 2595 2651 2601
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 5721 2635 5779 2641
rect 5721 2601 5733 2635
rect 5767 2632 5779 2635
rect 6822 2632 6828 2644
rect 5767 2604 6828 2632
rect 5767 2601 5779 2604
rect 5721 2595 5779 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 6914 2592 6920 2644
rect 6972 2632 6978 2644
rect 9769 2635 9827 2641
rect 6972 2604 7017 2632
rect 6972 2592 6978 2604
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 10410 2632 10416 2644
rect 9815 2604 10416 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 10689 2635 10747 2641
rect 10689 2601 10701 2635
rect 10735 2601 10747 2635
rect 10689 2595 10747 2601
rect 13173 2635 13231 2641
rect 13173 2601 13185 2635
rect 13219 2632 13231 2635
rect 13906 2632 13912 2644
rect 13219 2604 13912 2632
rect 13219 2601 13231 2604
rect 13173 2595 13231 2601
rect 1854 2524 1860 2576
rect 1912 2564 1918 2576
rect 2041 2567 2099 2573
rect 2041 2564 2053 2567
rect 1912 2536 2053 2564
rect 1912 2524 1918 2536
rect 2041 2533 2053 2536
rect 2087 2533 2099 2567
rect 8754 2564 8760 2576
rect 2041 2527 2099 2533
rect 8496 2536 8760 2564
rect 474 2456 480 2508
rect 532 2496 538 2508
rect 2777 2499 2835 2505
rect 2777 2496 2789 2499
rect 532 2468 2789 2496
rect 532 2456 538 2468
rect 2777 2465 2789 2468
rect 2823 2465 2835 2499
rect 2777 2459 2835 2465
rect 3694 2456 3700 2508
rect 3752 2496 3758 2508
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 3752 2468 4261 2496
rect 3752 2456 3758 2468
rect 4249 2465 4261 2468
rect 4295 2465 4307 2499
rect 5534 2496 5540 2508
rect 5495 2468 5540 2496
rect 4249 2459 4307 2465
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 8496 2505 8524 2536
rect 8754 2524 8760 2536
rect 8812 2524 8818 2576
rect 10704 2564 10732 2595
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 16114 2632 16120 2644
rect 16075 2604 16120 2632
rect 16114 2592 16120 2604
rect 16172 2592 16178 2644
rect 17494 2592 17500 2644
rect 17552 2632 17558 2644
rect 17589 2635 17647 2641
rect 17589 2632 17601 2635
rect 17552 2604 17601 2632
rect 17552 2592 17558 2604
rect 17589 2601 17601 2604
rect 17635 2601 17647 2635
rect 17589 2595 17647 2601
rect 18230 2592 18236 2644
rect 18288 2632 18294 2644
rect 18877 2635 18935 2641
rect 18877 2632 18889 2635
rect 18288 2604 18889 2632
rect 18288 2592 18294 2604
rect 18877 2601 18889 2604
rect 18923 2601 18935 2635
rect 18877 2595 18935 2601
rect 15289 2567 15347 2573
rect 15289 2564 15301 2567
rect 10704 2536 15301 2564
rect 15289 2533 15301 2536
rect 15335 2533 15347 2567
rect 15470 2564 15476 2576
rect 15431 2536 15476 2564
rect 15289 2527 15347 2533
rect 15470 2524 15476 2536
rect 15528 2524 15534 2576
rect 20898 2564 20904 2576
rect 20859 2536 20904 2564
rect 20898 2524 20904 2536
rect 20956 2524 20962 2576
rect 7101 2499 7159 2505
rect 7101 2496 7113 2499
rect 6972 2468 7113 2496
rect 6972 2456 6978 2468
rect 7101 2465 7113 2468
rect 7147 2465 7159 2499
rect 7101 2459 7159 2465
rect 8481 2499 8539 2505
rect 8481 2465 8493 2499
rect 8527 2465 8539 2499
rect 9585 2499 9643 2505
rect 9585 2496 9597 2499
rect 8481 2459 8539 2465
rect 8680 2468 9597 2496
rect 1854 2360 1860 2372
rect 1815 2332 1860 2360
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 8680 2369 8708 2468
rect 9585 2465 9597 2468
rect 9631 2465 9643 2499
rect 9585 2459 9643 2465
rect 10505 2499 10563 2505
rect 10505 2465 10517 2499
rect 10551 2496 10563 2499
rect 10594 2496 10600 2508
rect 10551 2468 10600 2496
rect 10551 2465 10563 2468
rect 10505 2459 10563 2465
rect 10594 2456 10600 2468
rect 10652 2456 10658 2508
rect 11149 2499 11207 2505
rect 11149 2465 11161 2499
rect 11195 2465 11207 2499
rect 11149 2459 11207 2465
rect 12805 2499 12863 2505
rect 12805 2465 12817 2499
rect 12851 2496 12863 2499
rect 13262 2496 13268 2508
rect 12851 2468 13268 2496
rect 12851 2465 12863 2468
rect 12805 2459 12863 2465
rect 11164 2428 11192 2459
rect 13262 2456 13268 2468
rect 13320 2456 13326 2508
rect 13817 2499 13875 2505
rect 13817 2465 13829 2499
rect 13863 2496 13875 2499
rect 14090 2496 14096 2508
rect 13863 2468 14096 2496
rect 13863 2465 13875 2468
rect 13817 2459 13875 2465
rect 14090 2456 14096 2468
rect 14148 2456 14154 2508
rect 15654 2456 15660 2508
rect 15712 2496 15718 2508
rect 15933 2499 15991 2505
rect 15933 2496 15945 2499
rect 15712 2468 15945 2496
rect 15712 2456 15718 2468
rect 15933 2465 15945 2468
rect 15979 2465 15991 2499
rect 15933 2459 15991 2465
rect 17034 2456 17040 2508
rect 17092 2496 17098 2508
rect 17773 2499 17831 2505
rect 17773 2496 17785 2499
rect 17092 2468 17785 2496
rect 17092 2456 17098 2468
rect 17773 2465 17785 2468
rect 17819 2465 17831 2499
rect 17773 2459 17831 2465
rect 18874 2456 18880 2508
rect 18932 2496 18938 2508
rect 19061 2499 19119 2505
rect 19061 2496 19073 2499
rect 18932 2468 19073 2496
rect 18932 2456 18938 2468
rect 19061 2465 19073 2468
rect 19107 2465 19119 2499
rect 19061 2459 19119 2465
rect 13722 2428 13728 2440
rect 11164 2400 13728 2428
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 8665 2363 8723 2369
rect 8665 2329 8677 2363
rect 8711 2329 8723 2363
rect 8665 2323 8723 2329
rect 13173 2363 13231 2369
rect 13173 2329 13185 2363
rect 13219 2360 13231 2363
rect 13633 2363 13691 2369
rect 13633 2360 13645 2363
rect 13219 2332 13645 2360
rect 13219 2329 13231 2332
rect 13173 2323 13231 2329
rect 13633 2329 13645 2332
rect 13679 2329 13691 2363
rect 20714 2360 20720 2372
rect 20675 2332 20720 2360
rect 13633 2323 13691 2329
rect 20714 2320 20720 2332
rect 20772 2320 20778 2372
rect 11333 2295 11391 2301
rect 11333 2261 11345 2295
rect 11379 2292 11391 2295
rect 13354 2292 13360 2304
rect 11379 2264 13360 2292
rect 11379 2261 11391 2264
rect 11333 2255 11391 2261
rect 13354 2252 13360 2264
rect 13412 2252 13418 2304
rect 1104 2202 21804 2224
rect 1104 2150 4432 2202
rect 4484 2150 4496 2202
rect 4548 2150 4560 2202
rect 4612 2150 4624 2202
rect 4676 2150 11332 2202
rect 11384 2150 11396 2202
rect 11448 2150 11460 2202
rect 11512 2150 11524 2202
rect 11576 2150 18232 2202
rect 18284 2150 18296 2202
rect 18348 2150 18360 2202
rect 18412 2150 18424 2202
rect 18476 2150 21804 2202
rect 1104 2128 21804 2150
<< via1 >>
rect 4432 22822 4484 22874
rect 4496 22822 4548 22874
rect 4560 22822 4612 22874
rect 4624 22822 4676 22874
rect 11332 22822 11384 22874
rect 11396 22822 11448 22874
rect 11460 22822 11512 22874
rect 11524 22822 11576 22874
rect 18232 22822 18284 22874
rect 18296 22822 18348 22874
rect 18360 22822 18412 22874
rect 18424 22822 18476 22874
rect 1492 22763 1544 22772
rect 1492 22729 1501 22763
rect 1501 22729 1535 22763
rect 1535 22729 1544 22763
rect 1492 22720 1544 22729
rect 940 22516 992 22568
rect 2780 22559 2832 22568
rect 2780 22525 2789 22559
rect 2789 22525 2823 22559
rect 2823 22525 2832 22559
rect 2780 22516 2832 22525
rect 4804 22516 4856 22568
rect 6000 22559 6052 22568
rect 6000 22525 6009 22559
rect 6009 22525 6043 22559
rect 6043 22525 6052 22559
rect 6000 22516 6052 22525
rect 7840 22559 7892 22568
rect 7840 22525 7849 22559
rect 7849 22525 7883 22559
rect 7883 22525 7892 22559
rect 7840 22516 7892 22525
rect 9680 22516 9732 22568
rect 12900 22559 12952 22568
rect 1584 22491 1636 22500
rect 1584 22457 1593 22491
rect 1593 22457 1627 22491
rect 1627 22457 1636 22491
rect 1584 22448 1636 22457
rect 11704 22448 11756 22500
rect 12900 22525 12909 22559
rect 12909 22525 12943 22559
rect 12943 22525 12952 22559
rect 12900 22516 12952 22525
rect 14740 22516 14792 22568
rect 16580 22516 16632 22568
rect 17960 22516 18012 22568
rect 19800 22516 19852 22568
rect 21088 22559 21140 22568
rect 21088 22525 21097 22559
rect 21097 22525 21131 22559
rect 21131 22525 21140 22559
rect 21088 22516 21140 22525
rect 1676 22380 1728 22432
rect 3424 22380 3476 22432
rect 5080 22380 5132 22432
rect 5724 22380 5776 22432
rect 8208 22380 8260 22432
rect 9680 22423 9732 22432
rect 9680 22389 9689 22423
rect 9689 22389 9723 22423
rect 9723 22389 9732 22423
rect 9680 22380 9732 22389
rect 10324 22380 10376 22432
rect 13084 22423 13136 22432
rect 13084 22389 13093 22423
rect 13093 22389 13127 22423
rect 13127 22389 13136 22423
rect 13084 22380 13136 22389
rect 15384 22380 15436 22432
rect 16028 22380 16080 22432
rect 16672 22380 16724 22432
rect 20168 22380 20220 22432
rect 21364 22380 21416 22432
rect 7882 22278 7934 22330
rect 7946 22278 7998 22330
rect 8010 22278 8062 22330
rect 8074 22278 8126 22330
rect 14782 22278 14834 22330
rect 14846 22278 14898 22330
rect 14910 22278 14962 22330
rect 14974 22278 15026 22330
rect 6828 22108 6880 22160
rect 7012 22040 7064 22092
rect 5172 22015 5224 22024
rect 5172 21981 5181 22015
rect 5181 21981 5215 22015
rect 5215 21981 5224 22015
rect 5172 21972 5224 21981
rect 5816 21972 5868 22024
rect 9680 22040 9732 22092
rect 12072 22040 12124 22092
rect 13084 22083 13136 22092
rect 13084 22049 13093 22083
rect 13093 22049 13127 22083
rect 13127 22049 13136 22083
rect 13084 22040 13136 22049
rect 16672 22083 16724 22092
rect 9772 21972 9824 22024
rect 10692 22015 10744 22024
rect 10692 21981 10701 22015
rect 10701 21981 10735 22015
rect 10735 21981 10744 22015
rect 10692 21972 10744 21981
rect 11060 21972 11112 22024
rect 12256 21972 12308 22024
rect 16672 22049 16681 22083
rect 16681 22049 16715 22083
rect 16715 22049 16724 22083
rect 16672 22040 16724 22049
rect 20812 22040 20864 22092
rect 21640 22040 21692 22092
rect 17592 22015 17644 22024
rect 15200 21904 15252 21956
rect 17592 21981 17601 22015
rect 17601 21981 17635 22015
rect 17635 21981 17644 22015
rect 17592 21972 17644 21981
rect 17684 21972 17736 22024
rect 6460 21836 6512 21888
rect 8484 21836 8536 21888
rect 10232 21836 10284 21888
rect 10968 21836 11020 21888
rect 13360 21836 13412 21888
rect 14648 21836 14700 21888
rect 16856 21879 16908 21888
rect 16856 21845 16865 21879
rect 16865 21845 16899 21879
rect 16899 21845 16908 21879
rect 16856 21836 16908 21845
rect 19984 21836 20036 21888
rect 4432 21734 4484 21786
rect 4496 21734 4548 21786
rect 4560 21734 4612 21786
rect 4624 21734 4676 21786
rect 11332 21734 11384 21786
rect 11396 21734 11448 21786
rect 11460 21734 11512 21786
rect 11524 21734 11576 21786
rect 18232 21734 18284 21786
rect 18296 21734 18348 21786
rect 18360 21734 18412 21786
rect 18424 21734 18476 21786
rect 1584 21632 1636 21684
rect 6828 21675 6880 21684
rect 6828 21641 6837 21675
rect 6837 21641 6871 21675
rect 6871 21641 6880 21675
rect 6828 21632 6880 21641
rect 3240 21564 3292 21616
rect 5172 21564 5224 21616
rect 8392 21632 8444 21684
rect 11060 21675 11112 21684
rect 11060 21641 11069 21675
rect 11069 21641 11103 21675
rect 11103 21641 11112 21675
rect 11060 21632 11112 21641
rect 12072 21675 12124 21684
rect 12072 21641 12081 21675
rect 12081 21641 12115 21675
rect 12115 21641 12124 21675
rect 12072 21632 12124 21641
rect 17592 21632 17644 21684
rect 10692 21564 10744 21616
rect 3424 21471 3476 21480
rect 3424 21437 3433 21471
rect 3433 21437 3467 21471
rect 3467 21437 3476 21471
rect 3424 21428 3476 21437
rect 5080 21471 5132 21480
rect 5080 21437 5089 21471
rect 5089 21437 5123 21471
rect 5123 21437 5132 21471
rect 5080 21428 5132 21437
rect 5724 21471 5776 21480
rect 5724 21437 5733 21471
rect 5733 21437 5767 21471
rect 5767 21437 5776 21471
rect 5724 21428 5776 21437
rect 7012 21471 7064 21480
rect 7012 21437 7021 21471
rect 7021 21437 7055 21471
rect 7055 21437 7064 21471
rect 7012 21428 7064 21437
rect 11060 21496 11112 21548
rect 11152 21428 11204 21480
rect 12256 21471 12308 21480
rect 12256 21437 12265 21471
rect 12265 21437 12299 21471
rect 12299 21437 12308 21471
rect 12256 21428 12308 21437
rect 14280 21564 14332 21616
rect 19984 21564 20036 21616
rect 14004 21496 14056 21548
rect 15108 21496 15160 21548
rect 16856 21496 16908 21548
rect 15384 21471 15436 21480
rect 5356 21360 5408 21412
rect 8484 21360 8536 21412
rect 3700 21292 3752 21344
rect 5448 21292 5500 21344
rect 5908 21335 5960 21344
rect 5908 21301 5917 21335
rect 5917 21301 5951 21335
rect 5951 21301 5960 21335
rect 5908 21292 5960 21301
rect 10600 21292 10652 21344
rect 10968 21360 11020 21412
rect 10876 21292 10928 21344
rect 15384 21437 15393 21471
rect 15393 21437 15427 21471
rect 15427 21437 15436 21471
rect 15384 21428 15436 21437
rect 16028 21471 16080 21480
rect 16028 21437 16037 21471
rect 16037 21437 16071 21471
rect 16071 21437 16080 21471
rect 16028 21428 16080 21437
rect 19340 21428 19392 21480
rect 19984 21428 20036 21480
rect 14648 21360 14700 21412
rect 18144 21360 18196 21412
rect 21088 21428 21140 21480
rect 15200 21292 15252 21344
rect 15844 21335 15896 21344
rect 15844 21301 15853 21335
rect 15853 21301 15887 21335
rect 15887 21301 15896 21335
rect 15844 21292 15896 21301
rect 19892 21335 19944 21344
rect 19892 21301 19901 21335
rect 19901 21301 19935 21335
rect 19935 21301 19944 21335
rect 19892 21292 19944 21301
rect 7882 21190 7934 21242
rect 7946 21190 7998 21242
rect 8010 21190 8062 21242
rect 8074 21190 8126 21242
rect 14782 21190 14834 21242
rect 14846 21190 14898 21242
rect 14910 21190 14962 21242
rect 14974 21190 15026 21242
rect 5816 21131 5868 21140
rect 5816 21097 5825 21131
rect 5825 21097 5859 21131
rect 5859 21097 5868 21131
rect 5816 21088 5868 21097
rect 9772 21088 9824 21140
rect 10876 21088 10928 21140
rect 18144 21131 18196 21140
rect 5724 21020 5776 21072
rect 6460 21020 6512 21072
rect 10968 21020 11020 21072
rect 5816 20952 5868 21004
rect 8208 20995 8260 21004
rect 8208 20961 8217 20995
rect 8217 20961 8251 20995
rect 8251 20961 8260 20995
rect 8208 20952 8260 20961
rect 10600 20995 10652 21004
rect 10600 20961 10609 20995
rect 10609 20961 10643 20995
rect 10643 20961 10652 20995
rect 10600 20952 10652 20961
rect 10784 20995 10836 21004
rect 10784 20961 10793 20995
rect 10793 20961 10827 20995
rect 10827 20961 10836 20995
rect 10784 20952 10836 20961
rect 11060 20995 11112 21004
rect 11060 20961 11069 20995
rect 11069 20961 11103 20995
rect 11103 20961 11112 20995
rect 11060 20952 11112 20961
rect 15568 21020 15620 21072
rect 18144 21097 18153 21131
rect 18153 21097 18187 21131
rect 18187 21097 18196 21131
rect 18144 21088 18196 21097
rect 15200 20995 15252 21004
rect 15200 20961 15209 20995
rect 15209 20961 15243 20995
rect 15243 20961 15252 20995
rect 15200 20952 15252 20961
rect 17500 20952 17552 21004
rect 20168 20995 20220 21004
rect 20168 20961 20177 20995
rect 20177 20961 20211 20995
rect 20211 20961 20220 20995
rect 20168 20952 20220 20961
rect 21180 20952 21232 21004
rect 6552 20884 6604 20936
rect 12348 20884 12400 20936
rect 15476 20927 15528 20936
rect 15476 20893 15485 20927
rect 15485 20893 15519 20927
rect 15519 20893 15528 20927
rect 15476 20884 15528 20893
rect 6092 20816 6144 20868
rect 11796 20748 11848 20800
rect 16948 20791 17000 20800
rect 16948 20757 16957 20791
rect 16957 20757 16991 20791
rect 16991 20757 17000 20791
rect 16948 20748 17000 20757
rect 19616 20748 19668 20800
rect 20628 20748 20680 20800
rect 4432 20646 4484 20698
rect 4496 20646 4548 20698
rect 4560 20646 4612 20698
rect 4624 20646 4676 20698
rect 11332 20646 11384 20698
rect 11396 20646 11448 20698
rect 11460 20646 11512 20698
rect 11524 20646 11576 20698
rect 18232 20646 18284 20698
rect 18296 20646 18348 20698
rect 18360 20646 18412 20698
rect 18424 20646 18476 20698
rect 14004 20587 14056 20596
rect 14004 20553 14013 20587
rect 14013 20553 14047 20587
rect 14047 20553 14056 20587
rect 14004 20544 14056 20553
rect 21088 20587 21140 20596
rect 21088 20553 21097 20587
rect 21097 20553 21131 20587
rect 21131 20553 21140 20587
rect 21088 20544 21140 20553
rect 6920 20519 6972 20528
rect 6920 20485 6929 20519
rect 6929 20485 6963 20519
rect 6963 20485 6972 20519
rect 6920 20476 6972 20485
rect 3240 20451 3292 20460
rect 3240 20417 3249 20451
rect 3249 20417 3283 20451
rect 3283 20417 3292 20451
rect 3240 20408 3292 20417
rect 4068 20408 4120 20460
rect 1400 20383 1452 20392
rect 1400 20349 1409 20383
rect 1409 20349 1443 20383
rect 1443 20349 1452 20383
rect 1400 20340 1452 20349
rect 6092 20408 6144 20460
rect 8392 20451 8444 20460
rect 8392 20417 8401 20451
rect 8401 20417 8435 20451
rect 8435 20417 8444 20451
rect 8392 20408 8444 20417
rect 5632 20383 5684 20392
rect 5632 20349 5641 20383
rect 5641 20349 5675 20383
rect 5675 20349 5684 20383
rect 5632 20340 5684 20349
rect 7012 20383 7064 20392
rect 7012 20349 7021 20383
rect 7021 20349 7055 20383
rect 7055 20349 7064 20383
rect 7012 20340 7064 20349
rect 7104 20383 7156 20392
rect 7104 20349 7113 20383
rect 7113 20349 7147 20383
rect 7147 20349 7156 20383
rect 11060 20476 11112 20528
rect 10968 20408 11020 20460
rect 7104 20340 7156 20349
rect 11152 20383 11204 20392
rect 11152 20349 11161 20383
rect 11161 20349 11195 20383
rect 11195 20349 11204 20383
rect 11152 20340 11204 20349
rect 11244 20340 11296 20392
rect 14556 20476 14608 20528
rect 19984 20408 20036 20460
rect 3516 20315 3568 20324
rect 3516 20281 3525 20315
rect 3525 20281 3559 20315
rect 3559 20281 3568 20315
rect 3516 20272 3568 20281
rect 4252 20272 4304 20324
rect 9404 20272 9456 20324
rect 2412 20204 2464 20256
rect 5540 20247 5592 20256
rect 5540 20213 5549 20247
rect 5549 20213 5583 20247
rect 5583 20213 5592 20247
rect 5540 20204 5592 20213
rect 10784 20204 10836 20256
rect 14464 20272 14516 20324
rect 15108 20340 15160 20392
rect 19340 20383 19392 20392
rect 19340 20349 19349 20383
rect 19349 20349 19383 20383
rect 19383 20349 19392 20383
rect 19340 20340 19392 20349
rect 15752 20272 15804 20324
rect 20628 20272 20680 20324
rect 14648 20204 14700 20256
rect 7882 20102 7934 20154
rect 7946 20102 7998 20154
rect 8010 20102 8062 20154
rect 8074 20102 8126 20154
rect 14782 20102 14834 20154
rect 14846 20102 14898 20154
rect 14910 20102 14962 20154
rect 14974 20102 15026 20154
rect 3516 20000 3568 20052
rect 5816 20000 5868 20052
rect 9404 20000 9456 20052
rect 14464 20000 14516 20052
rect 20628 20043 20680 20052
rect 5540 19932 5592 19984
rect 6184 19975 6236 19984
rect 6184 19941 6193 19975
rect 6193 19941 6227 19975
rect 6227 19941 6236 19975
rect 20628 20009 20637 20043
rect 20637 20009 20671 20043
rect 20671 20009 20680 20043
rect 20628 20000 20680 20009
rect 6184 19932 6236 19941
rect 15200 19932 15252 19984
rect 6368 19907 6420 19916
rect 6368 19873 6377 19907
rect 6377 19873 6411 19907
rect 6411 19873 6420 19907
rect 6368 19864 6420 19873
rect 6644 19864 6696 19916
rect 7104 19864 7156 19916
rect 8024 19907 8076 19916
rect 5632 19796 5684 19848
rect 8024 19873 8033 19907
rect 8033 19873 8067 19907
rect 8067 19873 8076 19907
rect 8024 19864 8076 19873
rect 9772 19864 9824 19916
rect 12440 19864 12492 19916
rect 14924 19907 14976 19916
rect 14924 19873 14933 19907
rect 14933 19873 14967 19907
rect 14967 19873 14976 19907
rect 14924 19864 14976 19873
rect 15752 19907 15804 19916
rect 13176 19839 13228 19848
rect 13176 19805 13185 19839
rect 13185 19805 13219 19839
rect 13219 19805 13228 19839
rect 13176 19796 13228 19805
rect 6552 19728 6604 19780
rect 8024 19728 8076 19780
rect 13820 19796 13872 19848
rect 14188 19796 14240 19848
rect 14648 19796 14700 19848
rect 15752 19873 15761 19907
rect 15761 19873 15795 19907
rect 15795 19873 15804 19907
rect 15752 19864 15804 19873
rect 16028 19907 16080 19916
rect 16028 19873 16037 19907
rect 16037 19873 16071 19907
rect 16071 19873 16080 19907
rect 16028 19864 16080 19873
rect 20812 19907 20864 19916
rect 20812 19873 20821 19907
rect 20821 19873 20855 19907
rect 20855 19873 20864 19907
rect 20812 19864 20864 19873
rect 13728 19728 13780 19780
rect 15476 19728 15528 19780
rect 5540 19660 5592 19712
rect 5724 19660 5776 19712
rect 7012 19660 7064 19712
rect 7748 19660 7800 19712
rect 8208 19660 8260 19712
rect 11704 19660 11756 19712
rect 14096 19660 14148 19712
rect 4432 19558 4484 19610
rect 4496 19558 4548 19610
rect 4560 19558 4612 19610
rect 4624 19558 4676 19610
rect 11332 19558 11384 19610
rect 11396 19558 11448 19610
rect 11460 19558 11512 19610
rect 11524 19558 11576 19610
rect 18232 19558 18284 19610
rect 18296 19558 18348 19610
rect 18360 19558 18412 19610
rect 18424 19558 18476 19610
rect 4252 19456 4304 19508
rect 6092 19456 6144 19508
rect 7104 19456 7156 19508
rect 14372 19456 14424 19508
rect 15200 19456 15252 19508
rect 16304 19456 16356 19508
rect 16120 19388 16172 19440
rect 12624 19363 12676 19372
rect 12624 19329 12633 19363
rect 12633 19329 12667 19363
rect 12667 19329 12676 19363
rect 12624 19320 12676 19329
rect 14096 19363 14148 19372
rect 14096 19329 14105 19363
rect 14105 19329 14139 19363
rect 14139 19329 14148 19363
rect 14096 19320 14148 19329
rect 14188 19363 14240 19372
rect 14188 19329 14197 19363
rect 14197 19329 14231 19363
rect 14231 19329 14240 19363
rect 14188 19320 14240 19329
rect 14464 19320 14516 19372
rect 2412 19295 2464 19304
rect 2412 19261 2421 19295
rect 2421 19261 2455 19295
rect 2455 19261 2464 19295
rect 2412 19252 2464 19261
rect 4896 19252 4948 19304
rect 5356 19252 5408 19304
rect 5632 19252 5684 19304
rect 6184 19252 6236 19304
rect 6460 19252 6512 19304
rect 7748 19295 7800 19304
rect 7748 19261 7757 19295
rect 7757 19261 7791 19295
rect 7791 19261 7800 19295
rect 7748 19252 7800 19261
rect 8024 19252 8076 19304
rect 12348 19295 12400 19304
rect 12348 19261 12357 19295
rect 12357 19261 12391 19295
rect 12391 19261 12400 19295
rect 12348 19252 12400 19261
rect 12440 19295 12492 19304
rect 12440 19261 12449 19295
rect 12449 19261 12483 19295
rect 12483 19261 12492 19295
rect 12440 19252 12492 19261
rect 13176 19252 13228 19304
rect 14280 19252 14332 19304
rect 14372 19295 14424 19304
rect 14372 19261 14381 19295
rect 14381 19261 14415 19295
rect 14415 19261 14424 19295
rect 14372 19252 14424 19261
rect 15108 19252 15160 19304
rect 15660 19295 15712 19304
rect 15660 19261 15669 19295
rect 15669 19261 15703 19295
rect 15703 19261 15712 19295
rect 15660 19252 15712 19261
rect 15936 19329 15945 19346
rect 15945 19329 15979 19346
rect 15979 19329 15988 19346
rect 15936 19294 15988 19329
rect 17684 19363 17736 19372
rect 17684 19329 17693 19363
rect 17693 19329 17727 19363
rect 17727 19329 17736 19363
rect 17684 19320 17736 19329
rect 17592 19252 17644 19304
rect 17868 19295 17920 19304
rect 17868 19261 17877 19295
rect 17877 19261 17911 19295
rect 17911 19261 17920 19295
rect 17868 19252 17920 19261
rect 17960 19295 18012 19304
rect 17960 19261 17969 19295
rect 17969 19261 18003 19295
rect 18003 19261 18012 19295
rect 17960 19252 18012 19261
rect 6644 19184 6696 19236
rect 2596 19159 2648 19168
rect 2596 19125 2605 19159
rect 2605 19125 2639 19159
rect 2639 19125 2648 19159
rect 2596 19116 2648 19125
rect 7656 19116 7708 19168
rect 12716 19227 12768 19236
rect 12716 19193 12725 19227
rect 12725 19193 12759 19227
rect 12759 19193 12768 19227
rect 12716 19184 12768 19193
rect 12808 19227 12860 19236
rect 12808 19193 12817 19227
rect 12817 19193 12851 19227
rect 12851 19193 12860 19227
rect 12808 19184 12860 19193
rect 12992 19184 13044 19236
rect 15660 19116 15712 19168
rect 19156 19252 19208 19304
rect 19616 19295 19668 19304
rect 19616 19261 19625 19295
rect 19625 19261 19659 19295
rect 19659 19261 19668 19295
rect 19616 19252 19668 19261
rect 19892 19184 19944 19236
rect 20444 19184 20496 19236
rect 18604 19159 18656 19168
rect 18604 19125 18613 19159
rect 18613 19125 18647 19159
rect 18647 19125 18656 19159
rect 18604 19116 18656 19125
rect 19524 19159 19576 19168
rect 19524 19125 19533 19159
rect 19533 19125 19567 19159
rect 19567 19125 19576 19159
rect 19524 19116 19576 19125
rect 7882 19014 7934 19066
rect 7946 19014 7998 19066
rect 8010 19014 8062 19066
rect 8074 19014 8126 19066
rect 14782 19014 14834 19066
rect 14846 19014 14898 19066
rect 14910 19014 14962 19066
rect 14974 19014 15026 19066
rect 12716 18912 12768 18964
rect 6000 18819 6052 18828
rect 6000 18785 6009 18819
rect 6009 18785 6043 18819
rect 6043 18785 6052 18819
rect 6000 18776 6052 18785
rect 6920 18776 6972 18828
rect 7380 18819 7432 18828
rect 7380 18785 7389 18819
rect 7389 18785 7423 18819
rect 7423 18785 7432 18819
rect 7380 18776 7432 18785
rect 7564 18776 7616 18828
rect 11704 18819 11756 18828
rect 11704 18785 11713 18819
rect 11713 18785 11747 18819
rect 11747 18785 11756 18819
rect 11704 18776 11756 18785
rect 12808 18844 12860 18896
rect 13176 18912 13228 18964
rect 13728 18844 13780 18896
rect 16304 18844 16356 18896
rect 20720 18844 20772 18896
rect 11980 18819 12032 18828
rect 11980 18785 11989 18819
rect 11989 18785 12023 18819
rect 12023 18785 12032 18819
rect 11980 18776 12032 18785
rect 12256 18819 12308 18828
rect 12256 18785 12265 18819
rect 12265 18785 12299 18819
rect 12299 18785 12308 18819
rect 12256 18776 12308 18785
rect 12992 18776 13044 18828
rect 13820 18819 13872 18828
rect 13820 18785 13829 18819
rect 13829 18785 13863 18819
rect 13863 18785 13872 18819
rect 13820 18776 13872 18785
rect 17316 18776 17368 18828
rect 17868 18776 17920 18828
rect 18788 18776 18840 18828
rect 19064 18819 19116 18828
rect 19064 18785 19073 18819
rect 19073 18785 19107 18819
rect 19107 18785 19116 18819
rect 19064 18776 19116 18785
rect 7748 18708 7800 18760
rect 8116 18708 8168 18760
rect 15568 18708 15620 18760
rect 5356 18572 5408 18624
rect 7012 18572 7064 18624
rect 7748 18572 7800 18624
rect 8208 18572 8260 18624
rect 15108 18572 15160 18624
rect 16948 18572 17000 18624
rect 17408 18572 17460 18624
rect 17684 18615 17736 18624
rect 17684 18581 17693 18615
rect 17693 18581 17727 18615
rect 17727 18581 17736 18615
rect 17684 18572 17736 18581
rect 4432 18470 4484 18522
rect 4496 18470 4548 18522
rect 4560 18470 4612 18522
rect 4624 18470 4676 18522
rect 11332 18470 11384 18522
rect 11396 18470 11448 18522
rect 11460 18470 11512 18522
rect 11524 18470 11576 18522
rect 18232 18470 18284 18522
rect 18296 18470 18348 18522
rect 18360 18470 18412 18522
rect 18424 18470 18476 18522
rect 6644 18368 6696 18420
rect 12072 18411 12124 18420
rect 12072 18377 12081 18411
rect 12081 18377 12115 18411
rect 12115 18377 12124 18411
rect 12072 18368 12124 18377
rect 12256 18368 12308 18420
rect 12808 18368 12860 18420
rect 16028 18368 16080 18420
rect 17316 18411 17368 18420
rect 17316 18377 17325 18411
rect 17325 18377 17359 18411
rect 17359 18377 17368 18411
rect 17316 18368 17368 18377
rect 17960 18368 18012 18420
rect 18788 18411 18840 18420
rect 18788 18377 18797 18411
rect 18797 18377 18831 18411
rect 18831 18377 18840 18411
rect 18788 18368 18840 18377
rect 4896 18164 4948 18216
rect 5356 18207 5408 18216
rect 5356 18173 5365 18207
rect 5365 18173 5399 18207
rect 5399 18173 5408 18207
rect 5356 18164 5408 18173
rect 6184 18300 6236 18352
rect 7656 18300 7708 18352
rect 8300 18232 8352 18284
rect 8852 18275 8904 18284
rect 8852 18241 8861 18275
rect 8861 18241 8895 18275
rect 8895 18241 8904 18275
rect 8852 18232 8904 18241
rect 19245 18300 19297 18352
rect 19524 18300 19576 18352
rect 9588 18232 9640 18284
rect 11980 18232 12032 18284
rect 7012 18207 7064 18216
rect 7012 18173 7021 18207
rect 7021 18173 7055 18207
rect 7055 18173 7064 18207
rect 7012 18164 7064 18173
rect 4620 18096 4672 18148
rect 5540 18139 5592 18148
rect 5540 18105 5549 18139
rect 5549 18105 5583 18139
rect 5583 18105 5592 18139
rect 5540 18096 5592 18105
rect 6092 18096 6144 18148
rect 6736 18096 6788 18148
rect 4988 18028 5040 18080
rect 6184 18028 6236 18080
rect 7288 18028 7340 18080
rect 7564 18028 7616 18080
rect 8116 18207 8168 18216
rect 8116 18173 8125 18207
rect 8125 18173 8159 18207
rect 8159 18173 8168 18207
rect 8392 18207 8444 18216
rect 8116 18164 8168 18173
rect 8392 18173 8401 18207
rect 8401 18173 8435 18207
rect 8435 18173 8444 18207
rect 8392 18164 8444 18173
rect 8300 18096 8352 18148
rect 9772 18164 9824 18216
rect 10508 18164 10560 18216
rect 11796 18164 11848 18216
rect 14096 18232 14148 18284
rect 17684 18232 17736 18284
rect 12164 18096 12216 18148
rect 14280 18164 14332 18216
rect 16212 18207 16264 18216
rect 16212 18173 16221 18207
rect 16221 18173 16255 18207
rect 16255 18173 16264 18207
rect 16212 18164 16264 18173
rect 17500 18207 17552 18216
rect 14096 18096 14148 18148
rect 16120 18096 16172 18148
rect 17500 18173 17509 18207
rect 17509 18173 17543 18207
rect 17543 18173 17552 18207
rect 17500 18164 17552 18173
rect 19616 18232 19668 18284
rect 19156 18207 19208 18216
rect 17592 18096 17644 18148
rect 8668 18028 8720 18080
rect 9772 18028 9824 18080
rect 10048 18071 10100 18080
rect 10048 18037 10057 18071
rect 10057 18037 10091 18071
rect 10091 18037 10100 18071
rect 10048 18028 10100 18037
rect 19156 18173 19165 18207
rect 19165 18173 19199 18207
rect 19199 18173 19208 18207
rect 19156 18164 19208 18173
rect 19524 18207 19576 18216
rect 19064 18096 19116 18148
rect 19248 18028 19300 18080
rect 19524 18173 19533 18207
rect 19533 18173 19567 18207
rect 19567 18173 19576 18207
rect 19524 18164 19576 18173
rect 20628 18164 20680 18216
rect 20720 18028 20772 18080
rect 20812 18028 20864 18080
rect 7882 17926 7934 17978
rect 7946 17926 7998 17978
rect 8010 17926 8062 17978
rect 8074 17926 8126 17978
rect 14782 17926 14834 17978
rect 14846 17926 14898 17978
rect 14910 17926 14962 17978
rect 14974 17926 15026 17978
rect 6000 17824 6052 17876
rect 4620 17756 4672 17808
rect 4988 17756 5040 17808
rect 6644 17756 6696 17808
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 4160 17688 4212 17740
rect 6092 17688 6144 17740
rect 7196 17756 7248 17808
rect 7564 17756 7616 17808
rect 8208 17824 8260 17876
rect 8852 17824 8904 17876
rect 12624 17824 12676 17876
rect 13912 17824 13964 17876
rect 9772 17799 9824 17808
rect 9772 17765 9781 17799
rect 9781 17765 9815 17799
rect 9815 17765 9824 17799
rect 9772 17756 9824 17765
rect 10048 17756 10100 17808
rect 11796 17756 11848 17808
rect 7656 17731 7708 17740
rect 7656 17697 7665 17731
rect 7665 17697 7699 17731
rect 7699 17697 7708 17731
rect 7656 17688 7708 17697
rect 7748 17731 7800 17740
rect 7748 17697 7758 17731
rect 7758 17697 7792 17731
rect 7792 17697 7800 17731
rect 7748 17688 7800 17697
rect 7196 17620 7248 17672
rect 7380 17620 7432 17672
rect 8484 17688 8536 17740
rect 9496 17731 9548 17740
rect 9496 17697 9505 17731
rect 9505 17697 9539 17731
rect 9539 17697 9548 17731
rect 9496 17688 9548 17697
rect 11980 17731 12032 17740
rect 11980 17697 11989 17731
rect 11989 17697 12023 17731
rect 12023 17697 12032 17731
rect 11980 17688 12032 17697
rect 12164 17756 12216 17808
rect 13820 17756 13872 17808
rect 13636 17688 13688 17740
rect 16212 17688 16264 17740
rect 16396 17688 16448 17740
rect 17500 17688 17552 17740
rect 19340 17688 19392 17740
rect 8024 17620 8076 17672
rect 12072 17663 12124 17672
rect 12072 17629 12081 17663
rect 12081 17629 12115 17663
rect 12115 17629 12124 17663
rect 12072 17620 12124 17629
rect 7656 17552 7708 17604
rect 13820 17620 13872 17672
rect 18880 17620 18932 17672
rect 20260 17731 20312 17740
rect 20260 17697 20269 17731
rect 20269 17697 20303 17731
rect 20303 17697 20312 17731
rect 20260 17688 20312 17697
rect 20444 17688 20496 17740
rect 14096 17552 14148 17604
rect 2320 17484 2372 17536
rect 6092 17484 6144 17536
rect 8300 17484 8352 17536
rect 8668 17484 8720 17536
rect 9588 17484 9640 17536
rect 14004 17484 14056 17536
rect 17316 17484 17368 17536
rect 18972 17527 19024 17536
rect 18972 17493 18981 17527
rect 18981 17493 19015 17527
rect 19015 17493 19024 17527
rect 18972 17484 19024 17493
rect 19616 17484 19668 17536
rect 4432 17382 4484 17434
rect 4496 17382 4548 17434
rect 4560 17382 4612 17434
rect 4624 17382 4676 17434
rect 11332 17382 11384 17434
rect 11396 17382 11448 17434
rect 11460 17382 11512 17434
rect 11524 17382 11576 17434
rect 18232 17382 18284 17434
rect 18296 17382 18348 17434
rect 18360 17382 18412 17434
rect 18424 17382 18476 17434
rect 8024 17323 8076 17332
rect 8024 17289 8033 17323
rect 8033 17289 8067 17323
rect 8067 17289 8076 17323
rect 8024 17280 8076 17289
rect 7012 17212 7064 17264
rect 7104 17187 7156 17196
rect 7104 17153 7113 17187
rect 7113 17153 7147 17187
rect 7147 17153 7156 17187
rect 7104 17144 7156 17153
rect 7288 17212 7340 17264
rect 6000 17076 6052 17128
rect 6736 17008 6788 17060
rect 7380 17076 7432 17128
rect 7564 17076 7616 17128
rect 8300 17280 8352 17332
rect 11888 17280 11940 17332
rect 19064 17280 19116 17332
rect 20260 17280 20312 17332
rect 8668 17119 8720 17128
rect 7656 17008 7708 17060
rect 8668 17085 8677 17119
rect 8677 17085 8711 17119
rect 8711 17085 8720 17119
rect 8668 17076 8720 17085
rect 15568 17076 15620 17128
rect 17408 17076 17460 17128
rect 17592 17119 17644 17128
rect 17592 17085 17601 17119
rect 17601 17085 17635 17119
rect 17635 17085 17644 17119
rect 18604 17144 18656 17196
rect 19248 17144 19300 17196
rect 19616 17187 19668 17196
rect 19616 17153 19625 17187
rect 19625 17153 19659 17187
rect 19659 17153 19668 17187
rect 19616 17144 19668 17153
rect 17592 17076 17644 17085
rect 18696 17119 18748 17128
rect 11796 17008 11848 17060
rect 12440 17051 12492 17060
rect 12440 17017 12449 17051
rect 12449 17017 12483 17051
rect 12483 17017 12492 17051
rect 12440 17008 12492 17017
rect 6828 16983 6880 16992
rect 6828 16949 6837 16983
rect 6837 16949 6871 16983
rect 6871 16949 6880 16983
rect 6828 16940 6880 16949
rect 8392 16940 8444 16992
rect 13912 16940 13964 16992
rect 15292 17008 15344 17060
rect 17684 17051 17736 17060
rect 17684 17017 17693 17051
rect 17693 17017 17727 17051
rect 17727 17017 17736 17051
rect 17684 17008 17736 17017
rect 15752 16940 15804 16992
rect 16396 16940 16448 16992
rect 16580 16940 16632 16992
rect 17500 16940 17552 16992
rect 18696 17085 18705 17119
rect 18705 17085 18739 17119
rect 18739 17085 18748 17119
rect 18696 17076 18748 17085
rect 19340 17119 19392 17128
rect 19340 17085 19349 17119
rect 19349 17085 19383 17119
rect 19383 17085 19392 17119
rect 19340 17076 19392 17085
rect 18972 17008 19024 17060
rect 20628 17008 20680 17060
rect 19064 16940 19116 16992
rect 7882 16838 7934 16890
rect 7946 16838 7998 16890
rect 8010 16838 8062 16890
rect 8074 16838 8126 16890
rect 14782 16838 14834 16890
rect 14846 16838 14898 16890
rect 14910 16838 14962 16890
rect 14974 16838 15026 16890
rect 2412 16736 2464 16788
rect 4252 16736 4304 16788
rect 11888 16736 11940 16788
rect 12164 16736 12216 16788
rect 13636 16736 13688 16788
rect 15292 16779 15344 16788
rect 12440 16668 12492 16720
rect 12808 16668 12860 16720
rect 15292 16745 15301 16779
rect 15301 16745 15335 16779
rect 15335 16745 15344 16779
rect 15292 16736 15344 16745
rect 16580 16711 16632 16720
rect 16580 16677 16589 16711
rect 16589 16677 16623 16711
rect 16623 16677 16632 16711
rect 16580 16668 16632 16677
rect 17316 16668 17368 16720
rect 18696 16736 18748 16788
rect 20628 16736 20680 16788
rect 1676 16643 1728 16652
rect 1676 16609 1685 16643
rect 1685 16609 1719 16643
rect 1719 16609 1728 16643
rect 1676 16600 1728 16609
rect 2320 16643 2372 16652
rect 2320 16609 2329 16643
rect 2329 16609 2363 16643
rect 2363 16609 2372 16643
rect 2320 16600 2372 16609
rect 6092 16600 6144 16652
rect 7656 16600 7708 16652
rect 11796 16643 11848 16652
rect 11796 16609 11805 16643
rect 11805 16609 11839 16643
rect 11839 16609 11848 16643
rect 11796 16600 11848 16609
rect 18972 16668 19024 16720
rect 13636 16643 13688 16652
rect 13636 16609 13645 16643
rect 13645 16609 13679 16643
rect 13679 16609 13688 16643
rect 13636 16600 13688 16609
rect 13912 16600 13964 16652
rect 14372 16600 14424 16652
rect 14648 16600 14700 16652
rect 15200 16600 15252 16652
rect 15476 16600 15528 16652
rect 15568 16600 15620 16652
rect 18880 16643 18932 16652
rect 18880 16609 18889 16643
rect 18889 16609 18923 16643
rect 18923 16609 18932 16643
rect 18880 16600 18932 16609
rect 19064 16600 19116 16652
rect 20904 16600 20956 16652
rect 13820 16507 13872 16516
rect 13820 16473 13829 16507
rect 13829 16473 13863 16507
rect 13863 16473 13872 16507
rect 13820 16464 13872 16473
rect 4432 16294 4484 16346
rect 4496 16294 4548 16346
rect 4560 16294 4612 16346
rect 4624 16294 4676 16346
rect 11332 16294 11384 16346
rect 11396 16294 11448 16346
rect 11460 16294 11512 16346
rect 11524 16294 11576 16346
rect 18232 16294 18284 16346
rect 18296 16294 18348 16346
rect 18360 16294 18412 16346
rect 18424 16294 18476 16346
rect 11796 16192 11848 16244
rect 12808 16235 12860 16244
rect 12808 16201 12817 16235
rect 12817 16201 12851 16235
rect 12851 16201 12860 16235
rect 12808 16192 12860 16201
rect 19156 16235 19208 16244
rect 19156 16201 19165 16235
rect 19165 16201 19199 16235
rect 19199 16201 19208 16235
rect 19156 16192 19208 16201
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 7564 16124 7616 16176
rect 17684 16124 17736 16176
rect 4160 16056 4212 16108
rect 5724 16056 5776 16108
rect 7472 16056 7524 16108
rect 8852 16056 8904 16108
rect 9680 16056 9732 16108
rect 2136 15988 2188 16040
rect 7104 16031 7156 16040
rect 7104 15997 7113 16031
rect 7113 15997 7147 16031
rect 7147 15997 7156 16031
rect 9036 16031 9088 16040
rect 7104 15988 7156 15997
rect 9036 15997 9045 16031
rect 9045 15997 9079 16031
rect 9079 15997 9088 16031
rect 9036 15988 9088 15997
rect 10508 16031 10560 16040
rect 10508 15997 10517 16031
rect 10517 15997 10551 16031
rect 10551 15997 10560 16031
rect 10508 15988 10560 15997
rect 10968 15988 11020 16040
rect 4344 15920 4396 15972
rect 4988 15852 5040 15904
rect 5632 15852 5684 15904
rect 6368 15852 6420 15904
rect 7288 15852 7340 15904
rect 9772 15852 9824 15904
rect 10784 15852 10836 15904
rect 16948 16056 17000 16108
rect 13820 15988 13872 16040
rect 14372 16031 14424 16040
rect 14372 15997 14381 16031
rect 14381 15997 14415 16031
rect 14415 15997 14424 16031
rect 14372 15988 14424 15997
rect 17592 15988 17644 16040
rect 18696 15988 18748 16040
rect 14004 15920 14056 15972
rect 15476 15920 15528 15972
rect 18604 15920 18656 15972
rect 13636 15852 13688 15904
rect 17408 15852 17460 15904
rect 20904 16031 20956 16040
rect 20904 15997 20913 16031
rect 20913 15997 20947 16031
rect 20947 15997 20956 16031
rect 20904 15988 20956 15997
rect 19984 15852 20036 15904
rect 7882 15750 7934 15802
rect 7946 15750 7998 15802
rect 8010 15750 8062 15802
rect 8074 15750 8126 15802
rect 14782 15750 14834 15802
rect 14846 15750 14898 15802
rect 14910 15750 14962 15802
rect 14974 15750 15026 15802
rect 4344 15648 4396 15700
rect 4988 15648 5040 15700
rect 7196 15648 7248 15700
rect 14096 15648 14148 15700
rect 17592 15648 17644 15700
rect 20904 15691 20956 15700
rect 20904 15657 20913 15691
rect 20913 15657 20947 15691
rect 20947 15657 20956 15691
rect 20904 15648 20956 15657
rect 5724 15580 5776 15632
rect 9772 15623 9824 15632
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 4896 15512 4948 15564
rect 5264 15555 5316 15564
rect 5264 15521 5273 15555
rect 5273 15521 5307 15555
rect 5307 15521 5316 15555
rect 5264 15512 5316 15521
rect 5632 15512 5684 15564
rect 6368 15555 6420 15564
rect 6368 15521 6377 15555
rect 6377 15521 6411 15555
rect 6411 15521 6420 15555
rect 6368 15512 6420 15521
rect 7012 15512 7064 15564
rect 7196 15555 7248 15564
rect 7196 15521 7205 15555
rect 7205 15521 7239 15555
rect 7239 15521 7248 15555
rect 7196 15512 7248 15521
rect 7288 15555 7340 15564
rect 9772 15589 9781 15623
rect 9781 15589 9815 15623
rect 9815 15589 9824 15623
rect 9772 15580 9824 15589
rect 10784 15580 10836 15632
rect 7288 15521 7302 15555
rect 7302 15521 7336 15555
rect 7336 15521 7340 15555
rect 7288 15512 7340 15521
rect 8208 15555 8260 15564
rect 8208 15521 8217 15555
rect 8217 15521 8251 15555
rect 8251 15521 8260 15555
rect 8208 15512 8260 15521
rect 8300 15555 8352 15564
rect 8300 15521 8309 15555
rect 8309 15521 8343 15555
rect 8343 15521 8352 15555
rect 8300 15512 8352 15521
rect 8944 15512 8996 15564
rect 9496 15555 9548 15564
rect 9496 15521 9505 15555
rect 9505 15521 9539 15555
rect 9539 15521 9548 15555
rect 9496 15512 9548 15521
rect 17040 15555 17092 15564
rect 8576 15444 8628 15496
rect 17040 15521 17049 15555
rect 17049 15521 17083 15555
rect 17083 15521 17092 15555
rect 17040 15512 17092 15521
rect 18788 15512 18840 15564
rect 21088 15555 21140 15564
rect 21088 15521 21097 15555
rect 21097 15521 21131 15555
rect 21131 15521 21140 15555
rect 21088 15512 21140 15521
rect 15292 15487 15344 15496
rect 8852 15376 8904 15428
rect 15292 15453 15301 15487
rect 15301 15453 15335 15487
rect 15335 15453 15344 15487
rect 15292 15444 15344 15453
rect 15384 15487 15436 15496
rect 15384 15453 15393 15487
rect 15393 15453 15427 15487
rect 15427 15453 15436 15487
rect 15384 15444 15436 15453
rect 1860 15308 1912 15360
rect 7472 15351 7524 15360
rect 7472 15317 7481 15351
rect 7481 15317 7515 15351
rect 7515 15317 7524 15351
rect 7472 15308 7524 15317
rect 9956 15308 10008 15360
rect 10140 15308 10192 15360
rect 14096 15308 14148 15360
rect 15568 15308 15620 15360
rect 17960 15308 18012 15360
rect 4432 15206 4484 15258
rect 4496 15206 4548 15258
rect 4560 15206 4612 15258
rect 4624 15206 4676 15258
rect 11332 15206 11384 15258
rect 11396 15206 11448 15258
rect 11460 15206 11512 15258
rect 11524 15206 11576 15258
rect 18232 15206 18284 15258
rect 18296 15206 18348 15258
rect 18360 15206 18412 15258
rect 18424 15206 18476 15258
rect 5264 15104 5316 15156
rect 5724 15104 5776 15156
rect 6644 15104 6696 15156
rect 8944 15147 8996 15156
rect 7012 15036 7064 15088
rect 8944 15113 8953 15147
rect 8953 15113 8987 15147
rect 8987 15113 8996 15147
rect 8944 15104 8996 15113
rect 9680 15104 9732 15156
rect 14004 15104 14056 15156
rect 15292 15104 15344 15156
rect 17040 15104 17092 15156
rect 17500 15147 17552 15156
rect 17500 15113 17509 15147
rect 17509 15113 17543 15147
rect 17543 15113 17552 15147
rect 17500 15104 17552 15113
rect 10968 15036 11020 15088
rect 1860 14943 1912 14952
rect 1860 14909 1869 14943
rect 1869 14909 1903 14943
rect 1903 14909 1912 14943
rect 1860 14900 1912 14909
rect 6736 14968 6788 15020
rect 7472 15011 7524 15020
rect 7472 14977 7481 15011
rect 7481 14977 7515 15011
rect 7515 14977 7524 15011
rect 7472 14968 7524 14977
rect 7564 14968 7616 15020
rect 9956 15011 10008 15020
rect 6828 14943 6880 14952
rect 2044 14807 2096 14816
rect 2044 14773 2053 14807
rect 2053 14773 2087 14807
rect 2087 14773 2096 14807
rect 2044 14764 2096 14773
rect 2320 14764 2372 14816
rect 3516 14764 3568 14816
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 6920 14900 6972 14952
rect 6184 14832 6236 14884
rect 7748 14900 7800 14952
rect 9036 14900 9088 14952
rect 9956 14977 9965 15011
rect 9965 14977 9999 15011
rect 9999 14977 10008 15011
rect 9956 14968 10008 14977
rect 6828 14764 6880 14816
rect 7564 14764 7616 14816
rect 9680 14900 9732 14952
rect 15200 15036 15252 15088
rect 15384 15036 15436 15088
rect 14648 14900 14700 14952
rect 15108 14900 15160 14952
rect 17960 14968 18012 15020
rect 10600 14832 10652 14884
rect 17316 14900 17368 14952
rect 18696 14943 18748 14952
rect 11428 14764 11480 14816
rect 12348 14807 12400 14816
rect 12348 14773 12357 14807
rect 12357 14773 12391 14807
rect 12391 14773 12400 14807
rect 12348 14764 12400 14773
rect 14556 14807 14608 14816
rect 14556 14773 14565 14807
rect 14565 14773 14599 14807
rect 14599 14773 14608 14807
rect 14556 14764 14608 14773
rect 16212 14764 16264 14816
rect 18696 14909 18705 14943
rect 18705 14909 18739 14943
rect 18739 14909 18748 14943
rect 18696 14900 18748 14909
rect 19984 14968 20036 15020
rect 19340 14943 19392 14952
rect 19340 14909 19349 14943
rect 19349 14909 19383 14943
rect 19383 14909 19392 14943
rect 19340 14900 19392 14909
rect 18788 14832 18840 14884
rect 19616 14875 19668 14884
rect 19616 14841 19625 14875
rect 19625 14841 19659 14875
rect 19659 14841 19668 14875
rect 19616 14832 19668 14841
rect 20628 14832 20680 14884
rect 19708 14764 19760 14816
rect 20260 14764 20312 14816
rect 7882 14662 7934 14714
rect 7946 14662 7998 14714
rect 8010 14662 8062 14714
rect 8074 14662 8126 14714
rect 14782 14662 14834 14714
rect 14846 14662 14898 14714
rect 14910 14662 14962 14714
rect 14974 14662 15026 14714
rect 6184 14603 6236 14612
rect 6184 14569 6193 14603
rect 6193 14569 6227 14603
rect 6227 14569 6236 14603
rect 6184 14560 6236 14569
rect 5632 14492 5684 14544
rect 6828 14560 6880 14612
rect 7196 14560 7248 14612
rect 8300 14560 8352 14612
rect 9036 14560 9088 14612
rect 9496 14560 9548 14612
rect 10600 14603 10652 14612
rect 10600 14569 10609 14603
rect 10609 14569 10643 14603
rect 10643 14569 10652 14603
rect 10600 14560 10652 14569
rect 12348 14560 12400 14612
rect 14648 14560 14700 14612
rect 7104 14492 7156 14544
rect 7564 14492 7616 14544
rect 7748 14492 7800 14544
rect 2320 14467 2372 14476
rect 2320 14433 2329 14467
rect 2329 14433 2363 14467
rect 2363 14433 2372 14467
rect 2320 14424 2372 14433
rect 6736 14467 6788 14476
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 2780 14399 2832 14408
rect 2780 14365 2789 14399
rect 2789 14365 2823 14399
rect 2823 14365 2832 14399
rect 3148 14399 3200 14408
rect 2780 14356 2832 14365
rect 3148 14365 3157 14399
rect 3157 14365 3191 14399
rect 3191 14365 3200 14399
rect 3148 14356 3200 14365
rect 6736 14433 6745 14467
rect 6745 14433 6779 14467
rect 6779 14433 6788 14467
rect 6736 14424 6788 14433
rect 7012 14424 7064 14476
rect 7472 14424 7524 14476
rect 8208 14424 8260 14476
rect 9680 14492 9732 14544
rect 11428 14535 11480 14544
rect 10140 14424 10192 14476
rect 11428 14501 11437 14535
rect 11437 14501 11471 14535
rect 11471 14501 11480 14535
rect 11428 14492 11480 14501
rect 14556 14492 14608 14544
rect 15016 14535 15068 14544
rect 15016 14501 15025 14535
rect 15025 14501 15059 14535
rect 15059 14501 15068 14535
rect 15016 14492 15068 14501
rect 15200 14560 15252 14612
rect 15752 14560 15804 14612
rect 19984 14603 20036 14612
rect 19984 14569 19993 14603
rect 19993 14569 20027 14603
rect 20027 14569 20036 14603
rect 19984 14560 20036 14569
rect 20260 14560 20312 14612
rect 17040 14492 17092 14544
rect 10784 14424 10836 14476
rect 15292 14467 15344 14476
rect 6644 14356 6696 14408
rect 11152 14399 11204 14408
rect 11152 14365 11161 14399
rect 11161 14365 11195 14399
rect 11195 14365 11204 14399
rect 11152 14356 11204 14365
rect 15292 14433 15301 14467
rect 15301 14433 15335 14467
rect 15335 14433 15344 14467
rect 15292 14424 15344 14433
rect 16212 14467 16264 14476
rect 16212 14433 16221 14467
rect 16221 14433 16255 14467
rect 16255 14433 16264 14467
rect 16212 14424 16264 14433
rect 16948 14467 17000 14476
rect 16948 14433 16957 14467
rect 16957 14433 16991 14467
rect 16991 14433 17000 14467
rect 16948 14424 17000 14433
rect 17960 14424 18012 14476
rect 18880 14492 18932 14544
rect 18604 14467 18656 14476
rect 15476 14356 15528 14408
rect 17408 14356 17460 14408
rect 17500 14356 17552 14408
rect 18604 14433 18613 14467
rect 18613 14433 18647 14467
rect 18647 14433 18656 14467
rect 18604 14424 18656 14433
rect 19524 14424 19576 14476
rect 20260 14424 20312 14476
rect 18788 14356 18840 14408
rect 17316 14288 17368 14340
rect 2320 14263 2372 14272
rect 2320 14229 2329 14263
rect 2329 14229 2363 14263
rect 2363 14229 2372 14263
rect 2320 14220 2372 14229
rect 3516 14220 3568 14272
rect 12900 14263 12952 14272
rect 12900 14229 12909 14263
rect 12909 14229 12943 14263
rect 12943 14229 12952 14263
rect 12900 14220 12952 14229
rect 14280 14220 14332 14272
rect 17960 14288 18012 14340
rect 18052 14220 18104 14272
rect 4432 14118 4484 14170
rect 4496 14118 4548 14170
rect 4560 14118 4612 14170
rect 4624 14118 4676 14170
rect 11332 14118 11384 14170
rect 11396 14118 11448 14170
rect 11460 14118 11512 14170
rect 11524 14118 11576 14170
rect 18232 14118 18284 14170
rect 18296 14118 18348 14170
rect 18360 14118 18412 14170
rect 18424 14118 18476 14170
rect 1952 14059 2004 14068
rect 1952 14025 1961 14059
rect 1961 14025 1995 14059
rect 1995 14025 2004 14059
rect 1952 14016 2004 14025
rect 2412 13923 2464 13932
rect 2412 13889 2421 13923
rect 2421 13889 2455 13923
rect 2455 13889 2464 13923
rect 2412 13880 2464 13889
rect 4804 14016 4856 14068
rect 8576 14059 8628 14068
rect 8576 14025 8585 14059
rect 8585 14025 8619 14059
rect 8619 14025 8628 14059
rect 8576 14016 8628 14025
rect 15016 14016 15068 14068
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 17500 14059 17552 14068
rect 17500 14025 17509 14059
rect 17509 14025 17543 14059
rect 17543 14025 17552 14059
rect 17500 14016 17552 14025
rect 19616 14016 19668 14068
rect 20628 14016 20680 14068
rect 3148 13923 3200 13932
rect 2228 13812 2280 13864
rect 3148 13889 3157 13923
rect 3157 13889 3191 13923
rect 3191 13889 3200 13923
rect 16948 13948 17000 14000
rect 3148 13880 3200 13889
rect 12256 13880 12308 13932
rect 14280 13923 14332 13932
rect 14280 13889 14289 13923
rect 14289 13889 14323 13923
rect 14323 13889 14332 13923
rect 14280 13880 14332 13889
rect 17316 13923 17368 13932
rect 17316 13889 17325 13923
rect 17325 13889 17359 13923
rect 17359 13889 17368 13923
rect 17316 13880 17368 13889
rect 2780 13812 2832 13864
rect 8944 13812 8996 13864
rect 10324 13812 10376 13864
rect 11152 13812 11204 13864
rect 11980 13812 12032 13864
rect 14004 13855 14056 13864
rect 14004 13821 14013 13855
rect 14013 13821 14047 13855
rect 14047 13821 14056 13855
rect 14004 13812 14056 13821
rect 17868 13812 17920 13864
rect 18052 13855 18104 13864
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 19248 13880 19300 13932
rect 19524 13812 19576 13864
rect 19708 13855 19760 13864
rect 19708 13821 19717 13855
rect 19717 13821 19751 13855
rect 19751 13821 19760 13855
rect 19708 13812 19760 13821
rect 20720 13812 20772 13864
rect 20996 13812 21048 13864
rect 5632 13744 5684 13796
rect 3516 13719 3568 13728
rect 3516 13685 3525 13719
rect 3525 13685 3559 13719
rect 3559 13685 3568 13719
rect 3516 13676 3568 13685
rect 5448 13676 5500 13728
rect 10692 13744 10744 13796
rect 15568 13744 15620 13796
rect 20260 13744 20312 13796
rect 9864 13719 9916 13728
rect 9864 13685 9873 13719
rect 9873 13685 9907 13719
rect 9907 13685 9916 13719
rect 9864 13676 9916 13685
rect 18604 13676 18656 13728
rect 7882 13574 7934 13626
rect 7946 13574 7998 13626
rect 8010 13574 8062 13626
rect 8074 13574 8126 13626
rect 14782 13574 14834 13626
rect 14846 13574 14898 13626
rect 14910 13574 14962 13626
rect 14974 13574 15026 13626
rect 2320 13472 2372 13524
rect 2780 13472 2832 13524
rect 6920 13472 6972 13524
rect 7748 13472 7800 13524
rect 9864 13515 9916 13524
rect 9864 13481 9873 13515
rect 9873 13481 9907 13515
rect 9907 13481 9916 13515
rect 9864 13472 9916 13481
rect 15108 13472 15160 13524
rect 15568 13515 15620 13524
rect 15568 13481 15577 13515
rect 15577 13481 15611 13515
rect 15611 13481 15620 13515
rect 15568 13472 15620 13481
rect 1952 13336 2004 13388
rect 4252 13404 4304 13456
rect 3332 13379 3384 13388
rect 3332 13345 3341 13379
rect 3341 13345 3375 13379
rect 3375 13345 3384 13379
rect 3332 13336 3384 13345
rect 6460 13336 6512 13388
rect 6644 13336 6696 13388
rect 7288 13336 7340 13388
rect 14556 13404 14608 13456
rect 16212 13447 16264 13456
rect 4804 13311 4856 13320
rect 4804 13277 4813 13311
rect 4813 13277 4847 13311
rect 4847 13277 4856 13311
rect 4804 13268 4856 13277
rect 5448 13268 5500 13320
rect 5632 13311 5684 13320
rect 5632 13277 5641 13311
rect 5641 13277 5675 13311
rect 5675 13277 5684 13311
rect 5632 13268 5684 13277
rect 3608 13132 3660 13184
rect 6828 13268 6880 13320
rect 10048 13336 10100 13388
rect 10508 13336 10560 13388
rect 9496 13268 9548 13320
rect 11152 13336 11204 13388
rect 16212 13413 16221 13447
rect 16221 13413 16255 13447
rect 16255 13413 16264 13447
rect 16212 13404 16264 13413
rect 17316 13404 17368 13456
rect 17960 13447 18012 13456
rect 17960 13413 17969 13447
rect 17969 13413 18003 13447
rect 18003 13413 18012 13447
rect 17960 13404 18012 13413
rect 15752 13379 15804 13388
rect 10784 13268 10836 13320
rect 12164 13311 12216 13320
rect 6736 13132 6788 13184
rect 6920 13175 6972 13184
rect 6920 13141 6929 13175
rect 6929 13141 6963 13175
rect 6963 13141 6972 13175
rect 6920 13132 6972 13141
rect 7104 13200 7156 13252
rect 9404 13200 9456 13252
rect 9588 13200 9640 13252
rect 10600 13200 10652 13252
rect 12164 13277 12173 13311
rect 12173 13277 12207 13311
rect 12207 13277 12216 13311
rect 12164 13268 12216 13277
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 12900 13200 12952 13252
rect 13544 13200 13596 13252
rect 14004 13200 14056 13252
rect 17960 13268 18012 13320
rect 19340 13268 19392 13320
rect 7564 13132 7616 13184
rect 10140 13132 10192 13184
rect 12624 13175 12676 13184
rect 12624 13141 12633 13175
rect 12633 13141 12667 13175
rect 12667 13141 12676 13175
rect 12624 13132 12676 13141
rect 4432 13030 4484 13082
rect 4496 13030 4548 13082
rect 4560 13030 4612 13082
rect 4624 13030 4676 13082
rect 11332 13030 11384 13082
rect 11396 13030 11448 13082
rect 11460 13030 11512 13082
rect 11524 13030 11576 13082
rect 18232 13030 18284 13082
rect 18296 13030 18348 13082
rect 18360 13030 18412 13082
rect 18424 13030 18476 13082
rect 1492 12971 1544 12980
rect 1492 12937 1501 12971
rect 1501 12937 1535 12971
rect 1535 12937 1544 12971
rect 1492 12928 1544 12937
rect 3332 12928 3384 12980
rect 9404 12971 9456 12980
rect 9404 12937 9413 12971
rect 9413 12937 9447 12971
rect 9447 12937 9456 12971
rect 9404 12928 9456 12937
rect 10692 12928 10744 12980
rect 6644 12860 6696 12912
rect 3608 12835 3660 12844
rect 3608 12801 3617 12835
rect 3617 12801 3651 12835
rect 3651 12801 3660 12835
rect 3608 12792 3660 12801
rect 7104 12792 7156 12844
rect 9496 12835 9548 12844
rect 4344 12724 4396 12776
rect 6828 12767 6880 12776
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 7564 12724 7616 12776
rect 7656 12724 7708 12776
rect 2412 12656 2464 12708
rect 3148 12699 3200 12708
rect 3148 12665 3157 12699
rect 3157 12665 3191 12699
rect 3191 12665 3200 12699
rect 3148 12656 3200 12665
rect 8392 12699 8444 12708
rect 8392 12665 8401 12699
rect 8401 12665 8435 12699
rect 8435 12665 8444 12699
rect 8392 12656 8444 12665
rect 9496 12801 9505 12835
rect 9505 12801 9539 12835
rect 9539 12801 9548 12835
rect 9496 12792 9548 12801
rect 11152 12860 11204 12912
rect 10784 12792 10836 12844
rect 12256 12835 12308 12844
rect 12256 12801 12265 12835
rect 12265 12801 12299 12835
rect 12299 12801 12308 12835
rect 12256 12792 12308 12801
rect 17960 12792 18012 12844
rect 18604 12792 18656 12844
rect 20260 12835 20312 12844
rect 20260 12801 20269 12835
rect 20269 12801 20303 12835
rect 20303 12801 20312 12835
rect 20260 12792 20312 12801
rect 9404 12767 9456 12776
rect 9404 12733 9413 12767
rect 9413 12733 9447 12767
rect 9447 12733 9456 12767
rect 9404 12724 9456 12733
rect 10600 12724 10652 12776
rect 11152 12767 11204 12776
rect 11152 12733 11161 12767
rect 11161 12733 11195 12767
rect 11195 12733 11204 12767
rect 11152 12724 11204 12733
rect 13544 12767 13596 12776
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 13544 12724 13596 12733
rect 21088 12767 21140 12776
rect 21088 12733 21097 12767
rect 21097 12733 21131 12767
rect 21131 12733 21140 12767
rect 21088 12724 21140 12733
rect 9588 12656 9640 12708
rect 12164 12656 12216 12708
rect 19984 12656 20036 12708
rect 7288 12588 7340 12640
rect 10968 12588 11020 12640
rect 12348 12588 12400 12640
rect 12532 12631 12584 12640
rect 12532 12597 12541 12631
rect 12541 12597 12575 12631
rect 12575 12597 12584 12631
rect 12900 12631 12952 12640
rect 12532 12588 12584 12597
rect 12900 12597 12909 12631
rect 12909 12597 12943 12631
rect 12943 12597 12952 12631
rect 12900 12588 12952 12597
rect 15108 12588 15160 12640
rect 20904 12631 20956 12640
rect 20904 12597 20913 12631
rect 20913 12597 20947 12631
rect 20947 12597 20956 12631
rect 20904 12588 20956 12597
rect 7882 12486 7934 12538
rect 7946 12486 7998 12538
rect 8010 12486 8062 12538
rect 8074 12486 8126 12538
rect 14782 12486 14834 12538
rect 14846 12486 14898 12538
rect 14910 12486 14962 12538
rect 14974 12486 15026 12538
rect 4344 12427 4396 12436
rect 4344 12393 4353 12427
rect 4353 12393 4387 12427
rect 4387 12393 4396 12427
rect 4344 12384 4396 12393
rect 12164 12384 12216 12436
rect 12256 12384 12308 12436
rect 12532 12384 12584 12436
rect 15108 12427 15160 12436
rect 15108 12393 15117 12427
rect 15117 12393 15151 12427
rect 15151 12393 15160 12427
rect 15108 12384 15160 12393
rect 15844 12384 15896 12436
rect 17316 12427 17368 12436
rect 17316 12393 17325 12427
rect 17325 12393 17359 12427
rect 17359 12393 17368 12427
rect 17316 12384 17368 12393
rect 19984 12427 20036 12436
rect 19984 12393 19993 12427
rect 19993 12393 20027 12427
rect 20027 12393 20036 12427
rect 19984 12384 20036 12393
rect 6092 12359 6144 12368
rect 6092 12325 6101 12359
rect 6101 12325 6135 12359
rect 6135 12325 6144 12359
rect 6092 12316 6144 12325
rect 6460 12359 6512 12368
rect 6460 12325 6469 12359
rect 6469 12325 6503 12359
rect 6503 12325 6512 12359
rect 6460 12316 6512 12325
rect 4160 12248 4212 12300
rect 7104 12248 7156 12300
rect 7748 12248 7800 12300
rect 7472 12180 7524 12232
rect 9496 12248 9548 12300
rect 10232 12291 10284 12300
rect 10232 12257 10241 12291
rect 10241 12257 10275 12291
rect 10275 12257 10284 12291
rect 10232 12248 10284 12257
rect 10416 12291 10468 12300
rect 10416 12257 10425 12291
rect 10425 12257 10459 12291
rect 10459 12257 10468 12291
rect 10416 12248 10468 12257
rect 10600 12248 10652 12300
rect 9864 12180 9916 12232
rect 10692 12180 10744 12232
rect 12164 12248 12216 12300
rect 12624 12291 12676 12300
rect 12624 12257 12633 12291
rect 12633 12257 12667 12291
rect 12667 12257 12676 12291
rect 12624 12248 12676 12257
rect 15752 12248 15804 12300
rect 20628 12248 20680 12300
rect 20812 12248 20864 12300
rect 12348 12180 12400 12232
rect 15568 12180 15620 12232
rect 15844 12112 15896 12164
rect 7380 12044 7432 12096
rect 10508 12044 10560 12096
rect 10968 12044 11020 12096
rect 14096 12044 14148 12096
rect 20720 12087 20772 12096
rect 20720 12053 20729 12087
rect 20729 12053 20763 12087
rect 20763 12053 20772 12087
rect 20720 12044 20772 12053
rect 4432 11942 4484 11994
rect 4496 11942 4548 11994
rect 4560 11942 4612 11994
rect 4624 11942 4676 11994
rect 11332 11942 11384 11994
rect 11396 11942 11448 11994
rect 11460 11942 11512 11994
rect 11524 11942 11576 11994
rect 18232 11942 18284 11994
rect 18296 11942 18348 11994
rect 18360 11942 18412 11994
rect 18424 11942 18476 11994
rect 7288 11840 7340 11892
rect 2228 11772 2280 11824
rect 4160 11772 4212 11824
rect 13268 11815 13320 11824
rect 13268 11781 13277 11815
rect 13277 11781 13311 11815
rect 13311 11781 13320 11815
rect 13268 11772 13320 11781
rect 2044 11704 2096 11756
rect 3148 11704 3200 11756
rect 3792 11704 3844 11756
rect 4344 11636 4396 11688
rect 7012 11704 7064 11756
rect 9864 11704 9916 11756
rect 10416 11704 10468 11756
rect 12900 11747 12952 11756
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 15568 11747 15620 11756
rect 7104 11636 7156 11688
rect 8484 11636 8536 11688
rect 6644 11568 6696 11620
rect 2596 11543 2648 11552
rect 2596 11509 2605 11543
rect 2605 11509 2639 11543
rect 2639 11509 2648 11543
rect 2596 11500 2648 11509
rect 4252 11500 4304 11552
rect 7564 11568 7616 11620
rect 8760 11679 8812 11688
rect 8760 11645 8769 11679
rect 8769 11645 8803 11679
rect 8803 11645 8812 11679
rect 8760 11636 8812 11645
rect 10692 11679 10744 11688
rect 10692 11645 10701 11679
rect 10701 11645 10735 11679
rect 10735 11645 10744 11679
rect 10692 11636 10744 11645
rect 13912 11679 13964 11688
rect 9680 11568 9732 11620
rect 10784 11568 10836 11620
rect 7748 11500 7800 11552
rect 9128 11500 9180 11552
rect 13912 11645 13921 11679
rect 13921 11645 13955 11679
rect 13955 11645 13964 11679
rect 13912 11636 13964 11645
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 15568 11704 15620 11713
rect 15660 11704 15712 11756
rect 20812 11704 20864 11756
rect 20720 11636 20772 11688
rect 20904 11679 20956 11688
rect 20904 11645 20913 11679
rect 20913 11645 20947 11679
rect 20947 11645 20956 11679
rect 20904 11636 20956 11645
rect 13728 11543 13780 11552
rect 13728 11509 13737 11543
rect 13737 11509 13771 11543
rect 13771 11509 13780 11543
rect 13728 11500 13780 11509
rect 16396 11500 16448 11552
rect 20720 11543 20772 11552
rect 20720 11509 20729 11543
rect 20729 11509 20763 11543
rect 20763 11509 20772 11543
rect 20720 11500 20772 11509
rect 7882 11398 7934 11450
rect 7946 11398 7998 11450
rect 8010 11398 8062 11450
rect 8074 11398 8126 11450
rect 14782 11398 14834 11450
rect 14846 11398 14898 11450
rect 14910 11398 14962 11450
rect 14974 11398 15026 11450
rect 4160 11296 4212 11348
rect 6460 11296 6512 11348
rect 12164 11296 12216 11348
rect 13268 11339 13320 11348
rect 13268 11305 13277 11339
rect 13277 11305 13311 11339
rect 13311 11305 13320 11339
rect 13268 11296 13320 11305
rect 2320 11160 2372 11212
rect 4252 11203 4304 11212
rect 4252 11169 4261 11203
rect 4261 11169 4295 11203
rect 4295 11169 4304 11203
rect 4252 11160 4304 11169
rect 4344 11160 4396 11212
rect 6460 11160 6512 11212
rect 6920 11160 6972 11212
rect 7840 11203 7892 11212
rect 7840 11169 7849 11203
rect 7849 11169 7883 11203
rect 7883 11169 7892 11203
rect 7840 11160 7892 11169
rect 5448 11092 5500 11144
rect 6092 11092 6144 11144
rect 6644 11135 6696 11144
rect 6644 11101 6653 11135
rect 6653 11101 6687 11135
rect 6687 11101 6696 11135
rect 6644 11092 6696 11101
rect 4160 11024 4212 11076
rect 7012 11092 7064 11144
rect 7196 11092 7248 11144
rect 7564 11135 7616 11144
rect 7564 11101 7573 11135
rect 7573 11101 7607 11135
rect 7607 11101 7616 11135
rect 7564 11092 7616 11101
rect 7656 11135 7708 11144
rect 7656 11101 7665 11135
rect 7665 11101 7699 11135
rect 7699 11101 7708 11135
rect 7656 11092 7708 11101
rect 8760 11160 8812 11212
rect 9312 11160 9364 11212
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9864 11203 9916 11212
rect 9680 11160 9732 11169
rect 9864 11169 9873 11203
rect 9873 11169 9907 11203
rect 9907 11169 9916 11203
rect 9864 11160 9916 11169
rect 10508 11228 10560 11280
rect 10692 11228 10744 11280
rect 20720 11228 20772 11280
rect 12900 11203 12952 11212
rect 12348 11092 12400 11144
rect 12900 11169 12909 11203
rect 12909 11169 12943 11203
rect 12943 11169 12952 11203
rect 12900 11160 12952 11169
rect 13728 11160 13780 11212
rect 16396 11203 16448 11212
rect 16396 11169 16405 11203
rect 16405 11169 16439 11203
rect 16439 11169 16448 11203
rect 16396 11160 16448 11169
rect 16764 11203 16816 11212
rect 16764 11169 16773 11203
rect 16773 11169 16807 11203
rect 16807 11169 16816 11203
rect 16764 11160 16816 11169
rect 15660 11092 15712 11144
rect 2688 10956 2740 11008
rect 13176 11024 13228 11076
rect 7104 10956 7156 11008
rect 7656 10956 7708 11008
rect 8484 10999 8536 11008
rect 8484 10965 8493 10999
rect 8493 10965 8527 10999
rect 8527 10965 8536 10999
rect 8484 10956 8536 10965
rect 15016 10999 15068 11008
rect 15016 10965 15025 10999
rect 15025 10965 15059 10999
rect 15059 10965 15068 10999
rect 15016 10956 15068 10965
rect 4432 10854 4484 10906
rect 4496 10854 4548 10906
rect 4560 10854 4612 10906
rect 4624 10854 4676 10906
rect 11332 10854 11384 10906
rect 11396 10854 11448 10906
rect 11460 10854 11512 10906
rect 11524 10854 11576 10906
rect 18232 10854 18284 10906
rect 18296 10854 18348 10906
rect 18360 10854 18412 10906
rect 18424 10854 18476 10906
rect 3792 10795 3844 10804
rect 3792 10761 3801 10795
rect 3801 10761 3835 10795
rect 3835 10761 3844 10795
rect 3792 10752 3844 10761
rect 6920 10752 6972 10804
rect 7472 10752 7524 10804
rect 8392 10752 8444 10804
rect 8484 10752 8536 10804
rect 10416 10752 10468 10804
rect 13912 10752 13964 10804
rect 20812 10752 20864 10804
rect 7380 10684 7432 10736
rect 2596 10616 2648 10668
rect 8484 10616 8536 10668
rect 2320 10548 2372 10600
rect 2688 10591 2740 10600
rect 2688 10557 2697 10591
rect 2697 10557 2731 10591
rect 2731 10557 2740 10591
rect 2688 10548 2740 10557
rect 4068 10548 4120 10600
rect 8760 10548 8812 10600
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 10876 10684 10928 10736
rect 13176 10659 13228 10668
rect 8484 10480 8536 10532
rect 11704 10548 11756 10600
rect 10508 10523 10560 10532
rect 10508 10489 10530 10523
rect 10530 10489 10560 10523
rect 10508 10480 10560 10489
rect 10968 10480 11020 10532
rect 13176 10625 13185 10659
rect 13185 10625 13219 10659
rect 13219 10625 13228 10659
rect 13176 10616 13228 10625
rect 13360 10659 13412 10668
rect 13360 10625 13369 10659
rect 13369 10625 13403 10659
rect 13403 10625 13412 10659
rect 13360 10616 13412 10625
rect 13268 10548 13320 10600
rect 15016 10684 15068 10736
rect 15476 10591 15528 10600
rect 2964 10412 3016 10464
rect 8668 10412 8720 10464
rect 10600 10412 10652 10464
rect 12532 10455 12584 10464
rect 12532 10421 12541 10455
rect 12541 10421 12575 10455
rect 12575 10421 12584 10455
rect 12532 10412 12584 10421
rect 13820 10455 13872 10464
rect 13820 10421 13829 10455
rect 13829 10421 13863 10455
rect 13863 10421 13872 10455
rect 13820 10412 13872 10421
rect 14648 10412 14700 10464
rect 15476 10557 15485 10591
rect 15485 10557 15519 10591
rect 15519 10557 15528 10591
rect 15476 10548 15528 10557
rect 20904 10591 20956 10600
rect 20904 10557 20913 10591
rect 20913 10557 20947 10591
rect 20947 10557 20956 10591
rect 20904 10548 20956 10557
rect 16764 10480 16816 10532
rect 7882 10310 7934 10362
rect 7946 10310 7998 10362
rect 8010 10310 8062 10362
rect 8074 10310 8126 10362
rect 14782 10310 14834 10362
rect 14846 10310 14898 10362
rect 14910 10310 14962 10362
rect 14974 10310 15026 10362
rect 1492 10251 1544 10260
rect 1492 10217 1501 10251
rect 1501 10217 1535 10251
rect 1535 10217 1544 10251
rect 1492 10208 1544 10217
rect 2320 10251 2372 10260
rect 2320 10217 2329 10251
rect 2329 10217 2363 10251
rect 2363 10217 2372 10251
rect 2320 10208 2372 10217
rect 2964 10251 3016 10260
rect 2964 10217 2973 10251
rect 2973 10217 3007 10251
rect 3007 10217 3016 10251
rect 2964 10208 3016 10217
rect 5908 10208 5960 10260
rect 7012 10208 7064 10260
rect 1768 10072 1820 10124
rect 2688 10072 2740 10124
rect 6920 10072 6972 10124
rect 15476 10208 15528 10260
rect 16764 10208 16816 10260
rect 20904 10251 20956 10260
rect 20904 10217 20913 10251
rect 20913 10217 20947 10251
rect 20947 10217 20956 10251
rect 20904 10208 20956 10217
rect 8852 10140 8904 10192
rect 10876 10140 10928 10192
rect 13912 10140 13964 10192
rect 9404 10072 9456 10124
rect 10508 10115 10560 10124
rect 10508 10081 10517 10115
rect 10517 10081 10551 10115
rect 10551 10081 10560 10115
rect 10508 10072 10560 10081
rect 10692 10115 10744 10124
rect 10692 10081 10701 10115
rect 10701 10081 10735 10115
rect 10735 10081 10744 10115
rect 10692 10072 10744 10081
rect 15752 10115 15804 10124
rect 15752 10081 15761 10115
rect 15761 10081 15795 10115
rect 15795 10081 15804 10115
rect 15752 10072 15804 10081
rect 21088 10115 21140 10124
rect 21088 10081 21097 10115
rect 21097 10081 21131 10115
rect 21131 10081 21140 10115
rect 21088 10072 21140 10081
rect 5448 10004 5500 10056
rect 3056 9911 3108 9920
rect 3056 9877 3065 9911
rect 3065 9877 3099 9911
rect 3099 9877 3108 9911
rect 3056 9868 3108 9877
rect 5540 9911 5592 9920
rect 5540 9877 5549 9911
rect 5549 9877 5583 9911
rect 5583 9877 5592 9911
rect 5540 9868 5592 9877
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 6644 9936 6696 9988
rect 7656 9936 7708 9988
rect 9588 10004 9640 10056
rect 12716 10004 12768 10056
rect 12808 9936 12860 9988
rect 7104 9868 7156 9920
rect 7564 9868 7616 9920
rect 9588 9911 9640 9920
rect 9588 9877 9597 9911
rect 9597 9877 9631 9911
rect 9631 9877 9640 9911
rect 9588 9868 9640 9877
rect 12900 9911 12952 9920
rect 12900 9877 12909 9911
rect 12909 9877 12943 9911
rect 12943 9877 12952 9911
rect 12900 9868 12952 9877
rect 4432 9766 4484 9818
rect 4496 9766 4548 9818
rect 4560 9766 4612 9818
rect 4624 9766 4676 9818
rect 11332 9766 11384 9818
rect 11396 9766 11448 9818
rect 11460 9766 11512 9818
rect 11524 9766 11576 9818
rect 18232 9766 18284 9818
rect 18296 9766 18348 9818
rect 18360 9766 18412 9818
rect 18424 9766 18476 9818
rect 6920 9664 6972 9716
rect 8852 9707 8904 9716
rect 8852 9673 8861 9707
rect 8861 9673 8895 9707
rect 8895 9673 8904 9707
rect 8852 9664 8904 9673
rect 3056 9528 3108 9580
rect 4160 9571 4212 9580
rect 4160 9537 4169 9571
rect 4169 9537 4203 9571
rect 4203 9537 4212 9571
rect 4160 9528 4212 9537
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 2044 9460 2096 9512
rect 5724 9460 5776 9512
rect 7656 9503 7708 9512
rect 2872 9392 2924 9444
rect 4068 9392 4120 9444
rect 4896 9392 4948 9444
rect 7656 9469 7665 9503
rect 7665 9469 7699 9503
rect 7699 9469 7708 9503
rect 7656 9460 7708 9469
rect 8668 9392 8720 9444
rect 9128 9460 9180 9512
rect 10508 9664 10560 9716
rect 15752 9664 15804 9716
rect 12532 9596 12584 9648
rect 9588 9528 9640 9580
rect 13820 9528 13872 9580
rect 15108 9571 15160 9580
rect 15108 9537 15117 9571
rect 15117 9537 15151 9571
rect 15151 9537 15160 9571
rect 15108 9528 15160 9537
rect 10692 9460 10744 9512
rect 10968 9460 11020 9512
rect 12716 9460 12768 9512
rect 9772 9392 9824 9444
rect 10416 9392 10468 9444
rect 15200 9392 15252 9444
rect 5264 9324 5316 9376
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 7288 9324 7340 9333
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 12440 9367 12492 9376
rect 12440 9333 12449 9367
rect 12449 9333 12483 9367
rect 12483 9333 12492 9367
rect 12440 9324 12492 9333
rect 12900 9367 12952 9376
rect 12900 9333 12909 9367
rect 12909 9333 12943 9367
rect 12943 9333 12952 9367
rect 12900 9324 12952 9333
rect 7882 9222 7934 9274
rect 7946 9222 7998 9274
rect 8010 9222 8062 9274
rect 8074 9222 8126 9274
rect 14782 9222 14834 9274
rect 14846 9222 14898 9274
rect 14910 9222 14962 9274
rect 14974 9222 15026 9274
rect 2044 9163 2096 9172
rect 2044 9129 2053 9163
rect 2053 9129 2087 9163
rect 2087 9129 2096 9163
rect 2044 9120 2096 9129
rect 7288 9120 7340 9172
rect 10324 9120 10376 9172
rect 12440 9120 12492 9172
rect 15752 9120 15804 9172
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 4160 8984 4212 9036
rect 5724 9052 5776 9104
rect 1676 8916 1728 8968
rect 4068 8916 4120 8968
rect 1492 8780 1544 8832
rect 3700 8848 3752 8900
rect 5540 8984 5592 9036
rect 6092 8984 6144 9036
rect 7564 9052 7616 9104
rect 9772 9052 9824 9104
rect 7104 9027 7156 9036
rect 7104 8993 7113 9027
rect 7113 8993 7147 9027
rect 7147 8993 7156 9027
rect 7104 8984 7156 8993
rect 9864 9027 9916 9036
rect 9864 8993 9873 9027
rect 9873 8993 9907 9027
rect 9907 8993 9916 9027
rect 9864 8984 9916 8993
rect 10232 8916 10284 8968
rect 10968 9052 11020 9104
rect 12900 8984 12952 9036
rect 16120 9027 16172 9036
rect 13268 8959 13320 8968
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 15108 8916 15160 8968
rect 16120 8993 16129 9027
rect 16129 8993 16163 9027
rect 16163 8993 16172 9027
rect 16120 8984 16172 8993
rect 21364 8984 21416 9036
rect 20628 8916 20680 8968
rect 9588 8848 9640 8900
rect 12716 8891 12768 8900
rect 5080 8780 5132 8832
rect 5264 8823 5316 8832
rect 5264 8789 5273 8823
rect 5273 8789 5307 8823
rect 5307 8789 5316 8823
rect 5264 8780 5316 8789
rect 7656 8823 7708 8832
rect 7656 8789 7665 8823
rect 7665 8789 7699 8823
rect 7699 8789 7708 8823
rect 7656 8780 7708 8789
rect 9496 8823 9548 8832
rect 9496 8789 9505 8823
rect 9505 8789 9539 8823
rect 9539 8789 9548 8823
rect 9496 8780 9548 8789
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 12716 8857 12725 8891
rect 12725 8857 12759 8891
rect 12759 8857 12768 8891
rect 12716 8848 12768 8857
rect 11888 8823 11940 8832
rect 11888 8789 11897 8823
rect 11897 8789 11931 8823
rect 11931 8789 11940 8823
rect 11888 8780 11940 8789
rect 20720 8823 20772 8832
rect 20720 8789 20729 8823
rect 20729 8789 20763 8823
rect 20763 8789 20772 8823
rect 20720 8780 20772 8789
rect 4432 8678 4484 8730
rect 4496 8678 4548 8730
rect 4560 8678 4612 8730
rect 4624 8678 4676 8730
rect 11332 8678 11384 8730
rect 11396 8678 11448 8730
rect 11460 8678 11512 8730
rect 11524 8678 11576 8730
rect 18232 8678 18284 8730
rect 18296 8678 18348 8730
rect 18360 8678 18412 8730
rect 18424 8678 18476 8730
rect 1676 8619 1728 8628
rect 1676 8585 1685 8619
rect 1685 8585 1719 8619
rect 1719 8585 1728 8619
rect 1676 8576 1728 8585
rect 4896 8619 4948 8628
rect 4896 8585 4905 8619
rect 4905 8585 4939 8619
rect 4939 8585 4948 8619
rect 4896 8576 4948 8585
rect 5080 8576 5132 8628
rect 5448 8576 5500 8628
rect 9588 8576 9640 8628
rect 9864 8619 9916 8628
rect 9864 8585 9873 8619
rect 9873 8585 9907 8619
rect 9907 8585 9916 8619
rect 9864 8576 9916 8585
rect 9772 8440 9824 8492
rect 13268 8483 13320 8492
rect 13268 8449 13277 8483
rect 13277 8449 13311 8483
rect 13311 8449 13320 8483
rect 13268 8440 13320 8449
rect 16120 8440 16172 8492
rect 20628 8576 20680 8628
rect 20720 8440 20772 8492
rect 1492 8415 1544 8424
rect 1492 8381 1501 8415
rect 1501 8381 1535 8415
rect 1535 8381 1544 8415
rect 1492 8372 1544 8381
rect 2044 8372 2096 8424
rect 2688 8415 2740 8424
rect 2688 8381 2697 8415
rect 2697 8381 2731 8415
rect 2731 8381 2740 8415
rect 2688 8372 2740 8381
rect 4068 8372 4120 8424
rect 5264 8372 5316 8424
rect 10876 8372 10928 8424
rect 12900 8372 12952 8424
rect 15476 8372 15528 8424
rect 2872 8304 2924 8356
rect 15108 8304 15160 8356
rect 20904 8415 20956 8424
rect 20904 8381 20913 8415
rect 20913 8381 20947 8415
rect 20947 8381 20956 8415
rect 20904 8372 20956 8381
rect 2964 8236 3016 8288
rect 10968 8279 11020 8288
rect 10968 8245 10977 8279
rect 10977 8245 11011 8279
rect 11011 8245 11020 8279
rect 10968 8236 11020 8245
rect 11060 8279 11112 8288
rect 11060 8245 11069 8279
rect 11069 8245 11103 8279
rect 11103 8245 11112 8279
rect 12624 8279 12676 8288
rect 11060 8236 11112 8245
rect 12624 8245 12633 8279
rect 12633 8245 12667 8279
rect 12667 8245 12676 8279
rect 12624 8236 12676 8245
rect 12992 8279 13044 8288
rect 12992 8245 13001 8279
rect 13001 8245 13035 8279
rect 13035 8245 13044 8279
rect 12992 8236 13044 8245
rect 16120 8304 16172 8356
rect 7882 8134 7934 8186
rect 7946 8134 7998 8186
rect 8010 8134 8062 8186
rect 8074 8134 8126 8186
rect 14782 8134 14834 8186
rect 14846 8134 14898 8186
rect 14910 8134 14962 8186
rect 14974 8134 15026 8186
rect 6092 8075 6144 8084
rect 6092 8041 6101 8075
rect 6101 8041 6135 8075
rect 6135 8041 6144 8075
rect 6092 8032 6144 8041
rect 9680 8032 9732 8084
rect 10876 8032 10928 8084
rect 12992 8075 13044 8084
rect 11152 7964 11204 8016
rect 7104 7896 7156 7948
rect 10232 7896 10284 7948
rect 10876 7896 10928 7948
rect 11888 7896 11940 7948
rect 12992 8041 13001 8075
rect 13001 8041 13035 8075
rect 13035 8041 13044 8075
rect 12992 8032 13044 8041
rect 15108 8032 15160 8084
rect 15476 8075 15528 8084
rect 15476 8041 15485 8075
rect 15485 8041 15519 8075
rect 15519 8041 15528 8075
rect 15476 8032 15528 8041
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 20904 8075 20956 8084
rect 20904 8041 20913 8075
rect 20913 8041 20947 8075
rect 20947 8041 20956 8075
rect 20904 8032 20956 8041
rect 13728 7896 13780 7948
rect 17960 7896 18012 7948
rect 21088 7939 21140 7948
rect 21088 7905 21097 7939
rect 21097 7905 21131 7939
rect 21131 7905 21140 7939
rect 21088 7896 21140 7905
rect 9772 7871 9824 7880
rect 9772 7837 9781 7871
rect 9781 7837 9815 7871
rect 9815 7837 9824 7871
rect 9772 7828 9824 7837
rect 12900 7828 12952 7880
rect 10324 7692 10376 7744
rect 11796 7735 11848 7744
rect 11796 7701 11805 7735
rect 11805 7701 11839 7735
rect 11839 7701 11848 7735
rect 11796 7692 11848 7701
rect 4432 7590 4484 7642
rect 4496 7590 4548 7642
rect 4560 7590 4612 7642
rect 4624 7590 4676 7642
rect 11332 7590 11384 7642
rect 11396 7590 11448 7642
rect 11460 7590 11512 7642
rect 11524 7590 11576 7642
rect 18232 7590 18284 7642
rect 18296 7590 18348 7642
rect 18360 7590 18412 7642
rect 18424 7590 18476 7642
rect 11796 7488 11848 7540
rect 13728 7531 13780 7540
rect 13728 7497 13737 7531
rect 13737 7497 13771 7531
rect 13771 7497 13780 7531
rect 13728 7488 13780 7497
rect 11060 7463 11112 7472
rect 11060 7429 11069 7463
rect 11069 7429 11103 7463
rect 11103 7429 11112 7463
rect 11060 7420 11112 7429
rect 10324 7352 10376 7404
rect 2964 7327 3016 7336
rect 2964 7293 2973 7327
rect 2973 7293 3007 7327
rect 3007 7293 3016 7327
rect 2964 7284 3016 7293
rect 4712 7284 4764 7336
rect 5448 7284 5500 7336
rect 5724 7327 5776 7336
rect 5724 7293 5733 7327
rect 5733 7293 5767 7327
rect 5767 7293 5776 7327
rect 5724 7284 5776 7293
rect 10876 7284 10928 7336
rect 11888 7352 11940 7404
rect 14096 7395 14148 7404
rect 14096 7361 14105 7395
rect 14105 7361 14139 7395
rect 14139 7361 14148 7395
rect 14096 7352 14148 7361
rect 13728 7327 13780 7336
rect 13728 7293 13737 7327
rect 13737 7293 13771 7327
rect 13771 7293 13780 7327
rect 13728 7284 13780 7293
rect 17776 7284 17828 7336
rect 2780 7148 2832 7200
rect 4804 7191 4856 7200
rect 4804 7157 4813 7191
rect 4813 7157 4847 7191
rect 4847 7157 4856 7191
rect 4804 7148 4856 7157
rect 10968 7216 11020 7268
rect 11152 7148 11204 7200
rect 12992 7216 13044 7268
rect 17500 7259 17552 7268
rect 17500 7225 17509 7259
rect 17509 7225 17543 7259
rect 17543 7225 17552 7259
rect 17500 7216 17552 7225
rect 7882 7046 7934 7098
rect 7946 7046 7998 7098
rect 8010 7046 8062 7098
rect 8074 7046 8126 7098
rect 14782 7046 14834 7098
rect 14846 7046 14898 7098
rect 14910 7046 14962 7098
rect 14974 7046 15026 7098
rect 7196 6944 7248 6996
rect 10876 6987 10928 6996
rect 10876 6953 10885 6987
rect 10885 6953 10919 6987
rect 10919 6953 10928 6987
rect 10876 6944 10928 6953
rect 11704 6944 11756 6996
rect 13176 6987 13228 6996
rect 13176 6953 13185 6987
rect 13185 6953 13219 6987
rect 13219 6953 13228 6987
rect 13176 6944 13228 6953
rect 2504 6808 2556 6860
rect 2596 6851 2648 6860
rect 2596 6817 2605 6851
rect 2605 6817 2639 6851
rect 2639 6817 2648 6851
rect 2596 6808 2648 6817
rect 6920 6808 6972 6860
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 4896 6783 4948 6792
rect 4896 6749 4905 6783
rect 4905 6749 4939 6783
rect 4939 6749 4948 6783
rect 4896 6740 4948 6749
rect 10232 6740 10284 6792
rect 12900 6876 12952 6928
rect 12992 6876 13044 6928
rect 19708 6808 19760 6860
rect 1768 6715 1820 6724
rect 1768 6681 1777 6715
rect 1777 6681 1811 6715
rect 1811 6681 1820 6715
rect 1768 6672 1820 6681
rect 2412 6715 2464 6724
rect 2412 6681 2421 6715
rect 2421 6681 2455 6715
rect 2455 6681 2464 6715
rect 2412 6672 2464 6681
rect 12716 6672 12768 6724
rect 20628 6740 20680 6792
rect 21180 6672 21232 6724
rect 11980 6604 12032 6656
rect 12256 6604 12308 6656
rect 4432 6502 4484 6554
rect 4496 6502 4548 6554
rect 4560 6502 4612 6554
rect 4624 6502 4676 6554
rect 11332 6502 11384 6554
rect 11396 6502 11448 6554
rect 11460 6502 11512 6554
rect 11524 6502 11576 6554
rect 18232 6502 18284 6554
rect 18296 6502 18348 6554
rect 18360 6502 18412 6554
rect 18424 6502 18476 6554
rect 2504 6400 2556 6452
rect 13176 6443 13228 6452
rect 2780 6264 2832 6316
rect 13176 6409 13185 6443
rect 13185 6409 13219 6443
rect 13219 6409 13228 6443
rect 13176 6400 13228 6409
rect 13728 6443 13780 6452
rect 13728 6409 13737 6443
rect 13737 6409 13771 6443
rect 13771 6409 13780 6443
rect 13728 6400 13780 6409
rect 19708 6443 19760 6452
rect 19708 6409 19717 6443
rect 19717 6409 19751 6443
rect 19751 6409 19760 6443
rect 19708 6400 19760 6409
rect 20628 6400 20680 6452
rect 4436 6239 4488 6248
rect 4436 6205 4445 6239
rect 4445 6205 4479 6239
rect 4479 6205 4488 6239
rect 4436 6196 4488 6205
rect 10232 6307 10284 6316
rect 10232 6273 10241 6307
rect 10241 6273 10275 6307
rect 10275 6273 10284 6307
rect 10232 6264 10284 6273
rect 12716 6264 12768 6316
rect 10416 6196 10468 6248
rect 2596 6128 2648 6180
rect 4068 6128 4120 6180
rect 5724 6128 5776 6180
rect 8208 6128 8260 6180
rect 12256 6196 12308 6248
rect 16212 6264 16264 6316
rect 18052 6264 18104 6316
rect 19708 6264 19760 6316
rect 13268 6196 13320 6248
rect 16120 6239 16172 6248
rect 4436 6060 4488 6112
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7288 6060 7340 6069
rect 8668 6060 8720 6112
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 12992 6128 13044 6180
rect 16120 6205 16129 6239
rect 16129 6205 16163 6239
rect 16163 6205 16172 6239
rect 16120 6196 16172 6205
rect 16488 6196 16540 6248
rect 20996 6196 21048 6248
rect 16580 6128 16632 6180
rect 17500 6128 17552 6180
rect 18604 6128 18656 6180
rect 10048 6060 10100 6069
rect 14648 6103 14700 6112
rect 14648 6069 14657 6103
rect 14657 6069 14691 6103
rect 14691 6069 14700 6103
rect 14648 6060 14700 6069
rect 7882 5958 7934 6010
rect 7946 5958 7998 6010
rect 8010 5958 8062 6010
rect 8074 5958 8126 6010
rect 14782 5958 14834 6010
rect 14846 5958 14898 6010
rect 14910 5958 14962 6010
rect 14974 5958 15026 6010
rect 9680 5856 9732 5908
rect 10416 5899 10468 5908
rect 7104 5788 7156 5840
rect 8208 5788 8260 5840
rect 1584 5763 1636 5772
rect 1584 5729 1593 5763
rect 1593 5729 1627 5763
rect 1627 5729 1636 5763
rect 1584 5720 1636 5729
rect 5724 5720 5776 5772
rect 6644 5763 6696 5772
rect 6644 5729 6653 5763
rect 6653 5729 6687 5763
rect 6687 5729 6696 5763
rect 6644 5720 6696 5729
rect 7288 5720 7340 5772
rect 8668 5720 8720 5772
rect 9496 5763 9548 5772
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 9496 5720 9548 5729
rect 10416 5865 10425 5899
rect 10425 5865 10459 5899
rect 10459 5865 10468 5899
rect 10416 5856 10468 5865
rect 14648 5856 14700 5908
rect 18052 5856 18104 5908
rect 10048 5788 10100 5840
rect 12624 5720 12676 5772
rect 18052 5720 18104 5772
rect 20904 5763 20956 5772
rect 20904 5729 20913 5763
rect 20913 5729 20947 5763
rect 20947 5729 20956 5763
rect 20904 5720 20956 5729
rect 4436 5652 4488 5704
rect 9864 5627 9916 5636
rect 9864 5593 9873 5627
rect 9873 5593 9907 5627
rect 9907 5593 9916 5627
rect 9864 5584 9916 5593
rect 12532 5652 12584 5704
rect 15660 5652 15712 5704
rect 15752 5652 15804 5704
rect 16488 5652 16540 5704
rect 17868 5695 17920 5704
rect 16396 5584 16448 5636
rect 17868 5661 17877 5695
rect 17877 5661 17911 5695
rect 17911 5661 17920 5695
rect 17868 5652 17920 5661
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 12256 5559 12308 5568
rect 12256 5525 12265 5559
rect 12265 5525 12299 5559
rect 12299 5525 12308 5559
rect 12256 5516 12308 5525
rect 4432 5414 4484 5466
rect 4496 5414 4548 5466
rect 4560 5414 4612 5466
rect 4624 5414 4676 5466
rect 11332 5414 11384 5466
rect 11396 5414 11448 5466
rect 11460 5414 11512 5466
rect 11524 5414 11576 5466
rect 18232 5414 18284 5466
rect 18296 5414 18348 5466
rect 18360 5414 18412 5466
rect 18424 5414 18476 5466
rect 1584 5312 1636 5364
rect 5724 5312 5776 5364
rect 6920 5355 6972 5364
rect 6920 5321 6929 5355
rect 6929 5321 6963 5355
rect 6963 5321 6972 5355
rect 6920 5312 6972 5321
rect 9680 5312 9732 5364
rect 9864 5312 9916 5364
rect 15752 5312 15804 5364
rect 18052 5312 18104 5364
rect 2504 5151 2556 5160
rect 2504 5117 2513 5151
rect 2513 5117 2547 5151
rect 2547 5117 2556 5151
rect 2504 5108 2556 5117
rect 9496 5176 9548 5228
rect 12624 5176 12676 5228
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 19708 5312 19760 5364
rect 20904 5355 20956 5364
rect 19248 5176 19300 5228
rect 20904 5321 20913 5355
rect 20913 5321 20947 5355
rect 20947 5321 20956 5355
rect 20904 5312 20956 5321
rect 7104 5151 7156 5160
rect 4068 5040 4120 5092
rect 7104 5117 7113 5151
rect 7113 5117 7147 5151
rect 7147 5117 7156 5151
rect 7104 5108 7156 5117
rect 2688 4972 2740 5024
rect 6000 5040 6052 5092
rect 8668 5040 8720 5092
rect 12532 5108 12584 5160
rect 15844 5151 15896 5160
rect 15844 5117 15853 5151
rect 15853 5117 15887 5151
rect 15887 5117 15896 5151
rect 15844 5108 15896 5117
rect 16120 5108 16172 5160
rect 16672 5108 16724 5160
rect 21088 5151 21140 5160
rect 16580 5040 16632 5092
rect 21088 5117 21097 5151
rect 21097 5117 21131 5151
rect 21131 5117 21140 5151
rect 21088 5108 21140 5117
rect 18144 5040 18196 5092
rect 18604 5040 18656 5092
rect 12256 4972 12308 5024
rect 17408 5015 17460 5024
rect 17408 4981 17417 5015
rect 17417 4981 17451 5015
rect 17451 4981 17460 5015
rect 17408 4972 17460 4981
rect 7882 4870 7934 4922
rect 7946 4870 7998 4922
rect 8010 4870 8062 4922
rect 8074 4870 8126 4922
rect 14782 4870 14834 4922
rect 14846 4870 14898 4922
rect 14910 4870 14962 4922
rect 14974 4870 15026 4922
rect 4068 4768 4120 4820
rect 6644 4811 6696 4820
rect 6644 4777 6653 4811
rect 6653 4777 6687 4811
rect 6687 4777 6696 4811
rect 6644 4768 6696 4777
rect 10692 4768 10744 4820
rect 11152 4768 11204 4820
rect 16396 4811 16448 4820
rect 16396 4777 16405 4811
rect 16405 4777 16439 4811
rect 16439 4777 16448 4811
rect 16396 4768 16448 4777
rect 6000 4632 6052 4684
rect 12532 4675 12584 4684
rect 12532 4641 12541 4675
rect 12541 4641 12575 4675
rect 12575 4641 12584 4675
rect 12532 4632 12584 4641
rect 13268 4675 13320 4684
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 13268 4632 13320 4641
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 10416 4607 10468 4616
rect 10416 4573 10425 4607
rect 10425 4573 10459 4607
rect 10459 4573 10468 4607
rect 10416 4564 10468 4573
rect 10784 4496 10836 4548
rect 11704 4539 11756 4548
rect 11704 4505 11713 4539
rect 11713 4505 11747 4539
rect 11747 4505 11756 4539
rect 11704 4496 11756 4505
rect 16212 4607 16264 4616
rect 16212 4573 16221 4607
rect 16221 4573 16255 4607
rect 16255 4573 16264 4607
rect 16212 4564 16264 4573
rect 17868 4700 17920 4752
rect 16672 4675 16724 4684
rect 16672 4641 16681 4675
rect 16681 4641 16715 4675
rect 16715 4641 16724 4675
rect 17224 4675 17276 4684
rect 16672 4632 16724 4641
rect 17224 4641 17233 4675
rect 17233 4641 17267 4675
rect 17267 4641 17276 4675
rect 17224 4632 17276 4641
rect 17408 4675 17460 4684
rect 17408 4641 17417 4675
rect 17417 4641 17451 4675
rect 17451 4641 17460 4675
rect 17408 4632 17460 4641
rect 18144 4632 18196 4684
rect 15844 4496 15896 4548
rect 4432 4326 4484 4378
rect 4496 4326 4548 4378
rect 4560 4326 4612 4378
rect 4624 4326 4676 4378
rect 11332 4326 11384 4378
rect 11396 4326 11448 4378
rect 11460 4326 11512 4378
rect 11524 4326 11576 4378
rect 18232 4326 18284 4378
rect 18296 4326 18348 4378
rect 18360 4326 18412 4378
rect 18424 4326 18476 4378
rect 11704 4224 11756 4276
rect 13268 4267 13320 4276
rect 13268 4233 13277 4267
rect 13277 4233 13311 4267
rect 13311 4233 13320 4267
rect 13268 4224 13320 4233
rect 15844 4224 15896 4276
rect 14096 4088 14148 4140
rect 2780 4020 2832 4072
rect 2872 4020 2924 4072
rect 7656 4020 7708 4072
rect 11152 4020 11204 4072
rect 12256 4063 12308 4072
rect 12256 4029 12265 4063
rect 12265 4029 12299 4063
rect 12299 4029 12308 4063
rect 12256 4020 12308 4029
rect 13636 4063 13688 4072
rect 13636 4029 13645 4063
rect 13645 4029 13679 4063
rect 13679 4029 13688 4063
rect 13636 4020 13688 4029
rect 15476 4020 15528 4072
rect 16212 4063 16264 4072
rect 16212 4029 16221 4063
rect 16221 4029 16255 4063
rect 16255 4029 16264 4063
rect 16212 4020 16264 4029
rect 19248 4020 19300 4072
rect 8668 3995 8720 4004
rect 8668 3961 8677 3995
rect 8677 3961 8711 3995
rect 8711 3961 8720 3995
rect 8668 3952 8720 3961
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 13912 3952 13964 4004
rect 10508 3884 10560 3936
rect 14188 3927 14240 3936
rect 14188 3893 14197 3927
rect 14197 3893 14231 3927
rect 14231 3893 14240 3927
rect 14188 3884 14240 3893
rect 20904 3884 20956 3936
rect 7882 3782 7934 3834
rect 7946 3782 7998 3834
rect 8010 3782 8062 3834
rect 8074 3782 8126 3834
rect 14782 3782 14834 3834
rect 14846 3782 14898 3834
rect 14910 3782 14962 3834
rect 14974 3782 15026 3834
rect 13268 3680 13320 3732
rect 15108 3723 15160 3732
rect 15108 3689 15117 3723
rect 15117 3689 15151 3723
rect 15151 3689 15160 3723
rect 15108 3680 15160 3689
rect 20996 3680 21048 3732
rect 6000 3655 6052 3664
rect 6000 3621 6009 3655
rect 6009 3621 6043 3655
rect 6043 3621 6052 3655
rect 6000 3612 6052 3621
rect 8668 3612 8720 3664
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 6920 3544 6972 3596
rect 7656 3587 7708 3596
rect 7656 3553 7665 3587
rect 7665 3553 7699 3587
rect 7699 3553 7708 3587
rect 7656 3544 7708 3553
rect 8576 3587 8628 3596
rect 8576 3553 8585 3587
rect 8585 3553 8619 3587
rect 8619 3553 8628 3587
rect 8576 3544 8628 3553
rect 10508 3587 10560 3596
rect 10508 3553 10517 3587
rect 10517 3553 10551 3587
rect 10551 3553 10560 3587
rect 10508 3544 10560 3553
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 12072 3544 12124 3596
rect 14188 3544 14240 3596
rect 20720 3544 20772 3596
rect 22100 3544 22152 3596
rect 13636 3476 13688 3528
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 2504 3340 2556 3392
rect 9312 3340 9364 3392
rect 9588 3340 9640 3392
rect 10692 3340 10744 3392
rect 4432 3238 4484 3290
rect 4496 3238 4548 3290
rect 4560 3238 4612 3290
rect 4624 3238 4676 3290
rect 11332 3238 11384 3290
rect 11396 3238 11448 3290
rect 11460 3238 11512 3290
rect 11524 3238 11576 3290
rect 18232 3238 18284 3290
rect 18296 3238 18348 3290
rect 18360 3238 18412 3290
rect 18424 3238 18476 3290
rect 1952 3136 2004 3188
rect 4896 3136 4948 3188
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 8576 3136 8628 3188
rect 9312 3179 9364 3188
rect 2320 2932 2372 2984
rect 2504 2975 2556 2984
rect 2504 2941 2513 2975
rect 2513 2941 2547 2975
rect 2547 2941 2556 2975
rect 2504 2932 2556 2941
rect 4436 2975 4488 2984
rect 4436 2941 4445 2975
rect 4445 2941 4479 2975
rect 4479 2941 4488 2975
rect 4436 2932 4488 2941
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 6828 2932 6880 2941
rect 9312 3145 9321 3179
rect 9321 3145 9355 3179
rect 9355 3145 9364 3179
rect 9312 3136 9364 3145
rect 9588 3000 9640 3052
rect 9864 3068 9916 3120
rect 10692 3043 10744 3052
rect 10692 3009 10701 3043
rect 10701 3009 10735 3043
rect 10735 3009 10744 3043
rect 10692 3000 10744 3009
rect 10784 3000 10836 3052
rect 15384 3136 15436 3188
rect 17960 3136 18012 3188
rect 20720 3179 20772 3188
rect 20720 3145 20729 3179
rect 20729 3145 20763 3179
rect 20763 3145 20772 3179
rect 20720 3136 20772 3145
rect 13912 3111 13964 3120
rect 13912 3077 13921 3111
rect 13921 3077 13955 3111
rect 13955 3077 13964 3111
rect 13912 3068 13964 3077
rect 17224 3068 17276 3120
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 10600 2975 10652 2984
rect 10600 2941 10609 2975
rect 10609 2941 10643 2975
rect 10643 2941 10652 2975
rect 10600 2932 10652 2941
rect 9772 2864 9824 2916
rect 12808 2864 12860 2916
rect 13360 2864 13412 2916
rect 16120 2975 16172 2984
rect 16120 2941 16129 2975
rect 16129 2941 16163 2975
rect 16163 2941 16172 2975
rect 16120 2932 16172 2941
rect 18236 2975 18288 2984
rect 18236 2941 18245 2975
rect 18245 2941 18279 2975
rect 18279 2941 18288 2975
rect 18236 2932 18288 2941
rect 20076 2975 20128 2984
rect 20076 2941 20085 2975
rect 20085 2941 20119 2975
rect 20119 2941 20128 2975
rect 20076 2932 20128 2941
rect 14096 2907 14148 2916
rect 14096 2873 14105 2907
rect 14105 2873 14139 2907
rect 14139 2873 14148 2907
rect 14096 2864 14148 2873
rect 17500 2907 17552 2916
rect 17500 2873 17509 2907
rect 17509 2873 17543 2907
rect 17543 2873 17552 2907
rect 17500 2864 17552 2873
rect 13268 2839 13320 2848
rect 13268 2805 13277 2839
rect 13277 2805 13311 2839
rect 13311 2805 13320 2839
rect 13268 2796 13320 2805
rect 7882 2694 7934 2746
rect 7946 2694 7998 2746
rect 8010 2694 8062 2746
rect 8074 2694 8126 2746
rect 14782 2694 14834 2746
rect 14846 2694 14898 2746
rect 14910 2694 14962 2746
rect 14974 2694 15026 2746
rect 2320 2592 2372 2644
rect 4436 2635 4488 2644
rect 4436 2601 4445 2635
rect 4445 2601 4479 2635
rect 4479 2601 4488 2635
rect 4436 2592 4488 2601
rect 6828 2592 6880 2644
rect 6920 2635 6972 2644
rect 6920 2601 6929 2635
rect 6929 2601 6963 2635
rect 6963 2601 6972 2635
rect 6920 2592 6972 2601
rect 10416 2592 10468 2644
rect 1860 2524 1912 2576
rect 480 2456 532 2508
rect 3700 2456 3752 2508
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 6920 2456 6972 2508
rect 8760 2524 8812 2576
rect 13912 2592 13964 2644
rect 16120 2635 16172 2644
rect 16120 2601 16129 2635
rect 16129 2601 16163 2635
rect 16163 2601 16172 2635
rect 16120 2592 16172 2601
rect 17500 2592 17552 2644
rect 18236 2592 18288 2644
rect 15476 2567 15528 2576
rect 15476 2533 15485 2567
rect 15485 2533 15519 2567
rect 15519 2533 15528 2567
rect 15476 2524 15528 2533
rect 20904 2567 20956 2576
rect 20904 2533 20913 2567
rect 20913 2533 20947 2567
rect 20947 2533 20956 2567
rect 20904 2524 20956 2533
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 10600 2456 10652 2508
rect 13268 2456 13320 2508
rect 14096 2456 14148 2508
rect 15660 2456 15712 2508
rect 17040 2456 17092 2508
rect 18880 2456 18932 2508
rect 13728 2388 13780 2440
rect 20720 2363 20772 2372
rect 20720 2329 20729 2363
rect 20729 2329 20763 2363
rect 20763 2329 20772 2363
rect 20720 2320 20772 2329
rect 13360 2252 13412 2304
rect 4432 2150 4484 2202
rect 4496 2150 4548 2202
rect 4560 2150 4612 2202
rect 4624 2150 4676 2202
rect 11332 2150 11384 2202
rect 11396 2150 11448 2202
rect 11460 2150 11512 2202
rect 11524 2150 11576 2202
rect 18232 2150 18284 2202
rect 18296 2150 18348 2202
rect 18360 2150 18412 2202
rect 18424 2150 18476 2202
<< metal2 >>
rect 938 24323 994 25123
rect 2778 24323 2834 25123
rect 4618 24323 4674 25123
rect 5998 24323 6054 25123
rect 7838 24323 7894 25123
rect 9678 24323 9734 25123
rect 11518 24323 11574 25123
rect 12898 24323 12954 25123
rect 14738 24323 14794 25123
rect 16578 24323 16634 25123
rect 17958 24323 18014 25123
rect 19798 24323 19854 25123
rect 21638 24323 21694 25123
rect 952 22574 980 24323
rect 1490 23216 1546 23225
rect 1490 23151 1546 23160
rect 1504 22778 1532 23151
rect 1492 22772 1544 22778
rect 1492 22714 1544 22720
rect 2792 22574 2820 24323
rect 4632 23066 4660 24323
rect 4632 23038 4844 23066
rect 4406 22876 4702 22896
rect 4462 22874 4486 22876
rect 4542 22874 4566 22876
rect 4622 22874 4646 22876
rect 4484 22822 4486 22874
rect 4548 22822 4560 22874
rect 4622 22822 4624 22874
rect 4462 22820 4486 22822
rect 4542 22820 4566 22822
rect 4622 22820 4646 22822
rect 4406 22800 4702 22820
rect 4816 22574 4844 23038
rect 6012 22574 6040 24323
rect 7852 22574 7880 24323
rect 9692 22574 9720 24323
rect 11532 23066 11560 24323
rect 11532 23038 11744 23066
rect 11306 22876 11602 22896
rect 11362 22874 11386 22876
rect 11442 22874 11466 22876
rect 11522 22874 11546 22876
rect 11384 22822 11386 22874
rect 11448 22822 11460 22874
rect 11522 22822 11524 22874
rect 11362 22820 11386 22822
rect 11442 22820 11466 22822
rect 11522 22820 11546 22822
rect 11306 22800 11602 22820
rect 940 22568 992 22574
rect 940 22510 992 22516
rect 2780 22568 2832 22574
rect 2780 22510 2832 22516
rect 4804 22568 4856 22574
rect 4804 22510 4856 22516
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 7840 22568 7892 22574
rect 7840 22510 7892 22516
rect 9680 22568 9732 22574
rect 9680 22510 9732 22516
rect 11716 22506 11744 23038
rect 12912 22574 12940 24323
rect 14752 22574 14780 24323
rect 16592 22574 16620 24323
rect 17972 22574 18000 24323
rect 18206 22876 18502 22896
rect 18262 22874 18286 22876
rect 18342 22874 18366 22876
rect 18422 22874 18446 22876
rect 18284 22822 18286 22874
rect 18348 22822 18360 22874
rect 18422 22822 18424 22874
rect 18262 22820 18286 22822
rect 18342 22820 18366 22822
rect 18422 22820 18446 22822
rect 18206 22800 18502 22820
rect 19812 22574 19840 24323
rect 21086 23216 21142 23225
rect 21086 23151 21142 23160
rect 21100 22574 21128 23151
rect 12900 22568 12952 22574
rect 12900 22510 12952 22516
rect 14740 22568 14792 22574
rect 14740 22510 14792 22516
rect 16580 22568 16632 22574
rect 16580 22510 16632 22516
rect 17960 22568 18012 22574
rect 17960 22510 18012 22516
rect 19800 22568 19852 22574
rect 19800 22510 19852 22516
rect 21088 22568 21140 22574
rect 21088 22510 21140 22516
rect 1584 22500 1636 22506
rect 1584 22442 1636 22448
rect 11704 22500 11756 22506
rect 11704 22442 11756 22448
rect 1596 21690 1624 22442
rect 1676 22432 1728 22438
rect 1676 22374 1728 22380
rect 3424 22432 3476 22438
rect 3424 22374 3476 22380
rect 5080 22432 5132 22438
rect 5080 22374 5132 22380
rect 5724 22432 5776 22438
rect 5724 22374 5776 22380
rect 8208 22432 8260 22438
rect 8208 22374 8260 22380
rect 9680 22432 9732 22438
rect 9680 22374 9732 22380
rect 10324 22432 10376 22438
rect 10324 22374 10376 22380
rect 13084 22432 13136 22438
rect 13084 22374 13136 22380
rect 15384 22432 15436 22438
rect 15384 22374 15436 22380
rect 16028 22432 16080 22438
rect 16028 22374 16080 22380
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 20168 22432 20220 22438
rect 20168 22374 20220 22380
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1398 20496 1454 20505
rect 1398 20431 1454 20440
rect 1412 20398 1440 20431
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1398 17776 1454 17785
rect 1398 17711 1400 17720
rect 1452 17711 1454 17720
rect 1400 17682 1452 17688
rect 1688 16658 1716 22374
rect 3240 21616 3292 21622
rect 3240 21558 3292 21564
rect 3252 20466 3280 21558
rect 3436 21486 3464 22374
rect 4406 21788 4702 21808
rect 4462 21786 4486 21788
rect 4542 21786 4566 21788
rect 4622 21786 4646 21788
rect 4484 21734 4486 21786
rect 4548 21734 4560 21786
rect 4622 21734 4624 21786
rect 4462 21732 4486 21734
rect 4542 21732 4566 21734
rect 4622 21732 4646 21734
rect 4406 21712 4702 21732
rect 5092 21486 5120 22374
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 5184 21622 5212 21966
rect 5172 21616 5224 21622
rect 5172 21558 5224 21564
rect 5736 21486 5764 22374
rect 7856 22332 8152 22352
rect 7912 22330 7936 22332
rect 7992 22330 8016 22332
rect 8072 22330 8096 22332
rect 7934 22278 7936 22330
rect 7998 22278 8010 22330
rect 8072 22278 8074 22330
rect 7912 22276 7936 22278
rect 7992 22276 8016 22278
rect 8072 22276 8096 22278
rect 7856 22256 8152 22276
rect 6828 22160 6880 22166
rect 6828 22102 6880 22108
rect 5816 22024 5868 22030
rect 5816 21966 5868 21972
rect 3424 21480 3476 21486
rect 3424 21422 3476 21428
rect 5080 21480 5132 21486
rect 5080 21422 5132 21428
rect 5724 21480 5776 21486
rect 5724 21422 5776 21428
rect 5356 21412 5408 21418
rect 5356 21354 5408 21360
rect 3700 21344 3752 21350
rect 3700 21286 3752 21292
rect 3240 20460 3292 20466
rect 3240 20402 3292 20408
rect 3516 20324 3568 20330
rect 3516 20266 3568 20272
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 2424 19310 2452 20198
rect 3528 20058 3556 20266
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 2412 19304 2464 19310
rect 2412 19246 2464 19252
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 2320 17536 2372 17542
rect 2320 17478 2372 17484
rect 2332 16658 2360 17478
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 2320 16652 2372 16658
rect 2320 16594 2372 16600
rect 2136 16040 2188 16046
rect 2136 15982 2188 15988
rect 1398 15736 1454 15745
rect 1398 15671 1454 15680
rect 1412 15570 1440 15671
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 1872 14958 1900 15302
rect 1860 14952 1912 14958
rect 1860 14894 1912 14900
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1964 14074 1992 14350
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 1964 13394 1992 14010
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1490 13016 1546 13025
rect 1490 12951 1492 12960
rect 1544 12951 1546 12960
rect 1492 12922 1544 12928
rect 2056 11762 2084 14758
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 1490 10296 1546 10305
rect 1490 10231 1492 10240
rect 1544 10231 1546 10240
rect 1492 10202 1544 10208
rect 1768 10124 1820 10130
rect 1768 10066 1820 10072
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1412 8265 1440 8978
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1504 8430 1532 8774
rect 1688 8634 1716 8910
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1492 8424 1544 8430
rect 1492 8366 1544 8372
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1780 6730 1808 10066
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 2056 9178 2084 9454
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2056 8430 2084 9114
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 2148 6914 2176 15982
rect 2320 14816 2372 14822
rect 2320 14758 2372 14764
rect 2332 14482 2360 14758
rect 2320 14476 2372 14482
rect 2320 14418 2372 14424
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 2228 13864 2280 13870
rect 2228 13806 2280 13812
rect 2240 11830 2268 13806
rect 2332 13530 2360 14214
rect 2424 13938 2452 16730
rect 2608 16574 2636 19110
rect 2516 16546 2636 16574
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 2228 11824 2280 11830
rect 2228 11766 2280 11772
rect 2332 11218 2360 13466
rect 2412 12708 2464 12714
rect 2412 12650 2464 12656
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2332 10266 2360 10542
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 1964 6886 2176 6914
rect 1768 6724 1820 6730
rect 1768 6666 1820 6672
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1492 5568 1544 5574
rect 1490 5536 1492 5545
rect 1544 5536 1546 5545
rect 1490 5471 1546 5480
rect 1596 5370 1624 5714
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1412 2825 1440 3538
rect 1398 2816 1454 2825
rect 1398 2751 1454 2760
rect 1872 2582 1900 3878
rect 1964 3194 1992 6886
rect 2424 6730 2452 12650
rect 2516 8242 2544 16546
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 2792 13870 2820 14350
rect 3160 13938 3188 14350
rect 3528 14278 3556 14758
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2792 13530 2820 13806
rect 3528 13734 3556 14214
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 3332 13388 3384 13394
rect 3332 13330 3384 13336
rect 3344 12986 3372 13330
rect 3608 13184 3660 13190
rect 3608 13126 3660 13132
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3620 12850 3648 13126
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3160 11762 3188 12650
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2608 10674 2636 11494
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2700 10606 2728 10950
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2700 10130 2728 10542
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2976 10266 3004 10406
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2700 8430 2728 10066
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 3068 9586 3096 9862
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2884 8362 2912 9386
rect 3712 8906 3740 21286
rect 4406 20700 4702 20720
rect 4462 20698 4486 20700
rect 4542 20698 4566 20700
rect 4622 20698 4646 20700
rect 4484 20646 4486 20698
rect 4548 20646 4560 20698
rect 4622 20646 4624 20698
rect 4462 20644 4486 20646
rect 4542 20644 4566 20646
rect 4622 20644 4646 20646
rect 4406 20624 4702 20644
rect 4068 20460 4120 20466
rect 4068 20402 4120 20408
rect 4080 19360 4108 20402
rect 4252 20324 4304 20330
rect 4252 20266 4304 20272
rect 4264 19514 4292 20266
rect 4406 19612 4702 19632
rect 4462 19610 4486 19612
rect 4542 19610 4566 19612
rect 4622 19610 4646 19612
rect 4484 19558 4486 19610
rect 4548 19558 4560 19610
rect 4622 19558 4624 19610
rect 4462 19556 4486 19558
rect 4542 19556 4566 19558
rect 4622 19556 4646 19558
rect 4406 19536 4702 19556
rect 4252 19508 4304 19514
rect 4252 19450 4304 19456
rect 4080 19332 4200 19360
rect 4172 17746 4200 19332
rect 5368 19310 5396 21354
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 4896 19304 4948 19310
rect 4896 19246 4948 19252
rect 5356 19304 5408 19310
rect 5356 19246 5408 19252
rect 4406 18524 4702 18544
rect 4462 18522 4486 18524
rect 4542 18522 4566 18524
rect 4622 18522 4646 18524
rect 4484 18470 4486 18522
rect 4548 18470 4560 18522
rect 4622 18470 4624 18522
rect 4462 18468 4486 18470
rect 4542 18468 4566 18470
rect 4622 18468 4646 18470
rect 4406 18448 4702 18468
rect 4908 18222 4936 19246
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5368 18222 5396 18566
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 5356 18216 5408 18222
rect 5356 18158 5408 18164
rect 4620 18148 4672 18154
rect 4620 18090 4672 18096
rect 4632 17814 4660 18090
rect 4620 17808 4672 17814
rect 4620 17750 4672 17756
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4172 16114 4200 17682
rect 4406 17436 4702 17456
rect 4462 17434 4486 17436
rect 4542 17434 4566 17436
rect 4622 17434 4646 17436
rect 4484 17382 4486 17434
rect 4548 17382 4560 17434
rect 4622 17382 4624 17434
rect 4462 17380 4486 17382
rect 4542 17380 4566 17382
rect 4622 17380 4646 17382
rect 4406 17360 4702 17380
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 4264 13462 4292 16730
rect 4406 16348 4702 16368
rect 4462 16346 4486 16348
rect 4542 16346 4566 16348
rect 4622 16346 4646 16348
rect 4484 16294 4486 16346
rect 4548 16294 4560 16346
rect 4622 16294 4624 16346
rect 4462 16292 4486 16294
rect 4542 16292 4566 16294
rect 4622 16292 4646 16294
rect 4406 16272 4702 16292
rect 4344 15972 4396 15978
rect 4344 15914 4396 15920
rect 4356 15706 4384 15914
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4908 15570 4936 18158
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 5000 17814 5028 18022
rect 4988 17808 5040 17814
rect 4988 17750 5040 17756
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 5000 15706 5028 15846
rect 4988 15700 5040 15706
rect 4988 15642 5040 15648
rect 4896 15564 4948 15570
rect 4896 15506 4948 15512
rect 5264 15564 5316 15570
rect 5264 15506 5316 15512
rect 4406 15260 4702 15280
rect 4462 15258 4486 15260
rect 4542 15258 4566 15260
rect 4622 15258 4646 15260
rect 4484 15206 4486 15258
rect 4548 15206 4560 15258
rect 4622 15206 4624 15258
rect 4462 15204 4486 15206
rect 4542 15204 4566 15206
rect 4622 15204 4646 15206
rect 4406 15184 4702 15204
rect 4406 14172 4702 14192
rect 4462 14170 4486 14172
rect 4542 14170 4566 14172
rect 4622 14170 4646 14172
rect 4484 14118 4486 14170
rect 4548 14118 4560 14170
rect 4622 14118 4624 14170
rect 4462 14116 4486 14118
rect 4542 14116 4566 14118
rect 4622 14116 4646 14118
rect 4406 14096 4702 14116
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 4816 13326 4844 14010
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4406 13084 4702 13104
rect 4462 13082 4486 13084
rect 4542 13082 4566 13084
rect 4622 13082 4646 13084
rect 4484 13030 4486 13082
rect 4548 13030 4560 13082
rect 4622 13030 4624 13082
rect 4462 13028 4486 13030
rect 4542 13028 4566 13030
rect 4622 13028 4646 13030
rect 4406 13008 4702 13028
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4356 12442 4384 12718
rect 4344 12436 4396 12442
rect 4908 12434 4936 15506
rect 5276 15162 5304 15506
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5460 13734 5488 21286
rect 5828 21146 5856 21966
rect 6460 21888 6512 21894
rect 6460 21830 6512 21836
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5816 21140 5868 21146
rect 5816 21082 5868 21088
rect 5724 21072 5776 21078
rect 5724 21014 5776 21020
rect 5632 20392 5684 20398
rect 5632 20334 5684 20340
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 5552 19990 5580 20198
rect 5540 19984 5592 19990
rect 5540 19926 5592 19932
rect 5644 19854 5672 20334
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5552 18154 5580 19654
rect 5644 19310 5672 19790
rect 5736 19718 5764 21014
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5828 20058 5856 20946
rect 5816 20052 5868 20058
rect 5816 19994 5868 20000
rect 5724 19712 5776 19718
rect 5724 19654 5776 19660
rect 5632 19304 5684 19310
rect 5632 19246 5684 19252
rect 5540 18148 5592 18154
rect 5540 18090 5592 18096
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5644 15570 5672 15846
rect 5736 15638 5764 16050
rect 5724 15632 5776 15638
rect 5724 15574 5776 15580
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 5644 14550 5672 15506
rect 5736 15162 5764 15574
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5632 14544 5684 14550
rect 5632 14486 5684 14492
rect 5632 13796 5684 13802
rect 5632 13738 5684 13744
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5644 13326 5672 13738
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 4344 12378 4396 12384
rect 4816 12406 4936 12434
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4172 11830 4200 12242
rect 4406 11996 4702 12016
rect 4462 11994 4486 11996
rect 4542 11994 4566 11996
rect 4622 11994 4646 11996
rect 4484 11942 4486 11994
rect 4548 11942 4560 11994
rect 4622 11942 4624 11994
rect 4462 11940 4486 11942
rect 4542 11940 4566 11942
rect 4622 11940 4646 11942
rect 4406 11920 4702 11940
rect 4160 11824 4212 11830
rect 4160 11766 4212 11772
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3804 10810 3832 11698
rect 4172 11354 4200 11766
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4264 11218 4292 11494
rect 4356 11218 4384 11630
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4080 9450 4108 10542
rect 4172 9586 4200 11018
rect 4406 10908 4702 10928
rect 4462 10906 4486 10908
rect 4542 10906 4566 10908
rect 4622 10906 4646 10908
rect 4484 10854 4486 10906
rect 4548 10854 4560 10906
rect 4622 10854 4624 10906
rect 4462 10852 4486 10854
rect 4542 10852 4566 10854
rect 4622 10852 4646 10854
rect 4406 10832 4702 10852
rect 4406 9820 4702 9840
rect 4462 9818 4486 9820
rect 4542 9818 4566 9820
rect 4622 9818 4646 9820
rect 4484 9766 4486 9818
rect 4548 9766 4560 9818
rect 4622 9766 4624 9818
rect 4462 9764 4486 9766
rect 4542 9764 4566 9766
rect 4622 9764 4646 9766
rect 4406 9744 4702 9764
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 4080 8974 4108 9386
rect 4172 9042 4200 9522
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3700 8900 3752 8906
rect 3700 8842 3752 8848
rect 4080 8430 4108 8910
rect 4406 8732 4702 8752
rect 4462 8730 4486 8732
rect 4542 8730 4566 8732
rect 4622 8730 4646 8732
rect 4484 8678 4486 8730
rect 4548 8678 4560 8730
rect 4622 8678 4624 8730
rect 4462 8676 4486 8678
rect 4542 8676 4566 8678
rect 4622 8676 4646 8678
rect 4406 8656 4702 8676
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2516 8214 2728 8242
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 2516 6458 2544 6802
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2608 6186 2636 6802
rect 2596 6180 2648 6186
rect 2596 6122 2648 6128
rect 2504 5160 2556 5166
rect 2608 5148 2636 6122
rect 2556 5120 2636 5148
rect 2504 5102 2556 5108
rect 2700 5030 2728 8214
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2792 6322 2820 7142
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 2792 4078 2820 6258
rect 2884 4078 2912 8298
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 7342 3004 8230
rect 4406 7644 4702 7664
rect 4462 7642 4486 7644
rect 4542 7642 4566 7644
rect 4622 7642 4646 7644
rect 4484 7590 4486 7642
rect 4548 7590 4560 7642
rect 4622 7590 4624 7642
rect 4462 7588 4486 7590
rect 4542 7588 4566 7590
rect 4622 7588 4646 7590
rect 4406 7568 4702 7588
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4724 6798 4752 7278
rect 4816 7206 4844 12406
rect 5460 11150 5488 13262
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5460 10062 5488 11086
rect 5920 10266 5948 21286
rect 6472 21078 6500 21830
rect 6840 21690 6868 22102
rect 7012 22092 7064 22098
rect 7012 22034 7064 22040
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 7024 21486 7052 22034
rect 7012 21480 7064 21486
rect 7012 21422 7064 21428
rect 7856 21244 8152 21264
rect 7912 21242 7936 21244
rect 7992 21242 8016 21244
rect 8072 21242 8096 21244
rect 7934 21190 7936 21242
rect 7998 21190 8010 21242
rect 8072 21190 8074 21242
rect 7912 21188 7936 21190
rect 7992 21188 8016 21190
rect 8072 21188 8096 21190
rect 7856 21168 8152 21188
rect 6460 21072 6512 21078
rect 6460 21014 6512 21020
rect 6092 20868 6144 20874
rect 6092 20810 6144 20816
rect 6104 20466 6132 20810
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 6104 19514 6132 20402
rect 6184 19984 6236 19990
rect 6184 19926 6236 19932
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 6196 19310 6224 19926
rect 6368 19916 6420 19922
rect 6472 19904 6500 21014
rect 8220 21010 8248 22374
rect 9692 22098 9720 22374
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 6552 20936 6604 20942
rect 6552 20878 6604 20884
rect 6420 19876 6500 19904
rect 6368 19858 6420 19864
rect 6472 19310 6500 19876
rect 6564 19786 6592 20878
rect 6920 20528 6972 20534
rect 6920 20470 6972 20476
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 6552 19780 6604 19786
rect 6552 19722 6604 19728
rect 6184 19304 6236 19310
rect 6184 19246 6236 19252
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 6656 19242 6684 19858
rect 6644 19236 6696 19242
rect 6644 19178 6696 19184
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 6012 17882 6040 18770
rect 6656 18426 6684 19178
rect 6932 18834 6960 20470
rect 8404 20466 8432 21626
rect 8496 21418 8524 21830
rect 8484 21412 8536 21418
rect 8484 21354 8536 21360
rect 9784 21146 9812 21966
rect 10232 21888 10284 21894
rect 10232 21830 10284 21836
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 7012 20392 7064 20398
rect 7012 20334 7064 20340
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 7024 19718 7052 20334
rect 7116 19922 7144 20334
rect 7856 20156 8152 20176
rect 7912 20154 7936 20156
rect 7992 20154 8016 20156
rect 8072 20154 8096 20156
rect 7934 20102 7936 20154
rect 7998 20102 8010 20154
rect 8072 20102 8074 20154
rect 7912 20100 7936 20102
rect 7992 20100 8016 20102
rect 8072 20100 8096 20102
rect 7856 20080 8152 20100
rect 7104 19916 7156 19922
rect 7104 19858 7156 19864
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 7116 19514 7144 19858
rect 8036 19786 8064 19858
rect 8024 19780 8076 19786
rect 8024 19722 8076 19728
rect 7748 19712 7800 19718
rect 7748 19654 7800 19660
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 7760 19310 7788 19654
rect 8036 19310 8064 19722
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 8220 19334 8248 19654
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 8024 19304 8076 19310
rect 8220 19306 8340 19334
rect 8024 19246 8076 19252
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 6920 18828 6972 18834
rect 6920 18770 6972 18776
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 6184 18352 6236 18358
rect 6184 18294 6236 18300
rect 6092 18148 6144 18154
rect 6092 18090 6144 18096
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 6012 17134 6040 17818
rect 6104 17746 6132 18090
rect 6196 18086 6224 18294
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6656 17814 6684 18362
rect 7024 18222 7052 18566
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 6736 18148 6788 18154
rect 6736 18090 6788 18096
rect 6644 17808 6696 17814
rect 6644 17750 6696 17756
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 6104 17542 6132 17682
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 6000 17128 6052 17134
rect 6000 17070 6052 17076
rect 6104 16658 6132 17478
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 6104 12374 6132 16594
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6380 15570 6408 15846
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6656 15162 6684 17750
rect 6748 17066 6776 18090
rect 7024 17270 7052 18158
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7196 17808 7248 17814
rect 7116 17756 7196 17762
rect 7116 17750 7248 17756
rect 7116 17734 7236 17750
rect 7012 17264 7064 17270
rect 7012 17206 7064 17212
rect 7116 17202 7144 17734
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 6736 17060 6788 17066
rect 6736 17002 6788 17008
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6840 15450 6868 16934
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 6748 15422 6868 15450
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6184 14884 6236 14890
rect 6184 14826 6236 14832
rect 6196 14618 6224 14826
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 6656 14414 6684 15098
rect 6748 15026 6776 15422
rect 7024 15094 7052 15506
rect 7012 15088 7064 15094
rect 7012 15030 7064 15036
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6840 14822 6868 14894
rect 6828 14816 6880 14822
rect 6748 14776 6828 14804
rect 6748 14482 6776 14776
rect 6828 14758 6880 14764
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6472 12374 6500 13330
rect 6656 12918 6684 13330
rect 6840 13326 6868 14554
rect 6932 13530 6960 14894
rect 7024 14482 7052 15030
rect 7116 14550 7144 15982
rect 7208 15706 7236 17614
rect 7300 17270 7328 18022
rect 7392 17678 7420 18770
rect 7576 18086 7604 18770
rect 7668 18358 7696 19110
rect 7760 18766 7788 19246
rect 7856 19068 8152 19088
rect 7912 19066 7936 19068
rect 7992 19066 8016 19068
rect 8072 19066 8096 19068
rect 7934 19014 7936 19066
rect 7998 19014 8010 19066
rect 8072 19014 8074 19066
rect 7912 19012 7936 19014
rect 7992 19012 8016 19014
rect 8072 19012 8096 19014
rect 7856 18992 8152 19012
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 8116 18760 8168 18766
rect 8116 18702 8168 18708
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7564 18080 7616 18086
rect 7564 18022 7616 18028
rect 7576 17814 7604 18022
rect 7564 17808 7616 17814
rect 7564 17750 7616 17756
rect 7668 17746 7696 18294
rect 7760 17746 7788 18566
rect 8128 18222 8156 18702
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 7856 17980 8152 18000
rect 7912 17978 7936 17980
rect 7992 17978 8016 17980
rect 8072 17978 8096 17980
rect 7934 17926 7936 17978
rect 7998 17926 8010 17978
rect 8072 17926 8074 17978
rect 7912 17924 7936 17926
rect 7992 17924 8016 17926
rect 8072 17924 8096 17926
rect 7856 17904 8152 17924
rect 8220 17882 8248 18566
rect 8312 18290 8340 19306
rect 8404 18306 8432 20402
rect 9404 20324 9456 20330
rect 9404 20266 9456 20272
rect 9416 20058 9444 20266
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 9784 19922 9812 21082
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 8300 18284 8352 18290
rect 8404 18278 8524 18306
rect 8300 18226 8352 18232
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 7656 17604 7708 17610
rect 7656 17546 7708 17552
rect 7288 17264 7340 17270
rect 7288 17206 7340 17212
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7300 15570 7328 15846
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7208 14618 7236 15506
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 7104 14544 7156 14550
rect 7104 14486 7156 14492
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6736 13184 6788 13190
rect 6840 13172 6868 13262
rect 7116 13258 7144 14486
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 6788 13144 6868 13172
rect 6736 13126 6788 13132
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6092 12368 6144 12374
rect 6092 12310 6144 12316
rect 6460 12368 6512 12374
rect 6460 12310 6512 12316
rect 6104 11150 6132 12310
rect 6656 11626 6684 12854
rect 6840 12782 6868 13144
rect 6920 13184 6972 13190
rect 6972 13132 7144 13138
rect 6920 13126 7144 13132
rect 6932 13110 7144 13126
rect 7116 12850 7144 13110
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6472 11218 6500 11290
rect 6460 11212 6512 11218
rect 6840 11200 6868 12718
rect 7116 12306 7144 12786
rect 7300 12646 7328 13330
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 6920 11212 6972 11218
rect 6840 11172 6920 11200
rect 6460 11154 6512 11160
rect 6920 11154 6972 11160
rect 7024 11150 7052 11698
rect 7116 11694 7144 12242
rect 7300 11898 7328 12582
rect 7392 12102 7420 17070
rect 7576 16182 7604 17070
rect 7668 17066 7696 17546
rect 8036 17338 8064 17614
rect 8312 17542 8340 18090
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 8312 17338 8340 17478
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 7668 16658 7696 17002
rect 8404 16998 8432 18158
rect 8496 17746 8524 18278
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8484 17740 8536 17746
rect 8484 17682 8536 17688
rect 8680 17542 8708 18022
rect 8864 17882 8892 18226
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 9496 17740 9548 17746
rect 9496 17682 9548 17688
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8680 17134 8708 17478
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 7856 16892 8152 16912
rect 7912 16890 7936 16892
rect 7992 16890 8016 16892
rect 8072 16890 8096 16892
rect 7934 16838 7936 16890
rect 7998 16838 8010 16890
rect 8072 16838 8074 16890
rect 7912 16836 7936 16838
rect 7992 16836 8016 16838
rect 8072 16836 8096 16838
rect 7856 16816 8152 16836
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7564 16176 7616 16182
rect 7564 16118 7616 16124
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7484 15366 7512 16050
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7576 15026 7604 16118
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7484 14482 7512 14962
rect 7576 14822 7604 14962
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7576 13190 7604 14486
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7576 12782 7604 13126
rect 7668 12782 7696 16594
rect 7856 15804 8152 15824
rect 7912 15802 7936 15804
rect 7992 15802 8016 15804
rect 8072 15802 8096 15804
rect 7934 15750 7936 15802
rect 7998 15750 8010 15802
rect 8072 15750 8074 15802
rect 7912 15748 7936 15750
rect 7992 15748 8016 15750
rect 8072 15748 8096 15750
rect 7856 15728 8152 15748
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7760 14550 7788 14894
rect 7856 14716 8152 14736
rect 7912 14714 7936 14716
rect 7992 14714 8016 14716
rect 8072 14714 8096 14716
rect 7934 14662 7936 14714
rect 7998 14662 8010 14714
rect 8072 14662 8074 14714
rect 7912 14660 7936 14662
rect 7992 14660 8016 14662
rect 8072 14660 8096 14662
rect 7856 14640 8152 14660
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 8220 14482 8248 15506
rect 8312 14618 8340 15506
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 7856 13628 8152 13648
rect 7912 13626 7936 13628
rect 7992 13626 8016 13628
rect 8072 13626 8096 13628
rect 7934 13574 7936 13626
rect 7998 13574 8010 13626
rect 8072 13574 8074 13626
rect 7912 13572 7936 13574
rect 7992 13572 8016 13574
rect 8072 13572 8096 13574
rect 7856 13552 8152 13572
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 4896 9444 4948 9450
rect 4896 9386 4948 9392
rect 4908 8634 4936 9386
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5276 8838 5304 9318
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5092 8634 5120 8774
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5276 8430 5304 8774
rect 5460 8634 5488 9998
rect 6656 9994 6684 11086
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6932 10130 6960 10746
rect 7024 10266 7052 11086
rect 7116 11014 7144 11630
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6644 9988 6696 9994
rect 6644 9930 6696 9936
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5552 9586 5580 9862
rect 6932 9722 6960 10066
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5552 9042 5580 9522
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5736 9110 5764 9454
rect 5724 9104 5776 9110
rect 5724 9046 5776 9052
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5460 7342 5488 8570
rect 6104 8090 6132 8978
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4406 6556 4702 6576
rect 4462 6554 4486 6556
rect 4542 6554 4566 6556
rect 4622 6554 4646 6556
rect 4484 6502 4486 6554
rect 4548 6502 4560 6554
rect 4622 6502 4624 6554
rect 4462 6500 4486 6502
rect 4542 6500 4566 6502
rect 4622 6500 4646 6502
rect 4406 6480 4702 6500
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 4080 5098 4108 6122
rect 4448 6118 4476 6190
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4448 5710 4476 6054
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4406 5468 4702 5488
rect 4462 5466 4486 5468
rect 4542 5466 4566 5468
rect 4622 5466 4646 5468
rect 4484 5414 4486 5466
rect 4548 5414 4560 5466
rect 4622 5414 4624 5466
rect 4462 5412 4486 5414
rect 4542 5412 4566 5414
rect 4622 5412 4646 5414
rect 4406 5392 4702 5412
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 4080 4826 4108 5034
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4406 4380 4702 4400
rect 4462 4378 4486 4380
rect 4542 4378 4566 4380
rect 4622 4378 4646 4380
rect 4484 4326 4486 4378
rect 4548 4326 4560 4378
rect 4622 4326 4624 4378
rect 4462 4324 4486 4326
rect 4542 4324 4566 4326
rect 4622 4324 4646 4326
rect 4406 4304 4702 4324
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 2516 2990 2544 3334
rect 4406 3292 4702 3312
rect 4462 3290 4486 3292
rect 4542 3290 4566 3292
rect 4622 3290 4646 3292
rect 4484 3238 4486 3290
rect 4548 3238 4560 3290
rect 4622 3238 4624 3290
rect 4462 3236 4486 3238
rect 4542 3236 4566 3238
rect 4622 3236 4646 3238
rect 4406 3216 4702 3236
rect 4908 3194 4936 6734
rect 5736 6186 5764 7278
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 5736 5778 5764 6122
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 5736 5370 5764 5714
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 6012 4690 6040 5034
rect 6656 4826 6684 5714
rect 6932 5370 6960 6802
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6012 3670 6040 4626
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 4436 2984 4488 2990
rect 4436 2926 4488 2932
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 2332 2650 2360 2926
rect 4448 2650 4476 2926
rect 6840 2650 6868 2926
rect 6932 2650 6960 3538
rect 7024 3194 7052 9998
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7116 9042 7144 9862
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7116 7954 7144 8978
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7208 7002 7236 11086
rect 7392 10742 7420 12038
rect 7484 10810 7512 12174
rect 7576 11626 7604 12718
rect 7760 12306 7788 13466
rect 8404 12714 8432 16934
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8588 14074 8616 15438
rect 8864 15434 8892 16050
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 8852 15428 8904 15434
rect 8852 15370 8904 15376
rect 8956 15162 8984 15506
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 8956 13870 8984 15098
rect 9048 14958 9076 15982
rect 9508 15570 9536 17682
rect 9600 17626 9628 18226
rect 9784 18222 9812 19858
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 9784 17814 9812 18022
rect 10060 17814 10088 18022
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 10048 17808 10100 17814
rect 10048 17750 10100 17756
rect 9600 17598 9720 17626
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9496 15564 9548 15570
rect 9496 15506 9548 15512
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 9048 14618 9076 14894
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 9508 13326 9536 14554
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9416 12986 9444 13194
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9416 12866 9444 12922
rect 9324 12838 9444 12866
rect 9508 12850 9536 13262
rect 9600 13258 9628 17478
rect 9692 16114 9720 17598
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 9692 15162 9720 16050
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9784 15638 9812 15846
rect 9772 15632 9824 15638
rect 9772 15574 9824 15580
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9968 15026 9996 15302
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9692 14550 9720 14894
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 10152 14482 10180 15302
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 10244 13682 10272 21830
rect 10336 13870 10364 22374
rect 13096 22098 13124 22374
rect 14756 22332 15052 22352
rect 14812 22330 14836 22332
rect 14892 22330 14916 22332
rect 14972 22330 14996 22332
rect 14834 22278 14836 22330
rect 14898 22278 14910 22330
rect 14972 22278 14974 22330
rect 14812 22276 14836 22278
rect 14892 22276 14916 22278
rect 14972 22276 14996 22278
rect 14756 22256 15052 22276
rect 12072 22092 12124 22098
rect 12072 22034 12124 22040
rect 13084 22092 13136 22098
rect 13084 22034 13136 22040
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 10704 21622 10732 21966
rect 10968 21888 11020 21894
rect 10968 21830 11020 21836
rect 10692 21616 10744 21622
rect 10692 21558 10744 21564
rect 10980 21418 11008 21830
rect 11072 21690 11100 21966
rect 11306 21788 11602 21808
rect 11362 21786 11386 21788
rect 11442 21786 11466 21788
rect 11522 21786 11546 21788
rect 11384 21734 11386 21786
rect 11448 21734 11460 21786
rect 11522 21734 11524 21786
rect 11362 21732 11386 21734
rect 11442 21732 11466 21734
rect 11522 21732 11546 21734
rect 11306 21712 11602 21732
rect 12084 21690 12112 22034
rect 12256 22024 12308 22030
rect 12256 21966 12308 21972
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 10968 21412 11020 21418
rect 10968 21354 11020 21360
rect 10600 21344 10652 21350
rect 10600 21286 10652 21292
rect 10876 21344 10928 21350
rect 10876 21286 10928 21292
rect 10612 21010 10640 21286
rect 10888 21146 10916 21286
rect 10876 21140 10928 21146
rect 10876 21082 10928 21088
rect 10980 21078 11008 21354
rect 10968 21072 11020 21078
rect 10968 21014 11020 21020
rect 10600 21004 10652 21010
rect 10600 20946 10652 20952
rect 10784 21004 10836 21010
rect 10784 20946 10836 20952
rect 10796 20262 10824 20946
rect 10980 20466 11008 21014
rect 11072 21010 11100 21490
rect 12268 21486 12296 21966
rect 15200 21956 15252 21962
rect 15200 21898 15252 21904
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 12256 21480 12308 21486
rect 12256 21422 12308 21428
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 11072 20534 11100 20946
rect 11060 20528 11112 20534
rect 11060 20470 11112 20476
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 11164 20398 11192 21422
rect 12348 20936 12400 20942
rect 12348 20878 12400 20884
rect 11796 20800 11848 20806
rect 11796 20742 11848 20748
rect 11306 20700 11602 20720
rect 11362 20698 11386 20700
rect 11442 20698 11466 20700
rect 11522 20698 11546 20700
rect 11384 20646 11386 20698
rect 11448 20646 11460 20698
rect 11522 20646 11524 20698
rect 11362 20644 11386 20646
rect 11442 20644 11466 20646
rect 11522 20644 11546 20646
rect 11306 20624 11602 20644
rect 11152 20392 11204 20398
rect 11244 20392 11296 20398
rect 11204 20352 11244 20380
rect 11152 20334 11204 20340
rect 11244 20334 11296 20340
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11306 19612 11602 19632
rect 11362 19610 11386 19612
rect 11442 19610 11466 19612
rect 11522 19610 11546 19612
rect 11384 19558 11386 19610
rect 11448 19558 11460 19610
rect 11522 19558 11524 19610
rect 11362 19556 11386 19558
rect 11442 19556 11466 19558
rect 11522 19556 11546 19558
rect 11306 19536 11602 19556
rect 11716 18834 11744 19654
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11306 18524 11602 18544
rect 11362 18522 11386 18524
rect 11442 18522 11466 18524
rect 11522 18522 11546 18524
rect 11384 18470 11386 18522
rect 11448 18470 11460 18522
rect 11522 18470 11524 18522
rect 11362 18468 11386 18470
rect 11442 18468 11466 18470
rect 11522 18468 11546 18470
rect 11306 18448 11602 18468
rect 11808 18222 11836 20742
rect 12360 19310 12388 20878
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 12452 19310 12480 19858
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 12622 19408 12678 19417
rect 12622 19343 12624 19352
rect 12676 19343 12678 19352
rect 12624 19314 12676 19320
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 11992 18408 12020 18770
rect 12268 18426 12296 18770
rect 11900 18380 12020 18408
rect 12072 18420 12124 18426
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 10520 16046 10548 18158
rect 11808 17814 11836 18158
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11306 17436 11602 17456
rect 11362 17434 11386 17436
rect 11442 17434 11466 17436
rect 11522 17434 11546 17436
rect 11384 17382 11386 17434
rect 11448 17382 11460 17434
rect 11522 17382 11524 17434
rect 11362 17380 11386 17382
rect 11442 17380 11466 17382
rect 11522 17380 11546 17382
rect 11306 17360 11602 17380
rect 11900 17338 11928 18380
rect 12072 18362 12124 18368
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 11992 17746 12020 18226
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 12084 17678 12112 18362
rect 12164 18148 12216 18154
rect 12164 18090 12216 18096
rect 12176 17814 12204 18090
rect 12636 17882 12664 19314
rect 13188 19310 13216 19790
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 12716 19236 12768 19242
rect 12716 19178 12768 19184
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12992 19236 13044 19242
rect 12992 19178 13044 19184
rect 12728 18970 12756 19178
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 12820 18902 12848 19178
rect 12808 18896 12860 18902
rect 12808 18838 12860 18844
rect 12820 18426 12848 18838
rect 13004 18834 13032 19178
rect 13188 18970 13216 19246
rect 13176 18964 13228 18970
rect 13176 18906 13228 18912
rect 12992 18828 13044 18834
rect 12992 18770 13044 18776
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12164 17808 12216 17814
rect 12164 17750 12216 17756
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11796 17060 11848 17066
rect 11796 17002 11848 17008
rect 11808 16658 11836 17002
rect 11900 16794 11928 17274
rect 12176 16794 12204 17750
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 12452 16726 12480 17002
rect 12440 16720 12492 16726
rect 12440 16662 12492 16668
rect 12808 16720 12860 16726
rect 12808 16662 12860 16668
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11306 16348 11602 16368
rect 11362 16346 11386 16348
rect 11442 16346 11466 16348
rect 11522 16346 11546 16348
rect 11384 16294 11386 16346
rect 11448 16294 11460 16346
rect 11522 16294 11524 16346
rect 11362 16292 11386 16294
rect 11442 16292 11466 16294
rect 11522 16292 11546 16294
rect 11306 16272 11602 16292
rect 11808 16250 11836 16594
rect 12820 16250 12848 16662
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10796 15638 10824 15846
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 10980 15094 11008 15982
rect 11306 15260 11602 15280
rect 11362 15258 11386 15260
rect 11442 15258 11466 15260
rect 11522 15258 11546 15260
rect 11384 15206 11386 15258
rect 11448 15206 11460 15258
rect 11522 15206 11524 15258
rect 11362 15204 11386 15206
rect 11442 15204 11466 15206
rect 11522 15204 11546 15206
rect 11306 15184 11602 15204
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 10600 14884 10652 14890
rect 10600 14826 10652 14832
rect 10612 14618 10640 14826
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 9876 13530 9904 13670
rect 10244 13654 10364 13682
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9496 12844 9548 12850
rect 8392 12708 8444 12714
rect 8392 12650 8444 12656
rect 7856 12540 8152 12560
rect 7912 12538 7936 12540
rect 7992 12538 8016 12540
rect 8072 12538 8096 12540
rect 7934 12486 7936 12538
rect 7998 12486 8010 12538
rect 8072 12486 8074 12538
rect 7912 12484 7936 12486
rect 7992 12484 8016 12486
rect 8072 12484 8096 12486
rect 7856 12464 8152 12484
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7564 11620 7616 11626
rect 7564 11562 7616 11568
rect 7576 11150 7604 11562
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7760 11234 7788 11494
rect 7856 11452 8152 11472
rect 7912 11450 7936 11452
rect 7992 11450 8016 11452
rect 8072 11450 8096 11452
rect 7934 11398 7936 11450
rect 7998 11398 8010 11450
rect 8072 11398 8074 11450
rect 7912 11396 7936 11398
rect 7992 11396 8016 11398
rect 8072 11396 8096 11398
rect 7856 11376 8152 11396
rect 7760 11218 7880 11234
rect 7760 11212 7892 11218
rect 7760 11206 7840 11212
rect 7840 11154 7892 11160
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7668 11014 7696 11086
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 8404 10810 8432 12650
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8496 11014 8524 11630
rect 8772 11218 8800 11630
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 10810 8524 10950
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 8404 10554 8432 10746
rect 8496 10674 8524 10746
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8772 10606 8800 11154
rect 9140 10674 9168 11494
rect 9324 11218 9352 12838
rect 9496 12786 9548 12792
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 8760 10600 8812 10606
rect 8404 10538 8524 10554
rect 8760 10542 8812 10548
rect 8404 10532 8536 10538
rect 8404 10526 8484 10532
rect 8484 10474 8536 10480
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 7856 10364 8152 10384
rect 7912 10362 7936 10364
rect 7992 10362 8016 10364
rect 8072 10362 8096 10364
rect 7934 10310 7936 10362
rect 7998 10310 8010 10362
rect 8072 10310 8074 10362
rect 7912 10308 7936 10310
rect 7992 10308 8016 10310
rect 8072 10308 8096 10310
rect 7856 10288 8152 10308
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 9178 7328 9318
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7576 9110 7604 9862
rect 7668 9518 7696 9930
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 8680 9450 8708 10406
rect 8852 10192 8904 10198
rect 8852 10134 8904 10140
rect 8864 9722 8892 10134
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 9140 9518 9168 10610
rect 9416 10130 9444 12718
rect 9508 12306 9536 12786
rect 9600 12714 9628 13194
rect 10060 13172 10088 13330
rect 10140 13184 10192 13190
rect 10060 13144 10140 13172
rect 10192 13144 10272 13172
rect 10140 13126 10192 13132
rect 9588 12708 9640 12714
rect 9588 12650 9640 12656
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9600 10062 9628 12650
rect 10244 12306 10272 13144
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9876 11762 9904 12174
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9692 11218 9720 11562
rect 9876 11218 9904 11698
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9600 9586 9628 9862
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 7856 9276 8152 9296
rect 7912 9274 7936 9276
rect 7992 9274 8016 9276
rect 8072 9274 8096 9276
rect 7934 9222 7936 9274
rect 7998 9222 8010 9274
rect 8072 9222 8074 9274
rect 7912 9220 7936 9222
rect 7992 9220 8016 9222
rect 8072 9220 8096 9222
rect 7856 9200 8152 9220
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7104 5840 7156 5846
rect 7104 5782 7156 5788
rect 7116 5166 7144 5782
rect 7300 5778 7328 6054
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7668 4078 7696 8774
rect 7856 8188 8152 8208
rect 7912 8186 7936 8188
rect 7992 8186 8016 8188
rect 8072 8186 8096 8188
rect 7934 8134 7936 8186
rect 7998 8134 8010 8186
rect 8072 8134 8074 8186
rect 7912 8132 7936 8134
rect 7992 8132 8016 8134
rect 8072 8132 8096 8134
rect 7856 8112 8152 8132
rect 7856 7100 8152 7120
rect 7912 7098 7936 7100
rect 7992 7098 8016 7100
rect 8072 7098 8096 7100
rect 7934 7046 7936 7098
rect 7998 7046 8010 7098
rect 8072 7046 8074 7098
rect 7912 7044 7936 7046
rect 7992 7044 8016 7046
rect 8072 7044 8096 7046
rect 7856 7024 8152 7044
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 7856 6012 8152 6032
rect 7912 6010 7936 6012
rect 7992 6010 8016 6012
rect 8072 6010 8096 6012
rect 7934 5958 7936 6010
rect 7998 5958 8010 6010
rect 8072 5958 8074 6010
rect 7912 5956 7936 5958
rect 7992 5956 8016 5958
rect 8072 5956 8096 5958
rect 7856 5936 8152 5956
rect 8220 5846 8248 6122
rect 8680 6118 8708 9386
rect 9600 8906 9628 9522
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 9508 5778 9536 8774
rect 9600 8634 9628 8842
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9692 8090 9720 9318
rect 9784 9110 9812 9386
rect 10336 9178 10364 13654
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10416 12300 10468 12306
rect 10520 12288 10548 13330
rect 10612 13258 10640 14554
rect 11440 14550 11468 14758
rect 12360 14618 12388 14758
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 11428 14544 11480 14550
rect 11428 14486 11480 14492
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10600 13252 10652 13258
rect 10600 13194 10652 13200
rect 10612 12782 10640 13194
rect 10704 12986 10732 13738
rect 10796 13326 10824 14418
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 11164 13870 11192 14350
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 11306 14172 11602 14192
rect 11362 14170 11386 14172
rect 11442 14170 11466 14172
rect 11522 14170 11546 14172
rect 11384 14118 11386 14170
rect 11448 14118 11460 14170
rect 11522 14118 11524 14170
rect 11362 14116 11386 14118
rect 11442 14116 11466 14118
rect 11522 14116 11546 14118
rect 11306 14096 11602 14116
rect 12256 13932 12308 13938
rect 12256 13874 12308 13880
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10796 12850 10824 13262
rect 11164 12918 11192 13330
rect 11306 13084 11602 13104
rect 11362 13082 11386 13084
rect 11442 13082 11466 13084
rect 11522 13082 11546 13084
rect 11384 13030 11386 13082
rect 11448 13030 11460 13082
rect 11522 13030 11524 13082
rect 11362 13028 11386 13030
rect 11442 13028 11466 13030
rect 11522 13028 11546 13030
rect 11306 13008 11602 13028
rect 11152 12912 11204 12918
rect 11152 12854 11204 12860
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10600 12776 10652 12782
rect 10652 12724 10732 12730
rect 10600 12718 10732 12724
rect 10612 12702 10732 12718
rect 10600 12300 10652 12306
rect 10520 12260 10600 12288
rect 10416 12242 10468 12248
rect 10600 12242 10652 12248
rect 10428 11762 10456 12242
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10520 11642 10548 12038
rect 10428 11614 10548 11642
rect 10428 10810 10456 11614
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10428 9450 10456 10746
rect 10520 10538 10548 11222
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 10520 10130 10548 10474
rect 10612 10470 10640 12242
rect 10704 12238 10732 12702
rect 10796 12434 10824 12786
rect 11164 12782 11192 12854
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10796 12406 10916 12434
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10704 11286 10732 11630
rect 10784 11620 10836 11626
rect 10784 11562 10836 11568
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10520 9722 10548 10066
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9784 8498 9812 9046
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9876 8634 9904 8978
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 10244 7954 10272 8910
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 8680 5098 8708 5714
rect 9508 5234 9536 5714
rect 9692 5370 9720 5850
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 7856 4924 8152 4944
rect 7912 4922 7936 4924
rect 7992 4922 8016 4924
rect 8072 4922 8096 4924
rect 7934 4870 7936 4922
rect 7998 4870 8010 4922
rect 8072 4870 8074 4922
rect 7912 4868 7936 4870
rect 7992 4868 8016 4870
rect 8072 4868 8096 4870
rect 7856 4848 8152 4868
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7668 3602 7696 4014
rect 8680 4010 8708 5034
rect 8668 4004 8720 4010
rect 8668 3946 8720 3952
rect 7856 3836 8152 3856
rect 7912 3834 7936 3836
rect 7992 3834 8016 3836
rect 8072 3834 8096 3836
rect 7934 3782 7936 3834
rect 7998 3782 8010 3834
rect 8072 3782 8074 3834
rect 7912 3780 7936 3782
rect 7992 3780 8016 3782
rect 8072 3780 8096 3782
rect 7856 3760 8152 3780
rect 8680 3670 8708 3946
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8588 3194 8616 3538
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9324 3194 9352 3334
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9600 3058 9628 3334
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9784 2922 9812 7822
rect 10244 6798 10272 7890
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10336 7410 10364 7686
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10244 6322 10272 6734
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10060 5846 10088 6054
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 9864 5636 9916 5642
rect 9864 5578 9916 5584
rect 9876 5370 9904 5578
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 10244 4622 10272 6258
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10428 5914 10456 6190
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9876 3126 9904 3470
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 7856 2748 8152 2768
rect 7912 2746 7936 2748
rect 7992 2746 8016 2748
rect 8072 2746 8096 2748
rect 7934 2694 7936 2746
rect 7998 2694 8010 2746
rect 8072 2694 8074 2746
rect 7912 2692 7936 2694
rect 7992 2692 8016 2694
rect 8072 2692 8096 2694
rect 7856 2672 8152 2692
rect 10428 2650 10456 4558
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10520 3602 10548 3878
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10612 2990 10640 10406
rect 10692 10124 10744 10130
rect 10796 10112 10824 11562
rect 10888 10826 10916 12406
rect 10980 12102 11008 12582
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 11306 11996 11602 12016
rect 11362 11994 11386 11996
rect 11442 11994 11466 11996
rect 11522 11994 11546 11996
rect 11384 11942 11386 11994
rect 11448 11942 11460 11994
rect 11522 11942 11524 11994
rect 11362 11940 11386 11942
rect 11442 11940 11466 11942
rect 11522 11940 11546 11942
rect 11306 11920 11602 11940
rect 11306 10908 11602 10928
rect 11362 10906 11386 10908
rect 11442 10906 11466 10908
rect 11522 10906 11546 10908
rect 11384 10854 11386 10906
rect 11448 10854 11460 10906
rect 11522 10854 11524 10906
rect 11362 10852 11386 10854
rect 11442 10852 11466 10854
rect 11522 10852 11546 10854
rect 11306 10832 11602 10852
rect 10888 10798 11008 10826
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 10888 10198 10916 10678
rect 10980 10538 11008 10798
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 10968 10532 11020 10538
rect 10968 10474 11020 10480
rect 10876 10192 10928 10198
rect 10876 10134 10928 10140
rect 10744 10084 10824 10112
rect 10692 10066 10744 10072
rect 10704 9518 10732 10066
rect 10980 9518 11008 10474
rect 11306 9820 11602 9840
rect 11362 9818 11386 9820
rect 11442 9818 11466 9820
rect 11522 9818 11546 9820
rect 11384 9766 11386 9818
rect 11448 9766 11460 9818
rect 11522 9766 11524 9818
rect 11362 9764 11386 9766
rect 11442 9764 11466 9766
rect 11522 9764 11546 9766
rect 11306 9744 11602 9764
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10980 9110 11008 9454
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10704 4826 10732 8774
rect 10888 8430 10916 8461
rect 10876 8424 10928 8430
rect 10980 8378 11008 9046
rect 11306 8732 11602 8752
rect 11362 8730 11386 8732
rect 11442 8730 11466 8732
rect 11522 8730 11546 8732
rect 11384 8678 11386 8730
rect 11448 8678 11460 8730
rect 11522 8678 11524 8730
rect 11362 8676 11386 8678
rect 11442 8676 11466 8678
rect 11522 8676 11546 8678
rect 11306 8656 11602 8676
rect 10928 8372 11008 8378
rect 10876 8366 11008 8372
rect 10888 8350 11008 8366
rect 10888 8090 10916 8350
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 10888 7342 10916 7890
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10888 7002 10916 7278
rect 10980 7274 11008 8230
rect 11072 7478 11100 8230
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 11164 7206 11192 7958
rect 11306 7644 11602 7664
rect 11362 7642 11386 7644
rect 11442 7642 11466 7644
rect 11522 7642 11546 7644
rect 11384 7590 11386 7642
rect 11448 7590 11460 7642
rect 11522 7590 11524 7642
rect 11362 7588 11386 7590
rect 11442 7588 11466 7590
rect 11522 7588 11546 7590
rect 11306 7568 11602 7588
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11716 7002 11744 10542
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11900 7954 11928 8774
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11808 7546 11836 7686
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11900 7410 11928 7890
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11992 6662 12020 13806
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12176 12714 12204 13262
rect 12268 12850 12296 13874
rect 12912 13258 12940 14214
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 12176 12442 12204 12650
rect 12268 12442 12296 12786
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 12360 12322 12388 12582
rect 12544 12442 12572 12582
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12176 12306 12388 12322
rect 12636 12306 12664 13126
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12164 12300 12388 12306
rect 12216 12294 12388 12300
rect 12624 12300 12676 12306
rect 12164 12242 12216 12248
rect 12624 12242 12676 12248
rect 12176 11354 12204 12242
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12360 11150 12388 12174
rect 12912 11762 12940 12582
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12912 11218 12940 11698
rect 13280 11354 13308 11766
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 13188 10674 13216 11018
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 13188 10418 13216 10610
rect 13280 10606 13308 11290
rect 13372 10674 13400 21830
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 14016 20602 14044 21490
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 13728 19780 13780 19786
rect 13728 19722 13780 19728
rect 13740 18902 13768 19722
rect 13728 18896 13780 18902
rect 13728 18838 13780 18844
rect 13832 18834 13860 19790
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14108 19378 14136 19654
rect 14200 19378 14228 19790
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13832 17814 13860 18770
rect 14108 18290 14136 19314
rect 14292 19310 14320 21558
rect 14660 21418 14688 21830
rect 15108 21548 15160 21554
rect 15108 21490 15160 21496
rect 14648 21412 14700 21418
rect 14648 21354 14700 21360
rect 14756 21244 15052 21264
rect 14812 21242 14836 21244
rect 14892 21242 14916 21244
rect 14972 21242 14996 21244
rect 14834 21190 14836 21242
rect 14898 21190 14910 21242
rect 14972 21190 14974 21242
rect 14812 21188 14836 21190
rect 14892 21188 14916 21190
rect 14972 21188 14996 21190
rect 14756 21168 15052 21188
rect 14556 20528 14608 20534
rect 14556 20470 14608 20476
rect 14464 20324 14516 20330
rect 14464 20266 14516 20272
rect 14476 20058 14504 20266
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14384 19310 14412 19450
rect 14476 19378 14504 19994
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14372 19304 14424 19310
rect 14568 19281 14596 20470
rect 15120 20398 15148 21490
rect 15212 21350 15240 21898
rect 15396 21486 15424 22374
rect 16040 21486 16068 22374
rect 16684 22098 16712 22374
rect 16672 22092 16724 22098
rect 16672 22034 16724 22040
rect 17592 22024 17644 22030
rect 17592 21966 17644 21972
rect 17684 22024 17736 22030
rect 17736 21984 17816 22012
rect 17684 21966 17736 21972
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 16868 21554 16896 21830
rect 17604 21690 17632 21966
rect 17592 21684 17644 21690
rect 17592 21626 17644 21632
rect 16856 21548 16908 21554
rect 16856 21490 16908 21496
rect 15384 21480 15436 21486
rect 15384 21422 15436 21428
rect 16028 21480 16080 21486
rect 16028 21422 16080 21428
rect 15200 21344 15252 21350
rect 15200 21286 15252 21292
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 15212 21010 15240 21286
rect 15568 21072 15620 21078
rect 15568 21014 15620 21020
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 15108 20392 15160 20398
rect 15108 20334 15160 20340
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14660 19854 14688 20198
rect 14756 20156 15052 20176
rect 14812 20154 14836 20156
rect 14892 20154 14916 20156
rect 14972 20154 14996 20156
rect 14834 20102 14836 20154
rect 14898 20102 14910 20154
rect 14972 20102 14974 20154
rect 14812 20100 14836 20102
rect 14892 20100 14916 20102
rect 14972 20100 14996 20102
rect 14756 20080 15052 20100
rect 15120 19938 15148 20334
rect 14936 19922 15148 19938
rect 15200 19984 15252 19990
rect 15200 19926 15252 19932
rect 14924 19916 15148 19922
rect 14976 19910 15148 19916
rect 14924 19858 14976 19864
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 15212 19514 15240 19926
rect 15488 19786 15516 20878
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15108 19304 15160 19310
rect 14372 19246 14424 19252
rect 14554 19272 14610 19281
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 14292 18222 14320 19246
rect 15108 19246 15160 19252
rect 15198 19272 15254 19281
rect 14554 19207 14610 19216
rect 14756 19068 15052 19088
rect 14812 19066 14836 19068
rect 14892 19066 14916 19068
rect 14972 19066 14996 19068
rect 14834 19014 14836 19066
rect 14898 19014 14910 19066
rect 14972 19014 14974 19066
rect 14812 19012 14836 19014
rect 14892 19012 14916 19014
rect 14972 19012 14996 19014
rect 14756 18992 15052 19012
rect 15120 18630 15148 19246
rect 15198 19207 15254 19216
rect 15108 18624 15160 18630
rect 15108 18566 15160 18572
rect 14280 18216 14332 18222
rect 14280 18158 14332 18164
rect 14096 18148 14148 18154
rect 14096 18090 14148 18096
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 13820 17808 13872 17814
rect 13820 17750 13872 17756
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 13648 16794 13676 17682
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 13648 16658 13676 16730
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13648 15910 13676 16594
rect 13832 16522 13860 17614
rect 13924 16998 13952 17818
rect 14108 17610 14136 18090
rect 14756 17980 15052 18000
rect 14812 17978 14836 17980
rect 14892 17978 14916 17980
rect 14972 17978 14996 17980
rect 14834 17926 14836 17978
rect 14898 17926 14910 17978
rect 14972 17926 14974 17978
rect 14812 17924 14836 17926
rect 14892 17924 14916 17926
rect 14972 17924 14996 17926
rect 14756 17904 15052 17924
rect 14096 17604 14148 17610
rect 14096 17546 14148 17552
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13924 16658 13952 16934
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13820 16516 13872 16522
rect 13820 16458 13872 16464
rect 13832 16046 13860 16458
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 14016 15978 14044 17478
rect 14004 15972 14056 15978
rect 14004 15914 14056 15920
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 14016 15162 14044 15914
rect 14108 15706 14136 17546
rect 14756 16892 15052 16912
rect 14812 16890 14836 16892
rect 14892 16890 14916 16892
rect 14972 16890 14996 16892
rect 14834 16838 14836 16890
rect 14898 16838 14910 16890
rect 14972 16838 14974 16890
rect 14812 16836 14836 16838
rect 14892 16836 14916 16838
rect 14972 16836 14996 16838
rect 14756 16816 15052 16836
rect 15212 16658 15240 19207
rect 15580 18766 15608 21014
rect 15752 20324 15804 20330
rect 15752 20266 15804 20272
rect 15764 19922 15792 20266
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 15660 19304 15712 19310
rect 15658 19272 15660 19281
rect 15712 19272 15714 19281
rect 15658 19207 15714 19216
rect 15672 19174 15700 19207
rect 15660 19168 15712 19174
rect 15764 19145 15792 19858
rect 15660 19110 15712 19116
rect 15750 19136 15806 19145
rect 15750 19071 15806 19080
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15580 17134 15608 18702
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 15304 16794 15332 17002
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15580 16658 15608 17070
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 14648 16652 14700 16658
rect 14648 16594 14700 16600
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 14384 16046 14412 16594
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 14004 15156 14056 15162
rect 14004 15098 14056 15104
rect 14108 15042 14136 15302
rect 14660 15065 14688 16594
rect 15488 15978 15516 16594
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 14756 15804 15052 15824
rect 14812 15802 14836 15804
rect 14892 15802 14916 15804
rect 14972 15802 14996 15804
rect 14834 15750 14836 15802
rect 14898 15750 14910 15802
rect 14972 15750 14974 15802
rect 14812 15748 14836 15750
rect 14892 15748 14916 15750
rect 14972 15748 14996 15750
rect 14756 15728 15052 15748
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15304 15162 15332 15438
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15396 15094 15424 15438
rect 15200 15088 15252 15094
rect 14016 15014 14136 15042
rect 14646 15056 14702 15065
rect 14016 13870 14044 15014
rect 15384 15088 15436 15094
rect 15200 15030 15252 15036
rect 15290 15056 15346 15065
rect 14646 14991 14702 15000
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14568 14550 14596 14758
rect 14660 14618 14688 14894
rect 14756 14716 15052 14736
rect 14812 14714 14836 14716
rect 14892 14714 14916 14716
rect 14972 14714 14996 14716
rect 14834 14662 14836 14714
rect 14898 14662 14910 14714
rect 14972 14662 14974 14714
rect 14812 14660 14836 14662
rect 14892 14660 14916 14662
rect 14972 14660 14996 14662
rect 14756 14640 15052 14660
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 15016 14544 15068 14550
rect 15016 14486 15068 14492
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14292 13938 14320 14214
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 14016 13258 14044 13806
rect 14568 13462 14596 14486
rect 15028 14074 15056 14486
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 14756 13628 15052 13648
rect 14812 13626 14836 13628
rect 14892 13626 14916 13628
rect 14972 13626 14996 13628
rect 14834 13574 14836 13626
rect 14898 13574 14910 13626
rect 14972 13574 14974 13626
rect 14812 13572 14836 13574
rect 14892 13572 14916 13574
rect 14972 13572 14996 13574
rect 14756 13552 15052 13572
rect 15120 13530 15148 14894
rect 15212 14618 15240 15030
rect 15384 15030 15436 15036
rect 15290 14991 15346 15000
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15304 14521 15332 14991
rect 15290 14512 15346 14521
rect 15290 14447 15292 14456
rect 15344 14447 15346 14456
rect 15292 14418 15344 14424
rect 15488 14414 15516 15914
rect 15580 15366 15608 16594
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15764 14618 15792 16934
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15580 13530 15608 13738
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 14556 13456 14608 13462
rect 14556 13398 14608 13404
rect 15764 13394 15792 14554
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 13556 12782 13584 13194
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 14756 12540 15052 12560
rect 14812 12538 14836 12540
rect 14892 12538 14916 12540
rect 14972 12538 14996 12540
rect 14834 12486 14836 12538
rect 14898 12486 14910 12538
rect 14972 12486 14974 12538
rect 14812 12484 14836 12486
rect 14892 12484 14916 12486
rect 14972 12484 14996 12486
rect 14756 12464 15052 12484
rect 15120 12442 15148 12582
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15764 12306 15792 13330
rect 15856 12442 15884 21286
rect 17500 21004 17552 21010
rect 17500 20946 17552 20952
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 15936 19346 15988 19352
rect 16040 19334 16068 19858
rect 16304 19508 16356 19514
rect 16304 19450 16356 19456
rect 16120 19440 16172 19446
rect 16120 19382 16172 19388
rect 15988 19306 16068 19334
rect 15936 19288 15988 19294
rect 16040 18426 16068 19306
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 16132 18154 16160 19382
rect 16316 18902 16344 19450
rect 16304 18896 16356 18902
rect 16304 18838 16356 18844
rect 16960 18630 16988 20742
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 17328 18426 17356 18770
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 16120 18148 16172 18154
rect 16120 18090 16172 18096
rect 16224 17746 16252 18158
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16408 16998 16436 17682
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16592 16726 16620 16934
rect 17328 16726 17356 17478
rect 17420 17134 17448 18566
rect 17512 18222 17540 20946
rect 17682 19408 17738 19417
rect 17682 19343 17684 19352
rect 17736 19343 17738 19352
rect 17684 19314 17736 19320
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17604 18612 17632 19246
rect 17684 18624 17736 18630
rect 17604 18584 17684 18612
rect 17684 18566 17736 18572
rect 17696 18290 17724 18566
rect 17684 18284 17736 18290
rect 17684 18226 17736 18232
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 17512 17746 17540 18158
rect 17592 18148 17644 18154
rect 17592 18090 17644 18096
rect 17500 17740 17552 17746
rect 17500 17682 17552 17688
rect 17604 17134 17632 18090
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 16580 16720 16632 16726
rect 16580 16662 16632 16668
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16224 14482 16252 14758
rect 16960 14482 16988 16050
rect 17420 15910 17448 17070
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 17052 15162 17080 15506
rect 17512 15162 17540 16934
rect 17604 16046 17632 17070
rect 17696 17066 17724 18226
rect 17684 17060 17736 17066
rect 17684 17002 17736 17008
rect 17696 16182 17724 17002
rect 17684 16176 17736 16182
rect 17684 16118 17736 16124
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17604 15706 17632 15982
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17052 14550 17080 15098
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17040 14544 17092 14550
rect 17040 14486 17092 14492
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 16224 13462 16252 14418
rect 16960 14006 16988 14418
rect 17328 14346 17356 14894
rect 17512 14414 17540 15098
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 17328 13938 17356 14282
rect 17420 14074 17448 14350
rect 17512 14074 17540 14350
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 17316 13456 17368 13462
rect 17316 13398 17368 13404
rect 17328 12442 17356 13398
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13740 11218 13768 11494
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13924 10810 13952 11630
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13820 10464 13872 10470
rect 12544 9654 12572 10406
rect 13188 10390 13308 10418
rect 13820 10406 13872 10412
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12728 9518 12756 9998
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12452 9178 12480 9318
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12728 8906 12756 9454
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 11306 6556 11602 6576
rect 11362 6554 11386 6556
rect 11442 6554 11466 6556
rect 11522 6554 11546 6556
rect 11384 6502 11386 6554
rect 11448 6502 11460 6554
rect 11522 6502 11524 6554
rect 11362 6500 11386 6502
rect 11442 6500 11466 6502
rect 11522 6500 11546 6502
rect 11306 6480 11602 6500
rect 12268 6254 12296 6598
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12636 5778 12664 8230
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12728 6322 12756 6666
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12256 5568 12308 5574
rect 12256 5510 12308 5516
rect 11306 5468 11602 5488
rect 11362 5466 11386 5468
rect 11442 5466 11466 5468
rect 11522 5466 11546 5468
rect 11384 5414 11386 5466
rect 11448 5414 11460 5466
rect 11522 5414 11524 5466
rect 11362 5412 11386 5414
rect 11442 5412 11466 5414
rect 11522 5412 11546 5414
rect 11306 5392 11602 5412
rect 12268 5030 12296 5510
rect 12544 5166 12572 5646
rect 12636 5234 12664 5714
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10704 3058 10732 3334
rect 10796 3058 10824 4490
rect 11164 4078 11192 4762
rect 11704 4548 11756 4554
rect 11704 4490 11756 4496
rect 11306 4380 11602 4400
rect 11362 4378 11386 4380
rect 11442 4378 11466 4380
rect 11522 4378 11546 4380
rect 11384 4326 11386 4378
rect 11448 4326 11460 4378
rect 11522 4326 11524 4378
rect 11362 4324 11386 4326
rect 11442 4324 11466 4326
rect 11522 4324 11546 4326
rect 11306 4304 11602 4324
rect 11716 4282 11744 4490
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 12268 4078 12296 4966
rect 12544 4690 12572 5102
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 12256 4072 12308 4078
rect 12256 4014 12308 4020
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11306 3292 11602 3312
rect 11362 3290 11386 3292
rect 11442 3290 11466 3292
rect 11522 3290 11546 3292
rect 11384 3238 11386 3290
rect 11448 3238 11460 3290
rect 11522 3238 11524 3290
rect 11362 3236 11386 3238
rect 11442 3236 11466 3238
rect 11522 3236 11546 3238
rect 11306 3216 11602 3236
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 12084 2774 12112 3538
rect 12820 2922 12848 9930
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12912 9382 12940 9862
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 9042 12940 9318
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 13280 8974 13308 10390
rect 13832 9586 13860 10406
rect 13924 10198 13952 10746
rect 13912 10192 13964 10198
rect 13912 10134 13964 10140
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13280 8498 13308 8910
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12912 7886 12940 8366
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 13004 8090 13032 8230
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12912 6934 12940 7822
rect 13740 7546 13768 7890
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 14108 7410 14136 12038
rect 15580 11762 15608 12174
rect 15844 12164 15896 12170
rect 15844 12106 15896 12112
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 14756 11452 15052 11472
rect 14812 11450 14836 11452
rect 14892 11450 14916 11452
rect 14972 11450 14996 11452
rect 14834 11398 14836 11450
rect 14898 11398 14910 11450
rect 14972 11398 14974 11450
rect 14812 11396 14836 11398
rect 14892 11396 14916 11398
rect 14972 11396 14996 11398
rect 14756 11376 15052 11396
rect 15672 11150 15700 11698
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 15028 10742 15056 10950
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 15476 10600 15528 10606
rect 15476 10542 15528 10548
rect 14648 10464 14700 10470
rect 14648 10406 14700 10412
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 12992 7268 13044 7274
rect 12992 7210 13044 7216
rect 13004 6934 13032 7210
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12992 6928 13044 6934
rect 12992 6870 13044 6876
rect 13004 6186 13032 6870
rect 13188 6458 13216 6938
rect 13740 6458 13768 7278
rect 14660 6914 14688 10406
rect 14756 10364 15052 10384
rect 14812 10362 14836 10364
rect 14892 10362 14916 10364
rect 14972 10362 14996 10364
rect 14834 10310 14836 10362
rect 14898 10310 14910 10362
rect 14972 10310 14974 10362
rect 14812 10308 14836 10310
rect 14892 10308 14916 10310
rect 14972 10308 14996 10310
rect 14756 10288 15052 10308
rect 15488 10266 15516 10542
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15764 9722 15792 10066
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 14756 9276 15052 9296
rect 14812 9274 14836 9276
rect 14892 9274 14916 9276
rect 14972 9274 14996 9276
rect 14834 9222 14836 9274
rect 14898 9222 14910 9274
rect 14972 9222 14974 9274
rect 14812 9220 14836 9222
rect 14892 9220 14916 9222
rect 14972 9220 14996 9222
rect 14756 9200 15052 9220
rect 15120 8974 15148 9522
rect 15200 9444 15252 9450
rect 15200 9386 15252 9392
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15212 8786 15240 9386
rect 15764 9178 15792 9658
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15120 8758 15240 8786
rect 15120 8362 15148 8758
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15108 8356 15160 8362
rect 15108 8298 15160 8304
rect 14756 8188 15052 8208
rect 14812 8186 14836 8188
rect 14892 8186 14916 8188
rect 14972 8186 14996 8188
rect 14834 8134 14836 8186
rect 14898 8134 14910 8186
rect 14972 8134 14974 8186
rect 14812 8132 14836 8134
rect 14892 8132 14916 8134
rect 14972 8132 14996 8134
rect 14756 8112 15052 8132
rect 15120 8090 15148 8298
rect 15488 8090 15516 8366
rect 15856 8090 15884 12106
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16408 11218 16436 11494
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16764 11212 16816 11218
rect 16764 11154 16816 11160
rect 16776 10538 16804 11154
rect 16764 10532 16816 10538
rect 16764 10474 16816 10480
rect 16776 10266 16804 10474
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16132 8498 16160 8978
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16132 8362 16160 8434
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 17788 7342 17816 21984
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 18206 21788 18502 21808
rect 18262 21786 18286 21788
rect 18342 21786 18366 21788
rect 18422 21786 18446 21788
rect 18284 21734 18286 21786
rect 18348 21734 18360 21786
rect 18422 21734 18424 21786
rect 18262 21732 18286 21734
rect 18342 21732 18366 21734
rect 18422 21732 18446 21734
rect 18206 21712 18502 21732
rect 19996 21622 20024 21830
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 19996 21486 20024 21558
rect 19340 21480 19392 21486
rect 19340 21422 19392 21428
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 18144 21412 18196 21418
rect 18144 21354 18196 21360
rect 18156 21146 18184 21354
rect 18144 21140 18196 21146
rect 18144 21082 18196 21088
rect 18206 20700 18502 20720
rect 18262 20698 18286 20700
rect 18342 20698 18366 20700
rect 18422 20698 18446 20700
rect 18284 20646 18286 20698
rect 18348 20646 18360 20698
rect 18422 20646 18424 20698
rect 18262 20644 18286 20646
rect 18342 20644 18366 20646
rect 18422 20644 18446 20646
rect 18206 20624 18502 20644
rect 19352 20398 19380 21422
rect 19892 21344 19944 21350
rect 19892 21286 19944 21292
rect 19616 20800 19668 20806
rect 19616 20742 19668 20748
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 18206 19612 18502 19632
rect 18262 19610 18286 19612
rect 18342 19610 18366 19612
rect 18422 19610 18446 19612
rect 18284 19558 18286 19610
rect 18348 19558 18360 19610
rect 18422 19558 18424 19610
rect 18262 19556 18286 19558
rect 18342 19556 18366 19558
rect 18422 19556 18446 19558
rect 18206 19536 18502 19556
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 17880 18834 17908 19246
rect 17868 18828 17920 18834
rect 17868 18770 17920 18776
rect 17972 18426 18000 19246
rect 18604 19168 18656 19174
rect 18602 19136 18604 19145
rect 18656 19136 18658 19145
rect 18602 19071 18658 19080
rect 18206 18524 18502 18544
rect 18262 18522 18286 18524
rect 18342 18522 18366 18524
rect 18422 18522 18446 18524
rect 18284 18470 18286 18522
rect 18348 18470 18360 18522
rect 18422 18470 18424 18522
rect 18262 18468 18286 18470
rect 18342 18468 18366 18470
rect 18422 18468 18446 18470
rect 18206 18448 18502 18468
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 18206 17436 18502 17456
rect 18262 17434 18286 17436
rect 18342 17434 18366 17436
rect 18422 17434 18446 17436
rect 18284 17382 18286 17434
rect 18348 17382 18360 17434
rect 18422 17382 18424 17434
rect 18262 17380 18286 17382
rect 18342 17380 18366 17382
rect 18422 17380 18446 17382
rect 18206 17360 18502 17380
rect 18616 17202 18644 19071
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 19064 18828 19116 18834
rect 19064 18770 19116 18776
rect 18800 18426 18828 18770
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 19076 18154 19104 18770
rect 19168 18222 19196 19246
rect 19245 18352 19297 18358
rect 19245 18294 19297 18300
rect 19257 18278 19288 18294
rect 19156 18216 19208 18222
rect 19156 18158 19208 18164
rect 19064 18148 19116 18154
rect 19064 18090 19116 18096
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18708 16794 18736 17070
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18206 16348 18502 16368
rect 18262 16346 18286 16348
rect 18342 16346 18366 16348
rect 18422 16346 18446 16348
rect 18284 16294 18286 16346
rect 18348 16294 18360 16346
rect 18422 16294 18424 16346
rect 18262 16292 18286 16294
rect 18342 16292 18366 16294
rect 18422 16292 18446 16294
rect 18206 16272 18502 16292
rect 18708 16046 18736 16730
rect 18892 16658 18920 17614
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18984 17066 19012 17478
rect 19076 17338 19104 18090
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 18972 17060 19024 17066
rect 18972 17002 19024 17008
rect 18984 16726 19012 17002
rect 19064 16992 19116 16998
rect 19064 16934 19116 16940
rect 18972 16720 19024 16726
rect 18972 16662 19024 16668
rect 19076 16658 19104 16934
rect 18880 16652 18932 16658
rect 18880 16594 18932 16600
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18604 15972 18656 15978
rect 18604 15914 18656 15920
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17972 15026 18000 15302
rect 18206 15260 18502 15280
rect 18262 15258 18286 15260
rect 18342 15258 18366 15260
rect 18422 15258 18446 15260
rect 18284 15206 18286 15258
rect 18348 15206 18360 15258
rect 18422 15206 18424 15258
rect 18262 15204 18286 15206
rect 18342 15204 18366 15206
rect 18422 15204 18446 15206
rect 18206 15184 18502 15204
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17972 14498 18000 14962
rect 17880 14482 18000 14498
rect 18616 14482 18644 15914
rect 18708 14958 18736 15982
rect 18788 15564 18840 15570
rect 18788 15506 18840 15512
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18800 14890 18828 15506
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 17880 14476 18012 14482
rect 17880 14470 17960 14476
rect 17880 13870 17908 14470
rect 17960 14418 18012 14424
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18800 14414 18828 14826
rect 18892 14550 18920 16594
rect 19168 16250 19196 18158
rect 19260 18086 19288 18278
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19352 17898 19380 20334
rect 19628 19310 19656 20742
rect 19616 19304 19668 19310
rect 19616 19246 19668 19252
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19536 18358 19564 19110
rect 19524 18352 19576 18358
rect 19524 18294 19576 18300
rect 19536 18222 19564 18294
rect 19628 18290 19656 19246
rect 19904 19242 19932 21286
rect 19996 20466 20024 21422
rect 20180 21010 20208 22374
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 20168 21004 20220 21010
rect 20168 20946 20220 20952
rect 20628 20800 20680 20806
rect 20628 20742 20680 20748
rect 20640 20505 20668 20742
rect 20626 20496 20682 20505
rect 19984 20460 20036 20466
rect 20626 20431 20682 20440
rect 19984 20402 20036 20408
rect 20628 20324 20680 20330
rect 20628 20266 20680 20272
rect 20640 20058 20668 20266
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20824 19922 20852 22034
rect 21088 21480 21140 21486
rect 21088 21422 21140 21428
rect 21100 20602 21128 21422
rect 21180 21004 21232 21010
rect 21180 20946 21232 20952
rect 21088 20596 21140 20602
rect 21088 20538 21140 20544
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 19892 19236 19944 19242
rect 19892 19178 19944 19184
rect 20444 19236 20496 19242
rect 20444 19178 20496 19184
rect 19616 18284 19668 18290
rect 19616 18226 19668 18232
rect 19524 18216 19576 18222
rect 19524 18158 19576 18164
rect 19352 17870 19472 17898
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19352 17218 19380 17682
rect 19260 17202 19380 17218
rect 19248 17196 19380 17202
rect 19300 17190 19380 17196
rect 19248 17138 19300 17144
rect 19156 16244 19208 16250
rect 19156 16186 19208 16192
rect 18880 14544 18932 14550
rect 19260 14521 19288 17138
rect 19340 17128 19392 17134
rect 19444 17082 19472 17870
rect 20456 17746 20484 19178
rect 20720 18896 20772 18902
rect 20720 18838 20772 18844
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 20640 17785 20668 18158
rect 20732 18086 20760 18838
rect 20824 18170 20852 19858
rect 20824 18142 20944 18170
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20812 18080 20864 18086
rect 20812 18022 20864 18028
rect 20626 17776 20682 17785
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20444 17740 20496 17746
rect 20626 17711 20682 17720
rect 20444 17682 20496 17688
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19628 17202 19656 17478
rect 20272 17338 20300 17682
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19392 17076 19472 17082
rect 19340 17070 19472 17076
rect 19352 17054 19472 17070
rect 20628 17060 20680 17066
rect 19352 14958 19380 17054
rect 20628 17002 20680 17008
rect 20640 16794 20668 17002
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20732 16250 20760 18022
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19996 15026 20024 15846
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 18880 14486 18932 14492
rect 19246 14512 19302 14521
rect 19246 14447 19302 14456
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 17960 14340 18012 14346
rect 17960 14282 18012 14288
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17972 13462 18000 14282
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 18064 13870 18092 14214
rect 18206 14172 18502 14192
rect 18262 14170 18286 14172
rect 18342 14170 18366 14172
rect 18422 14170 18446 14172
rect 18284 14118 18286 14170
rect 18348 14118 18360 14170
rect 18422 14118 18424 14170
rect 18262 14116 18286 14118
rect 18342 14116 18366 14118
rect 18422 14116 18446 14118
rect 18206 14096 18502 14116
rect 19260 13938 19288 14447
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18604 13728 18656 13734
rect 18604 13670 18656 13676
rect 17960 13456 18012 13462
rect 17960 13398 18012 13404
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17972 12850 18000 13262
rect 18206 13084 18502 13104
rect 18262 13082 18286 13084
rect 18342 13082 18366 13084
rect 18422 13082 18446 13084
rect 18284 13030 18286 13082
rect 18348 13030 18360 13082
rect 18422 13030 18424 13082
rect 18262 13028 18286 13030
rect 18342 13028 18366 13030
rect 18422 13028 18446 13030
rect 18206 13008 18502 13028
rect 18616 12850 18644 13670
rect 19352 13326 19380 14894
rect 19616 14884 19668 14890
rect 19616 14826 19668 14832
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19536 13870 19564 14418
rect 19628 14074 19656 14826
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19720 13870 19748 14758
rect 19996 14618 20024 14962
rect 20628 14884 20680 14890
rect 20628 14826 20680 14832
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20272 14618 20300 14758
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19708 13864 19760 13870
rect 19708 13806 19760 13812
rect 20272 13802 20300 14418
rect 20640 14074 20668 14826
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20720 13864 20772 13870
rect 20640 13812 20720 13818
rect 20640 13806 20772 13812
rect 20260 13796 20312 13802
rect 20260 13738 20312 13744
rect 20640 13790 20760 13806
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 20272 12850 20300 13738
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 19996 12442 20024 12650
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 20640 12306 20668 13790
rect 20824 12306 20852 18022
rect 20916 16658 20944 18142
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20916 16130 20944 16594
rect 20916 16102 21036 16130
rect 20904 16040 20956 16046
rect 20904 15982 20956 15988
rect 20916 15706 20944 15982
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 21008 13870 21036 16102
rect 21086 15736 21142 15745
rect 21086 15671 21142 15680
rect 21100 15570 21128 15671
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 21086 13016 21142 13025
rect 21086 12951 21142 12960
rect 21100 12782 21128 12951
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 18206 11996 18502 12016
rect 18262 11994 18286 11996
rect 18342 11994 18366 11996
rect 18422 11994 18446 11996
rect 18284 11942 18286 11994
rect 18348 11942 18360 11994
rect 18422 11942 18424 11994
rect 18262 11940 18286 11942
rect 18342 11940 18366 11942
rect 18422 11940 18446 11942
rect 18206 11920 18502 11940
rect 20732 11694 20760 12038
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20732 11286 20760 11494
rect 20720 11280 20772 11286
rect 20720 11222 20772 11228
rect 18206 10908 18502 10928
rect 18262 10906 18286 10908
rect 18342 10906 18366 10908
rect 18422 10906 18446 10908
rect 18284 10854 18286 10906
rect 18348 10854 18360 10906
rect 18422 10854 18424 10906
rect 18262 10852 18286 10854
rect 18342 10852 18366 10854
rect 18422 10852 18446 10854
rect 18206 10832 18502 10852
rect 20824 10810 20852 11698
rect 20916 11694 20944 12582
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 20904 10600 20956 10606
rect 20904 10542 20956 10548
rect 20916 10266 20944 10542
rect 21086 10296 21142 10305
rect 20904 10260 20956 10266
rect 21086 10231 21142 10240
rect 20904 10202 20956 10208
rect 21100 10130 21128 10231
rect 21088 10124 21140 10130
rect 21088 10066 21140 10072
rect 18206 9820 18502 9840
rect 18262 9818 18286 9820
rect 18342 9818 18366 9820
rect 18422 9818 18446 9820
rect 18284 9766 18286 9818
rect 18348 9766 18360 9818
rect 18422 9766 18424 9818
rect 18262 9764 18286 9766
rect 18342 9764 18366 9766
rect 18422 9764 18446 9766
rect 18206 9744 18502 9764
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 18206 8732 18502 8752
rect 18262 8730 18286 8732
rect 18342 8730 18366 8732
rect 18422 8730 18446 8732
rect 18284 8678 18286 8730
rect 18348 8678 18360 8730
rect 18422 8678 18424 8730
rect 18262 8676 18286 8678
rect 18342 8676 18366 8678
rect 18422 8676 18446 8678
rect 18206 8656 18502 8676
rect 20640 8634 20668 8910
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20732 8498 20760 8774
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20904 8424 20956 8430
rect 20904 8366 20956 8372
rect 20916 8090 20944 8366
rect 21086 8256 21142 8265
rect 21086 8191 21142 8200
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 21100 7954 21128 8191
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 21088 7948 21140 7954
rect 21088 7890 21140 7896
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 17500 7268 17552 7274
rect 17500 7210 17552 7216
rect 14756 7100 15052 7120
rect 14812 7098 14836 7100
rect 14892 7098 14916 7100
rect 14972 7098 14996 7100
rect 14834 7046 14836 7098
rect 14898 7046 14910 7098
rect 14972 7046 14974 7098
rect 14812 7044 14836 7046
rect 14892 7044 14916 7046
rect 14972 7044 14996 7046
rect 14756 7024 15052 7044
rect 14660 6886 15148 6914
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13188 6338 13216 6394
rect 13188 6310 13308 6338
rect 13280 6254 13308 6310
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14660 5914 14688 6054
rect 14756 6012 15052 6032
rect 14812 6010 14836 6012
rect 14892 6010 14916 6012
rect 14972 6010 14996 6012
rect 14834 5958 14836 6010
rect 14898 5958 14910 6010
rect 14972 5958 14974 6010
rect 14812 5956 14836 5958
rect 14892 5956 14916 5958
rect 14972 5956 14996 5958
rect 14756 5936 15052 5956
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14756 4924 15052 4944
rect 14812 4922 14836 4924
rect 14892 4922 14916 4924
rect 14972 4922 14996 4924
rect 14834 4870 14836 4922
rect 14898 4870 14910 4922
rect 14972 4870 14974 4922
rect 14812 4868 14836 4870
rect 14892 4868 14916 4870
rect 14972 4868 14996 4870
rect 14756 4848 15052 4868
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13280 4282 13308 4626
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13280 3738 13308 4218
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13648 3534 13676 4014
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13924 3126 13952 3946
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 13360 2916 13412 2922
rect 13360 2858 13412 2864
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 11992 2746 12112 2774
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 1860 2576 1912 2582
rect 1860 2518 1912 2524
rect 8760 2576 8812 2582
rect 8760 2518 8812 2524
rect 480 2508 532 2514
rect 480 2450 532 2456
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 492 800 520 2450
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 1872 800 1900 2314
rect 3712 800 3740 2450
rect 4406 2204 4702 2224
rect 4462 2202 4486 2204
rect 4542 2202 4566 2204
rect 4622 2202 4646 2204
rect 4484 2150 4486 2202
rect 4548 2150 4560 2202
rect 4622 2150 4624 2202
rect 4462 2148 4486 2150
rect 4542 2148 4566 2150
rect 4622 2148 4646 2150
rect 4406 2128 4702 2148
rect 5552 800 5580 2450
rect 6932 800 6960 2450
rect 8772 800 8800 2518
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 10612 800 10640 2450
rect 11306 2204 11602 2224
rect 11362 2202 11386 2204
rect 11442 2202 11466 2204
rect 11522 2202 11546 2204
rect 11384 2150 11386 2202
rect 11448 2150 11460 2202
rect 11522 2150 11524 2202
rect 11362 2148 11386 2150
rect 11442 2148 11466 2150
rect 11522 2148 11546 2150
rect 11306 2128 11602 2148
rect 11992 800 12020 2746
rect 13280 2514 13308 2790
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 13372 2310 13400 2858
rect 13924 2650 13952 3062
rect 14108 2922 14136 4082
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 14200 3602 14228 3878
rect 14756 3836 15052 3856
rect 14812 3834 14836 3836
rect 14892 3834 14916 3836
rect 14972 3834 14996 3836
rect 14834 3782 14836 3834
rect 14898 3782 14910 3834
rect 14972 3782 14974 3834
rect 14812 3780 14836 3782
rect 14892 3780 14916 3782
rect 14972 3780 14996 3782
rect 14756 3760 15052 3780
rect 15120 3738 15148 6886
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15672 5234 15700 5646
rect 15764 5370 15792 5646
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 16132 5166 16160 6190
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 15856 4554 15884 5102
rect 16224 4622 16252 6258
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16500 5710 16528 6190
rect 17512 6186 17540 7210
rect 16580 6180 16632 6186
rect 16580 6122 16632 6128
rect 17500 6180 17552 6186
rect 17500 6122 17552 6128
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16396 5636 16448 5642
rect 16396 5578 16448 5584
rect 16408 4826 16436 5578
rect 16592 5098 16620 6122
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16684 4690 16712 5102
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17420 4690 17448 4966
rect 17880 4758 17908 5646
rect 17868 4752 17920 4758
rect 17868 4694 17920 4700
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 15856 4282 15884 4490
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 16224 4078 16252 4558
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15396 3194 15424 3470
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15396 3058 15424 3130
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 14096 2916 14148 2922
rect 14096 2858 14148 2864
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 14108 2514 14136 2858
rect 14756 2748 15052 2768
rect 14812 2746 14836 2748
rect 14892 2746 14916 2748
rect 14972 2746 14996 2748
rect 14834 2694 14836 2746
rect 14898 2694 14910 2746
rect 14972 2694 14974 2746
rect 14812 2692 14836 2694
rect 14892 2692 14916 2694
rect 14972 2692 14996 2694
rect 14756 2672 15052 2692
rect 15488 2582 15516 4014
rect 17236 3126 17264 4626
rect 17972 3194 18000 7890
rect 18206 7644 18502 7664
rect 18262 7642 18286 7644
rect 18342 7642 18366 7644
rect 18422 7642 18446 7644
rect 18284 7590 18286 7642
rect 18348 7590 18360 7642
rect 18422 7590 18424 7642
rect 18262 7588 18286 7590
rect 18342 7588 18366 7590
rect 18422 7588 18446 7590
rect 18206 7568 18502 7588
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 18206 6556 18502 6576
rect 18262 6554 18286 6556
rect 18342 6554 18366 6556
rect 18422 6554 18446 6556
rect 18284 6502 18286 6554
rect 18348 6502 18360 6554
rect 18422 6502 18424 6554
rect 18262 6500 18286 6502
rect 18342 6500 18366 6502
rect 18422 6500 18446 6502
rect 18206 6480 18502 6500
rect 19720 6458 19748 6802
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20640 6458 20668 6734
rect 21192 6730 21220 20946
rect 21376 9042 21404 22374
rect 21652 22098 21680 24323
rect 21640 22092 21692 22098
rect 21640 22034 21692 22040
rect 21364 9036 21416 9042
rect 21364 8978 21416 8984
rect 21180 6724 21232 6730
rect 21180 6666 21232 6672
rect 19708 6452 19760 6458
rect 19708 6394 19760 6400
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 19720 6322 19748 6394
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 18064 5914 18092 6258
rect 18604 6180 18656 6186
rect 18604 6122 18656 6128
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 18064 5370 18092 5714
rect 18206 5468 18502 5488
rect 18262 5466 18286 5468
rect 18342 5466 18366 5468
rect 18422 5466 18446 5468
rect 18284 5414 18286 5466
rect 18348 5414 18360 5466
rect 18422 5414 18424 5466
rect 18262 5412 18286 5414
rect 18342 5412 18366 5414
rect 18422 5412 18446 5414
rect 18206 5392 18502 5412
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 18616 5098 18644 6122
rect 19720 5370 19748 6258
rect 20996 6248 21048 6254
rect 20996 6190 21048 6196
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 20916 5370 20944 5714
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 18156 4690 18184 5034
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 18206 4380 18502 4400
rect 18262 4378 18286 4380
rect 18342 4378 18366 4380
rect 18422 4378 18446 4380
rect 18284 4326 18286 4378
rect 18348 4326 18360 4378
rect 18422 4326 18424 4378
rect 18262 4324 18286 4326
rect 18342 4324 18366 4326
rect 18422 4324 18446 4326
rect 18206 4304 18502 4324
rect 19260 4078 19288 5170
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 18206 3292 18502 3312
rect 18262 3290 18286 3292
rect 18342 3290 18366 3292
rect 18422 3290 18446 3292
rect 18284 3238 18286 3290
rect 18348 3238 18360 3290
rect 18422 3238 18424 3290
rect 18262 3236 18286 3238
rect 18342 3236 18366 3238
rect 18422 3236 18446 3238
rect 18206 3216 18502 3236
rect 20732 3194 20760 3538
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 20720 3188 20772 3194
rect 20720 3130 20772 3136
rect 17224 3120 17276 3126
rect 17224 3062 17276 3068
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 18236 2984 18288 2990
rect 18236 2926 18288 2932
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 16132 2650 16160 2926
rect 17500 2916 17552 2922
rect 17500 2858 17552 2864
rect 17512 2650 17540 2858
rect 18248 2650 18276 2926
rect 20088 2825 20116 2926
rect 20074 2816 20130 2825
rect 20074 2751 20130 2760
rect 16120 2644 16172 2650
rect 16120 2586 16172 2592
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 18236 2644 18288 2650
rect 18236 2586 18288 2592
rect 20916 2582 20944 3878
rect 21008 3738 21036 6190
rect 21086 5536 21142 5545
rect 21086 5471 21142 5480
rect 21100 5166 21128 5471
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 20996 3732 21048 3738
rect 20996 3674 21048 3680
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 15476 2576 15528 2582
rect 15476 2518 15528 2524
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 15660 2508 15712 2514
rect 15660 2450 15712 2456
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 13740 1442 13768 2382
rect 13740 1414 13860 1442
rect 13832 800 13860 1414
rect 15672 800 15700 2450
rect 17052 800 17080 2450
rect 18206 2204 18502 2224
rect 18262 2202 18286 2204
rect 18342 2202 18366 2204
rect 18422 2202 18446 2204
rect 18284 2150 18286 2202
rect 18348 2150 18360 2202
rect 18422 2150 18424 2202
rect 18262 2148 18286 2150
rect 18342 2148 18366 2150
rect 18422 2148 18446 2150
rect 18206 2128 18502 2148
rect 18892 800 18920 2450
rect 20720 2372 20772 2378
rect 20720 2314 20772 2320
rect 20732 800 20760 2314
rect 22112 800 22140 3538
rect 478 0 534 800
rect 1858 0 1914 800
rect 3698 0 3754 800
rect 5538 0 5594 800
rect 6918 0 6974 800
rect 8758 0 8814 800
rect 10598 0 10654 800
rect 11978 0 12034 800
rect 13818 0 13874 800
rect 15658 0 15714 800
rect 17038 0 17094 800
rect 18878 0 18934 800
rect 20718 0 20774 800
rect 22098 0 22154 800
<< via2 >>
rect 1490 23160 1546 23216
rect 4406 22874 4462 22876
rect 4486 22874 4542 22876
rect 4566 22874 4622 22876
rect 4646 22874 4702 22876
rect 4406 22822 4432 22874
rect 4432 22822 4462 22874
rect 4486 22822 4496 22874
rect 4496 22822 4542 22874
rect 4566 22822 4612 22874
rect 4612 22822 4622 22874
rect 4646 22822 4676 22874
rect 4676 22822 4702 22874
rect 4406 22820 4462 22822
rect 4486 22820 4542 22822
rect 4566 22820 4622 22822
rect 4646 22820 4702 22822
rect 11306 22874 11362 22876
rect 11386 22874 11442 22876
rect 11466 22874 11522 22876
rect 11546 22874 11602 22876
rect 11306 22822 11332 22874
rect 11332 22822 11362 22874
rect 11386 22822 11396 22874
rect 11396 22822 11442 22874
rect 11466 22822 11512 22874
rect 11512 22822 11522 22874
rect 11546 22822 11576 22874
rect 11576 22822 11602 22874
rect 11306 22820 11362 22822
rect 11386 22820 11442 22822
rect 11466 22820 11522 22822
rect 11546 22820 11602 22822
rect 18206 22874 18262 22876
rect 18286 22874 18342 22876
rect 18366 22874 18422 22876
rect 18446 22874 18502 22876
rect 18206 22822 18232 22874
rect 18232 22822 18262 22874
rect 18286 22822 18296 22874
rect 18296 22822 18342 22874
rect 18366 22822 18412 22874
rect 18412 22822 18422 22874
rect 18446 22822 18476 22874
rect 18476 22822 18502 22874
rect 18206 22820 18262 22822
rect 18286 22820 18342 22822
rect 18366 22820 18422 22822
rect 18446 22820 18502 22822
rect 21086 23160 21142 23216
rect 1398 20440 1454 20496
rect 1398 17740 1454 17776
rect 1398 17720 1400 17740
rect 1400 17720 1452 17740
rect 1452 17720 1454 17740
rect 4406 21786 4462 21788
rect 4486 21786 4542 21788
rect 4566 21786 4622 21788
rect 4646 21786 4702 21788
rect 4406 21734 4432 21786
rect 4432 21734 4462 21786
rect 4486 21734 4496 21786
rect 4496 21734 4542 21786
rect 4566 21734 4612 21786
rect 4612 21734 4622 21786
rect 4646 21734 4676 21786
rect 4676 21734 4702 21786
rect 4406 21732 4462 21734
rect 4486 21732 4542 21734
rect 4566 21732 4622 21734
rect 4646 21732 4702 21734
rect 7856 22330 7912 22332
rect 7936 22330 7992 22332
rect 8016 22330 8072 22332
rect 8096 22330 8152 22332
rect 7856 22278 7882 22330
rect 7882 22278 7912 22330
rect 7936 22278 7946 22330
rect 7946 22278 7992 22330
rect 8016 22278 8062 22330
rect 8062 22278 8072 22330
rect 8096 22278 8126 22330
rect 8126 22278 8152 22330
rect 7856 22276 7912 22278
rect 7936 22276 7992 22278
rect 8016 22276 8072 22278
rect 8096 22276 8152 22278
rect 1398 15680 1454 15736
rect 1490 12980 1546 13016
rect 1490 12960 1492 12980
rect 1492 12960 1544 12980
rect 1544 12960 1546 12980
rect 1490 10260 1546 10296
rect 1490 10240 1492 10260
rect 1492 10240 1544 10260
rect 1544 10240 1546 10260
rect 1398 8200 1454 8256
rect 1490 5516 1492 5536
rect 1492 5516 1544 5536
rect 1544 5516 1546 5536
rect 1490 5480 1546 5516
rect 1398 2760 1454 2816
rect 4406 20698 4462 20700
rect 4486 20698 4542 20700
rect 4566 20698 4622 20700
rect 4646 20698 4702 20700
rect 4406 20646 4432 20698
rect 4432 20646 4462 20698
rect 4486 20646 4496 20698
rect 4496 20646 4542 20698
rect 4566 20646 4612 20698
rect 4612 20646 4622 20698
rect 4646 20646 4676 20698
rect 4676 20646 4702 20698
rect 4406 20644 4462 20646
rect 4486 20644 4542 20646
rect 4566 20644 4622 20646
rect 4646 20644 4702 20646
rect 4406 19610 4462 19612
rect 4486 19610 4542 19612
rect 4566 19610 4622 19612
rect 4646 19610 4702 19612
rect 4406 19558 4432 19610
rect 4432 19558 4462 19610
rect 4486 19558 4496 19610
rect 4496 19558 4542 19610
rect 4566 19558 4612 19610
rect 4612 19558 4622 19610
rect 4646 19558 4676 19610
rect 4676 19558 4702 19610
rect 4406 19556 4462 19558
rect 4486 19556 4542 19558
rect 4566 19556 4622 19558
rect 4646 19556 4702 19558
rect 4406 18522 4462 18524
rect 4486 18522 4542 18524
rect 4566 18522 4622 18524
rect 4646 18522 4702 18524
rect 4406 18470 4432 18522
rect 4432 18470 4462 18522
rect 4486 18470 4496 18522
rect 4496 18470 4542 18522
rect 4566 18470 4612 18522
rect 4612 18470 4622 18522
rect 4646 18470 4676 18522
rect 4676 18470 4702 18522
rect 4406 18468 4462 18470
rect 4486 18468 4542 18470
rect 4566 18468 4622 18470
rect 4646 18468 4702 18470
rect 4406 17434 4462 17436
rect 4486 17434 4542 17436
rect 4566 17434 4622 17436
rect 4646 17434 4702 17436
rect 4406 17382 4432 17434
rect 4432 17382 4462 17434
rect 4486 17382 4496 17434
rect 4496 17382 4542 17434
rect 4566 17382 4612 17434
rect 4612 17382 4622 17434
rect 4646 17382 4676 17434
rect 4676 17382 4702 17434
rect 4406 17380 4462 17382
rect 4486 17380 4542 17382
rect 4566 17380 4622 17382
rect 4646 17380 4702 17382
rect 4406 16346 4462 16348
rect 4486 16346 4542 16348
rect 4566 16346 4622 16348
rect 4646 16346 4702 16348
rect 4406 16294 4432 16346
rect 4432 16294 4462 16346
rect 4486 16294 4496 16346
rect 4496 16294 4542 16346
rect 4566 16294 4612 16346
rect 4612 16294 4622 16346
rect 4646 16294 4676 16346
rect 4676 16294 4702 16346
rect 4406 16292 4462 16294
rect 4486 16292 4542 16294
rect 4566 16292 4622 16294
rect 4646 16292 4702 16294
rect 4406 15258 4462 15260
rect 4486 15258 4542 15260
rect 4566 15258 4622 15260
rect 4646 15258 4702 15260
rect 4406 15206 4432 15258
rect 4432 15206 4462 15258
rect 4486 15206 4496 15258
rect 4496 15206 4542 15258
rect 4566 15206 4612 15258
rect 4612 15206 4622 15258
rect 4646 15206 4676 15258
rect 4676 15206 4702 15258
rect 4406 15204 4462 15206
rect 4486 15204 4542 15206
rect 4566 15204 4622 15206
rect 4646 15204 4702 15206
rect 4406 14170 4462 14172
rect 4486 14170 4542 14172
rect 4566 14170 4622 14172
rect 4646 14170 4702 14172
rect 4406 14118 4432 14170
rect 4432 14118 4462 14170
rect 4486 14118 4496 14170
rect 4496 14118 4542 14170
rect 4566 14118 4612 14170
rect 4612 14118 4622 14170
rect 4646 14118 4676 14170
rect 4676 14118 4702 14170
rect 4406 14116 4462 14118
rect 4486 14116 4542 14118
rect 4566 14116 4622 14118
rect 4646 14116 4702 14118
rect 4406 13082 4462 13084
rect 4486 13082 4542 13084
rect 4566 13082 4622 13084
rect 4646 13082 4702 13084
rect 4406 13030 4432 13082
rect 4432 13030 4462 13082
rect 4486 13030 4496 13082
rect 4496 13030 4542 13082
rect 4566 13030 4612 13082
rect 4612 13030 4622 13082
rect 4646 13030 4676 13082
rect 4676 13030 4702 13082
rect 4406 13028 4462 13030
rect 4486 13028 4542 13030
rect 4566 13028 4622 13030
rect 4646 13028 4702 13030
rect 4406 11994 4462 11996
rect 4486 11994 4542 11996
rect 4566 11994 4622 11996
rect 4646 11994 4702 11996
rect 4406 11942 4432 11994
rect 4432 11942 4462 11994
rect 4486 11942 4496 11994
rect 4496 11942 4542 11994
rect 4566 11942 4612 11994
rect 4612 11942 4622 11994
rect 4646 11942 4676 11994
rect 4676 11942 4702 11994
rect 4406 11940 4462 11942
rect 4486 11940 4542 11942
rect 4566 11940 4622 11942
rect 4646 11940 4702 11942
rect 4406 10906 4462 10908
rect 4486 10906 4542 10908
rect 4566 10906 4622 10908
rect 4646 10906 4702 10908
rect 4406 10854 4432 10906
rect 4432 10854 4462 10906
rect 4486 10854 4496 10906
rect 4496 10854 4542 10906
rect 4566 10854 4612 10906
rect 4612 10854 4622 10906
rect 4646 10854 4676 10906
rect 4676 10854 4702 10906
rect 4406 10852 4462 10854
rect 4486 10852 4542 10854
rect 4566 10852 4622 10854
rect 4646 10852 4702 10854
rect 4406 9818 4462 9820
rect 4486 9818 4542 9820
rect 4566 9818 4622 9820
rect 4646 9818 4702 9820
rect 4406 9766 4432 9818
rect 4432 9766 4462 9818
rect 4486 9766 4496 9818
rect 4496 9766 4542 9818
rect 4566 9766 4612 9818
rect 4612 9766 4622 9818
rect 4646 9766 4676 9818
rect 4676 9766 4702 9818
rect 4406 9764 4462 9766
rect 4486 9764 4542 9766
rect 4566 9764 4622 9766
rect 4646 9764 4702 9766
rect 4406 8730 4462 8732
rect 4486 8730 4542 8732
rect 4566 8730 4622 8732
rect 4646 8730 4702 8732
rect 4406 8678 4432 8730
rect 4432 8678 4462 8730
rect 4486 8678 4496 8730
rect 4496 8678 4542 8730
rect 4566 8678 4612 8730
rect 4612 8678 4622 8730
rect 4646 8678 4676 8730
rect 4676 8678 4702 8730
rect 4406 8676 4462 8678
rect 4486 8676 4542 8678
rect 4566 8676 4622 8678
rect 4646 8676 4702 8678
rect 4406 7642 4462 7644
rect 4486 7642 4542 7644
rect 4566 7642 4622 7644
rect 4646 7642 4702 7644
rect 4406 7590 4432 7642
rect 4432 7590 4462 7642
rect 4486 7590 4496 7642
rect 4496 7590 4542 7642
rect 4566 7590 4612 7642
rect 4612 7590 4622 7642
rect 4646 7590 4676 7642
rect 4676 7590 4702 7642
rect 4406 7588 4462 7590
rect 4486 7588 4542 7590
rect 4566 7588 4622 7590
rect 4646 7588 4702 7590
rect 7856 21242 7912 21244
rect 7936 21242 7992 21244
rect 8016 21242 8072 21244
rect 8096 21242 8152 21244
rect 7856 21190 7882 21242
rect 7882 21190 7912 21242
rect 7936 21190 7946 21242
rect 7946 21190 7992 21242
rect 8016 21190 8062 21242
rect 8062 21190 8072 21242
rect 8096 21190 8126 21242
rect 8126 21190 8152 21242
rect 7856 21188 7912 21190
rect 7936 21188 7992 21190
rect 8016 21188 8072 21190
rect 8096 21188 8152 21190
rect 7856 20154 7912 20156
rect 7936 20154 7992 20156
rect 8016 20154 8072 20156
rect 8096 20154 8152 20156
rect 7856 20102 7882 20154
rect 7882 20102 7912 20154
rect 7936 20102 7946 20154
rect 7946 20102 7992 20154
rect 8016 20102 8062 20154
rect 8062 20102 8072 20154
rect 8096 20102 8126 20154
rect 8126 20102 8152 20154
rect 7856 20100 7912 20102
rect 7936 20100 7992 20102
rect 8016 20100 8072 20102
rect 8096 20100 8152 20102
rect 7856 19066 7912 19068
rect 7936 19066 7992 19068
rect 8016 19066 8072 19068
rect 8096 19066 8152 19068
rect 7856 19014 7882 19066
rect 7882 19014 7912 19066
rect 7936 19014 7946 19066
rect 7946 19014 7992 19066
rect 8016 19014 8062 19066
rect 8062 19014 8072 19066
rect 8096 19014 8126 19066
rect 8126 19014 8152 19066
rect 7856 19012 7912 19014
rect 7936 19012 7992 19014
rect 8016 19012 8072 19014
rect 8096 19012 8152 19014
rect 7856 17978 7912 17980
rect 7936 17978 7992 17980
rect 8016 17978 8072 17980
rect 8096 17978 8152 17980
rect 7856 17926 7882 17978
rect 7882 17926 7912 17978
rect 7936 17926 7946 17978
rect 7946 17926 7992 17978
rect 8016 17926 8062 17978
rect 8062 17926 8072 17978
rect 8096 17926 8126 17978
rect 8126 17926 8152 17978
rect 7856 17924 7912 17926
rect 7936 17924 7992 17926
rect 8016 17924 8072 17926
rect 8096 17924 8152 17926
rect 7856 16890 7912 16892
rect 7936 16890 7992 16892
rect 8016 16890 8072 16892
rect 8096 16890 8152 16892
rect 7856 16838 7882 16890
rect 7882 16838 7912 16890
rect 7936 16838 7946 16890
rect 7946 16838 7992 16890
rect 8016 16838 8062 16890
rect 8062 16838 8072 16890
rect 8096 16838 8126 16890
rect 8126 16838 8152 16890
rect 7856 16836 7912 16838
rect 7936 16836 7992 16838
rect 8016 16836 8072 16838
rect 8096 16836 8152 16838
rect 7856 15802 7912 15804
rect 7936 15802 7992 15804
rect 8016 15802 8072 15804
rect 8096 15802 8152 15804
rect 7856 15750 7882 15802
rect 7882 15750 7912 15802
rect 7936 15750 7946 15802
rect 7946 15750 7992 15802
rect 8016 15750 8062 15802
rect 8062 15750 8072 15802
rect 8096 15750 8126 15802
rect 8126 15750 8152 15802
rect 7856 15748 7912 15750
rect 7936 15748 7992 15750
rect 8016 15748 8072 15750
rect 8096 15748 8152 15750
rect 7856 14714 7912 14716
rect 7936 14714 7992 14716
rect 8016 14714 8072 14716
rect 8096 14714 8152 14716
rect 7856 14662 7882 14714
rect 7882 14662 7912 14714
rect 7936 14662 7946 14714
rect 7946 14662 7992 14714
rect 8016 14662 8062 14714
rect 8062 14662 8072 14714
rect 8096 14662 8126 14714
rect 8126 14662 8152 14714
rect 7856 14660 7912 14662
rect 7936 14660 7992 14662
rect 8016 14660 8072 14662
rect 8096 14660 8152 14662
rect 7856 13626 7912 13628
rect 7936 13626 7992 13628
rect 8016 13626 8072 13628
rect 8096 13626 8152 13628
rect 7856 13574 7882 13626
rect 7882 13574 7912 13626
rect 7936 13574 7946 13626
rect 7946 13574 7992 13626
rect 8016 13574 8062 13626
rect 8062 13574 8072 13626
rect 8096 13574 8126 13626
rect 8126 13574 8152 13626
rect 7856 13572 7912 13574
rect 7936 13572 7992 13574
rect 8016 13572 8072 13574
rect 8096 13572 8152 13574
rect 4406 6554 4462 6556
rect 4486 6554 4542 6556
rect 4566 6554 4622 6556
rect 4646 6554 4702 6556
rect 4406 6502 4432 6554
rect 4432 6502 4462 6554
rect 4486 6502 4496 6554
rect 4496 6502 4542 6554
rect 4566 6502 4612 6554
rect 4612 6502 4622 6554
rect 4646 6502 4676 6554
rect 4676 6502 4702 6554
rect 4406 6500 4462 6502
rect 4486 6500 4542 6502
rect 4566 6500 4622 6502
rect 4646 6500 4702 6502
rect 4406 5466 4462 5468
rect 4486 5466 4542 5468
rect 4566 5466 4622 5468
rect 4646 5466 4702 5468
rect 4406 5414 4432 5466
rect 4432 5414 4462 5466
rect 4486 5414 4496 5466
rect 4496 5414 4542 5466
rect 4566 5414 4612 5466
rect 4612 5414 4622 5466
rect 4646 5414 4676 5466
rect 4676 5414 4702 5466
rect 4406 5412 4462 5414
rect 4486 5412 4542 5414
rect 4566 5412 4622 5414
rect 4646 5412 4702 5414
rect 4406 4378 4462 4380
rect 4486 4378 4542 4380
rect 4566 4378 4622 4380
rect 4646 4378 4702 4380
rect 4406 4326 4432 4378
rect 4432 4326 4462 4378
rect 4486 4326 4496 4378
rect 4496 4326 4542 4378
rect 4566 4326 4612 4378
rect 4612 4326 4622 4378
rect 4646 4326 4676 4378
rect 4676 4326 4702 4378
rect 4406 4324 4462 4326
rect 4486 4324 4542 4326
rect 4566 4324 4622 4326
rect 4646 4324 4702 4326
rect 4406 3290 4462 3292
rect 4486 3290 4542 3292
rect 4566 3290 4622 3292
rect 4646 3290 4702 3292
rect 4406 3238 4432 3290
rect 4432 3238 4462 3290
rect 4486 3238 4496 3290
rect 4496 3238 4542 3290
rect 4566 3238 4612 3290
rect 4612 3238 4622 3290
rect 4646 3238 4676 3290
rect 4676 3238 4702 3290
rect 4406 3236 4462 3238
rect 4486 3236 4542 3238
rect 4566 3236 4622 3238
rect 4646 3236 4702 3238
rect 14756 22330 14812 22332
rect 14836 22330 14892 22332
rect 14916 22330 14972 22332
rect 14996 22330 15052 22332
rect 14756 22278 14782 22330
rect 14782 22278 14812 22330
rect 14836 22278 14846 22330
rect 14846 22278 14892 22330
rect 14916 22278 14962 22330
rect 14962 22278 14972 22330
rect 14996 22278 15026 22330
rect 15026 22278 15052 22330
rect 14756 22276 14812 22278
rect 14836 22276 14892 22278
rect 14916 22276 14972 22278
rect 14996 22276 15052 22278
rect 11306 21786 11362 21788
rect 11386 21786 11442 21788
rect 11466 21786 11522 21788
rect 11546 21786 11602 21788
rect 11306 21734 11332 21786
rect 11332 21734 11362 21786
rect 11386 21734 11396 21786
rect 11396 21734 11442 21786
rect 11466 21734 11512 21786
rect 11512 21734 11522 21786
rect 11546 21734 11576 21786
rect 11576 21734 11602 21786
rect 11306 21732 11362 21734
rect 11386 21732 11442 21734
rect 11466 21732 11522 21734
rect 11546 21732 11602 21734
rect 11306 20698 11362 20700
rect 11386 20698 11442 20700
rect 11466 20698 11522 20700
rect 11546 20698 11602 20700
rect 11306 20646 11332 20698
rect 11332 20646 11362 20698
rect 11386 20646 11396 20698
rect 11396 20646 11442 20698
rect 11466 20646 11512 20698
rect 11512 20646 11522 20698
rect 11546 20646 11576 20698
rect 11576 20646 11602 20698
rect 11306 20644 11362 20646
rect 11386 20644 11442 20646
rect 11466 20644 11522 20646
rect 11546 20644 11602 20646
rect 11306 19610 11362 19612
rect 11386 19610 11442 19612
rect 11466 19610 11522 19612
rect 11546 19610 11602 19612
rect 11306 19558 11332 19610
rect 11332 19558 11362 19610
rect 11386 19558 11396 19610
rect 11396 19558 11442 19610
rect 11466 19558 11512 19610
rect 11512 19558 11522 19610
rect 11546 19558 11576 19610
rect 11576 19558 11602 19610
rect 11306 19556 11362 19558
rect 11386 19556 11442 19558
rect 11466 19556 11522 19558
rect 11546 19556 11602 19558
rect 11306 18522 11362 18524
rect 11386 18522 11442 18524
rect 11466 18522 11522 18524
rect 11546 18522 11602 18524
rect 11306 18470 11332 18522
rect 11332 18470 11362 18522
rect 11386 18470 11396 18522
rect 11396 18470 11442 18522
rect 11466 18470 11512 18522
rect 11512 18470 11522 18522
rect 11546 18470 11576 18522
rect 11576 18470 11602 18522
rect 11306 18468 11362 18470
rect 11386 18468 11442 18470
rect 11466 18468 11522 18470
rect 11546 18468 11602 18470
rect 12622 19372 12678 19408
rect 12622 19352 12624 19372
rect 12624 19352 12676 19372
rect 12676 19352 12678 19372
rect 11306 17434 11362 17436
rect 11386 17434 11442 17436
rect 11466 17434 11522 17436
rect 11546 17434 11602 17436
rect 11306 17382 11332 17434
rect 11332 17382 11362 17434
rect 11386 17382 11396 17434
rect 11396 17382 11442 17434
rect 11466 17382 11512 17434
rect 11512 17382 11522 17434
rect 11546 17382 11576 17434
rect 11576 17382 11602 17434
rect 11306 17380 11362 17382
rect 11386 17380 11442 17382
rect 11466 17380 11522 17382
rect 11546 17380 11602 17382
rect 11306 16346 11362 16348
rect 11386 16346 11442 16348
rect 11466 16346 11522 16348
rect 11546 16346 11602 16348
rect 11306 16294 11332 16346
rect 11332 16294 11362 16346
rect 11386 16294 11396 16346
rect 11396 16294 11442 16346
rect 11466 16294 11512 16346
rect 11512 16294 11522 16346
rect 11546 16294 11576 16346
rect 11576 16294 11602 16346
rect 11306 16292 11362 16294
rect 11386 16292 11442 16294
rect 11466 16292 11522 16294
rect 11546 16292 11602 16294
rect 11306 15258 11362 15260
rect 11386 15258 11442 15260
rect 11466 15258 11522 15260
rect 11546 15258 11602 15260
rect 11306 15206 11332 15258
rect 11332 15206 11362 15258
rect 11386 15206 11396 15258
rect 11396 15206 11442 15258
rect 11466 15206 11512 15258
rect 11512 15206 11522 15258
rect 11546 15206 11576 15258
rect 11576 15206 11602 15258
rect 11306 15204 11362 15206
rect 11386 15204 11442 15206
rect 11466 15204 11522 15206
rect 11546 15204 11602 15206
rect 7856 12538 7912 12540
rect 7936 12538 7992 12540
rect 8016 12538 8072 12540
rect 8096 12538 8152 12540
rect 7856 12486 7882 12538
rect 7882 12486 7912 12538
rect 7936 12486 7946 12538
rect 7946 12486 7992 12538
rect 8016 12486 8062 12538
rect 8062 12486 8072 12538
rect 8096 12486 8126 12538
rect 8126 12486 8152 12538
rect 7856 12484 7912 12486
rect 7936 12484 7992 12486
rect 8016 12484 8072 12486
rect 8096 12484 8152 12486
rect 7856 11450 7912 11452
rect 7936 11450 7992 11452
rect 8016 11450 8072 11452
rect 8096 11450 8152 11452
rect 7856 11398 7882 11450
rect 7882 11398 7912 11450
rect 7936 11398 7946 11450
rect 7946 11398 7992 11450
rect 8016 11398 8062 11450
rect 8062 11398 8072 11450
rect 8096 11398 8126 11450
rect 8126 11398 8152 11450
rect 7856 11396 7912 11398
rect 7936 11396 7992 11398
rect 8016 11396 8072 11398
rect 8096 11396 8152 11398
rect 7856 10362 7912 10364
rect 7936 10362 7992 10364
rect 8016 10362 8072 10364
rect 8096 10362 8152 10364
rect 7856 10310 7882 10362
rect 7882 10310 7912 10362
rect 7936 10310 7946 10362
rect 7946 10310 7992 10362
rect 8016 10310 8062 10362
rect 8062 10310 8072 10362
rect 8096 10310 8126 10362
rect 8126 10310 8152 10362
rect 7856 10308 7912 10310
rect 7936 10308 7992 10310
rect 8016 10308 8072 10310
rect 8096 10308 8152 10310
rect 7856 9274 7912 9276
rect 7936 9274 7992 9276
rect 8016 9274 8072 9276
rect 8096 9274 8152 9276
rect 7856 9222 7882 9274
rect 7882 9222 7912 9274
rect 7936 9222 7946 9274
rect 7946 9222 7992 9274
rect 8016 9222 8062 9274
rect 8062 9222 8072 9274
rect 8096 9222 8126 9274
rect 8126 9222 8152 9274
rect 7856 9220 7912 9222
rect 7936 9220 7992 9222
rect 8016 9220 8072 9222
rect 8096 9220 8152 9222
rect 7856 8186 7912 8188
rect 7936 8186 7992 8188
rect 8016 8186 8072 8188
rect 8096 8186 8152 8188
rect 7856 8134 7882 8186
rect 7882 8134 7912 8186
rect 7936 8134 7946 8186
rect 7946 8134 7992 8186
rect 8016 8134 8062 8186
rect 8062 8134 8072 8186
rect 8096 8134 8126 8186
rect 8126 8134 8152 8186
rect 7856 8132 7912 8134
rect 7936 8132 7992 8134
rect 8016 8132 8072 8134
rect 8096 8132 8152 8134
rect 7856 7098 7912 7100
rect 7936 7098 7992 7100
rect 8016 7098 8072 7100
rect 8096 7098 8152 7100
rect 7856 7046 7882 7098
rect 7882 7046 7912 7098
rect 7936 7046 7946 7098
rect 7946 7046 7992 7098
rect 8016 7046 8062 7098
rect 8062 7046 8072 7098
rect 8096 7046 8126 7098
rect 8126 7046 8152 7098
rect 7856 7044 7912 7046
rect 7936 7044 7992 7046
rect 8016 7044 8072 7046
rect 8096 7044 8152 7046
rect 7856 6010 7912 6012
rect 7936 6010 7992 6012
rect 8016 6010 8072 6012
rect 8096 6010 8152 6012
rect 7856 5958 7882 6010
rect 7882 5958 7912 6010
rect 7936 5958 7946 6010
rect 7946 5958 7992 6010
rect 8016 5958 8062 6010
rect 8062 5958 8072 6010
rect 8096 5958 8126 6010
rect 8126 5958 8152 6010
rect 7856 5956 7912 5958
rect 7936 5956 7992 5958
rect 8016 5956 8072 5958
rect 8096 5956 8152 5958
rect 11306 14170 11362 14172
rect 11386 14170 11442 14172
rect 11466 14170 11522 14172
rect 11546 14170 11602 14172
rect 11306 14118 11332 14170
rect 11332 14118 11362 14170
rect 11386 14118 11396 14170
rect 11396 14118 11442 14170
rect 11466 14118 11512 14170
rect 11512 14118 11522 14170
rect 11546 14118 11576 14170
rect 11576 14118 11602 14170
rect 11306 14116 11362 14118
rect 11386 14116 11442 14118
rect 11466 14116 11522 14118
rect 11546 14116 11602 14118
rect 11306 13082 11362 13084
rect 11386 13082 11442 13084
rect 11466 13082 11522 13084
rect 11546 13082 11602 13084
rect 11306 13030 11332 13082
rect 11332 13030 11362 13082
rect 11386 13030 11396 13082
rect 11396 13030 11442 13082
rect 11466 13030 11512 13082
rect 11512 13030 11522 13082
rect 11546 13030 11576 13082
rect 11576 13030 11602 13082
rect 11306 13028 11362 13030
rect 11386 13028 11442 13030
rect 11466 13028 11522 13030
rect 11546 13028 11602 13030
rect 7856 4922 7912 4924
rect 7936 4922 7992 4924
rect 8016 4922 8072 4924
rect 8096 4922 8152 4924
rect 7856 4870 7882 4922
rect 7882 4870 7912 4922
rect 7936 4870 7946 4922
rect 7946 4870 7992 4922
rect 8016 4870 8062 4922
rect 8062 4870 8072 4922
rect 8096 4870 8126 4922
rect 8126 4870 8152 4922
rect 7856 4868 7912 4870
rect 7936 4868 7992 4870
rect 8016 4868 8072 4870
rect 8096 4868 8152 4870
rect 7856 3834 7912 3836
rect 7936 3834 7992 3836
rect 8016 3834 8072 3836
rect 8096 3834 8152 3836
rect 7856 3782 7882 3834
rect 7882 3782 7912 3834
rect 7936 3782 7946 3834
rect 7946 3782 7992 3834
rect 8016 3782 8062 3834
rect 8062 3782 8072 3834
rect 8096 3782 8126 3834
rect 8126 3782 8152 3834
rect 7856 3780 7912 3782
rect 7936 3780 7992 3782
rect 8016 3780 8072 3782
rect 8096 3780 8152 3782
rect 7856 2746 7912 2748
rect 7936 2746 7992 2748
rect 8016 2746 8072 2748
rect 8096 2746 8152 2748
rect 7856 2694 7882 2746
rect 7882 2694 7912 2746
rect 7936 2694 7946 2746
rect 7946 2694 7992 2746
rect 8016 2694 8062 2746
rect 8062 2694 8072 2746
rect 8096 2694 8126 2746
rect 8126 2694 8152 2746
rect 7856 2692 7912 2694
rect 7936 2692 7992 2694
rect 8016 2692 8072 2694
rect 8096 2692 8152 2694
rect 11306 11994 11362 11996
rect 11386 11994 11442 11996
rect 11466 11994 11522 11996
rect 11546 11994 11602 11996
rect 11306 11942 11332 11994
rect 11332 11942 11362 11994
rect 11386 11942 11396 11994
rect 11396 11942 11442 11994
rect 11466 11942 11512 11994
rect 11512 11942 11522 11994
rect 11546 11942 11576 11994
rect 11576 11942 11602 11994
rect 11306 11940 11362 11942
rect 11386 11940 11442 11942
rect 11466 11940 11522 11942
rect 11546 11940 11602 11942
rect 11306 10906 11362 10908
rect 11386 10906 11442 10908
rect 11466 10906 11522 10908
rect 11546 10906 11602 10908
rect 11306 10854 11332 10906
rect 11332 10854 11362 10906
rect 11386 10854 11396 10906
rect 11396 10854 11442 10906
rect 11466 10854 11512 10906
rect 11512 10854 11522 10906
rect 11546 10854 11576 10906
rect 11576 10854 11602 10906
rect 11306 10852 11362 10854
rect 11386 10852 11442 10854
rect 11466 10852 11522 10854
rect 11546 10852 11602 10854
rect 11306 9818 11362 9820
rect 11386 9818 11442 9820
rect 11466 9818 11522 9820
rect 11546 9818 11602 9820
rect 11306 9766 11332 9818
rect 11332 9766 11362 9818
rect 11386 9766 11396 9818
rect 11396 9766 11442 9818
rect 11466 9766 11512 9818
rect 11512 9766 11522 9818
rect 11546 9766 11576 9818
rect 11576 9766 11602 9818
rect 11306 9764 11362 9766
rect 11386 9764 11442 9766
rect 11466 9764 11522 9766
rect 11546 9764 11602 9766
rect 11306 8730 11362 8732
rect 11386 8730 11442 8732
rect 11466 8730 11522 8732
rect 11546 8730 11602 8732
rect 11306 8678 11332 8730
rect 11332 8678 11362 8730
rect 11386 8678 11396 8730
rect 11396 8678 11442 8730
rect 11466 8678 11512 8730
rect 11512 8678 11522 8730
rect 11546 8678 11576 8730
rect 11576 8678 11602 8730
rect 11306 8676 11362 8678
rect 11386 8676 11442 8678
rect 11466 8676 11522 8678
rect 11546 8676 11602 8678
rect 11306 7642 11362 7644
rect 11386 7642 11442 7644
rect 11466 7642 11522 7644
rect 11546 7642 11602 7644
rect 11306 7590 11332 7642
rect 11332 7590 11362 7642
rect 11386 7590 11396 7642
rect 11396 7590 11442 7642
rect 11466 7590 11512 7642
rect 11512 7590 11522 7642
rect 11546 7590 11576 7642
rect 11576 7590 11602 7642
rect 11306 7588 11362 7590
rect 11386 7588 11442 7590
rect 11466 7588 11522 7590
rect 11546 7588 11602 7590
rect 14756 21242 14812 21244
rect 14836 21242 14892 21244
rect 14916 21242 14972 21244
rect 14996 21242 15052 21244
rect 14756 21190 14782 21242
rect 14782 21190 14812 21242
rect 14836 21190 14846 21242
rect 14846 21190 14892 21242
rect 14916 21190 14962 21242
rect 14962 21190 14972 21242
rect 14996 21190 15026 21242
rect 15026 21190 15052 21242
rect 14756 21188 14812 21190
rect 14836 21188 14892 21190
rect 14916 21188 14972 21190
rect 14996 21188 15052 21190
rect 14756 20154 14812 20156
rect 14836 20154 14892 20156
rect 14916 20154 14972 20156
rect 14996 20154 15052 20156
rect 14756 20102 14782 20154
rect 14782 20102 14812 20154
rect 14836 20102 14846 20154
rect 14846 20102 14892 20154
rect 14916 20102 14962 20154
rect 14962 20102 14972 20154
rect 14996 20102 15026 20154
rect 15026 20102 15052 20154
rect 14756 20100 14812 20102
rect 14836 20100 14892 20102
rect 14916 20100 14972 20102
rect 14996 20100 15052 20102
rect 14554 19216 14610 19272
rect 14756 19066 14812 19068
rect 14836 19066 14892 19068
rect 14916 19066 14972 19068
rect 14996 19066 15052 19068
rect 14756 19014 14782 19066
rect 14782 19014 14812 19066
rect 14836 19014 14846 19066
rect 14846 19014 14892 19066
rect 14916 19014 14962 19066
rect 14962 19014 14972 19066
rect 14996 19014 15026 19066
rect 15026 19014 15052 19066
rect 14756 19012 14812 19014
rect 14836 19012 14892 19014
rect 14916 19012 14972 19014
rect 14996 19012 15052 19014
rect 15198 19216 15254 19272
rect 14756 17978 14812 17980
rect 14836 17978 14892 17980
rect 14916 17978 14972 17980
rect 14996 17978 15052 17980
rect 14756 17926 14782 17978
rect 14782 17926 14812 17978
rect 14836 17926 14846 17978
rect 14846 17926 14892 17978
rect 14916 17926 14962 17978
rect 14962 17926 14972 17978
rect 14996 17926 15026 17978
rect 15026 17926 15052 17978
rect 14756 17924 14812 17926
rect 14836 17924 14892 17926
rect 14916 17924 14972 17926
rect 14996 17924 15052 17926
rect 14756 16890 14812 16892
rect 14836 16890 14892 16892
rect 14916 16890 14972 16892
rect 14996 16890 15052 16892
rect 14756 16838 14782 16890
rect 14782 16838 14812 16890
rect 14836 16838 14846 16890
rect 14846 16838 14892 16890
rect 14916 16838 14962 16890
rect 14962 16838 14972 16890
rect 14996 16838 15026 16890
rect 15026 16838 15052 16890
rect 14756 16836 14812 16838
rect 14836 16836 14892 16838
rect 14916 16836 14972 16838
rect 14996 16836 15052 16838
rect 15658 19252 15660 19272
rect 15660 19252 15712 19272
rect 15712 19252 15714 19272
rect 15658 19216 15714 19252
rect 15750 19080 15806 19136
rect 14756 15802 14812 15804
rect 14836 15802 14892 15804
rect 14916 15802 14972 15804
rect 14996 15802 15052 15804
rect 14756 15750 14782 15802
rect 14782 15750 14812 15802
rect 14836 15750 14846 15802
rect 14846 15750 14892 15802
rect 14916 15750 14962 15802
rect 14962 15750 14972 15802
rect 14996 15750 15026 15802
rect 15026 15750 15052 15802
rect 14756 15748 14812 15750
rect 14836 15748 14892 15750
rect 14916 15748 14972 15750
rect 14996 15748 15052 15750
rect 14646 15000 14702 15056
rect 14756 14714 14812 14716
rect 14836 14714 14892 14716
rect 14916 14714 14972 14716
rect 14996 14714 15052 14716
rect 14756 14662 14782 14714
rect 14782 14662 14812 14714
rect 14836 14662 14846 14714
rect 14846 14662 14892 14714
rect 14916 14662 14962 14714
rect 14962 14662 14972 14714
rect 14996 14662 15026 14714
rect 15026 14662 15052 14714
rect 14756 14660 14812 14662
rect 14836 14660 14892 14662
rect 14916 14660 14972 14662
rect 14996 14660 15052 14662
rect 14756 13626 14812 13628
rect 14836 13626 14892 13628
rect 14916 13626 14972 13628
rect 14996 13626 15052 13628
rect 14756 13574 14782 13626
rect 14782 13574 14812 13626
rect 14836 13574 14846 13626
rect 14846 13574 14892 13626
rect 14916 13574 14962 13626
rect 14962 13574 14972 13626
rect 14996 13574 15026 13626
rect 15026 13574 15052 13626
rect 14756 13572 14812 13574
rect 14836 13572 14892 13574
rect 14916 13572 14972 13574
rect 14996 13572 15052 13574
rect 15290 15000 15346 15056
rect 15290 14476 15346 14512
rect 15290 14456 15292 14476
rect 15292 14456 15344 14476
rect 15344 14456 15346 14476
rect 14756 12538 14812 12540
rect 14836 12538 14892 12540
rect 14916 12538 14972 12540
rect 14996 12538 15052 12540
rect 14756 12486 14782 12538
rect 14782 12486 14812 12538
rect 14836 12486 14846 12538
rect 14846 12486 14892 12538
rect 14916 12486 14962 12538
rect 14962 12486 14972 12538
rect 14996 12486 15026 12538
rect 15026 12486 15052 12538
rect 14756 12484 14812 12486
rect 14836 12484 14892 12486
rect 14916 12484 14972 12486
rect 14996 12484 15052 12486
rect 17682 19372 17738 19408
rect 17682 19352 17684 19372
rect 17684 19352 17736 19372
rect 17736 19352 17738 19372
rect 11306 6554 11362 6556
rect 11386 6554 11442 6556
rect 11466 6554 11522 6556
rect 11546 6554 11602 6556
rect 11306 6502 11332 6554
rect 11332 6502 11362 6554
rect 11386 6502 11396 6554
rect 11396 6502 11442 6554
rect 11466 6502 11512 6554
rect 11512 6502 11522 6554
rect 11546 6502 11576 6554
rect 11576 6502 11602 6554
rect 11306 6500 11362 6502
rect 11386 6500 11442 6502
rect 11466 6500 11522 6502
rect 11546 6500 11602 6502
rect 11306 5466 11362 5468
rect 11386 5466 11442 5468
rect 11466 5466 11522 5468
rect 11546 5466 11602 5468
rect 11306 5414 11332 5466
rect 11332 5414 11362 5466
rect 11386 5414 11396 5466
rect 11396 5414 11442 5466
rect 11466 5414 11512 5466
rect 11512 5414 11522 5466
rect 11546 5414 11576 5466
rect 11576 5414 11602 5466
rect 11306 5412 11362 5414
rect 11386 5412 11442 5414
rect 11466 5412 11522 5414
rect 11546 5412 11602 5414
rect 11306 4378 11362 4380
rect 11386 4378 11442 4380
rect 11466 4378 11522 4380
rect 11546 4378 11602 4380
rect 11306 4326 11332 4378
rect 11332 4326 11362 4378
rect 11386 4326 11396 4378
rect 11396 4326 11442 4378
rect 11466 4326 11512 4378
rect 11512 4326 11522 4378
rect 11546 4326 11576 4378
rect 11576 4326 11602 4378
rect 11306 4324 11362 4326
rect 11386 4324 11442 4326
rect 11466 4324 11522 4326
rect 11546 4324 11602 4326
rect 11306 3290 11362 3292
rect 11386 3290 11442 3292
rect 11466 3290 11522 3292
rect 11546 3290 11602 3292
rect 11306 3238 11332 3290
rect 11332 3238 11362 3290
rect 11386 3238 11396 3290
rect 11396 3238 11442 3290
rect 11466 3238 11512 3290
rect 11512 3238 11522 3290
rect 11546 3238 11576 3290
rect 11576 3238 11602 3290
rect 11306 3236 11362 3238
rect 11386 3236 11442 3238
rect 11466 3236 11522 3238
rect 11546 3236 11602 3238
rect 14756 11450 14812 11452
rect 14836 11450 14892 11452
rect 14916 11450 14972 11452
rect 14996 11450 15052 11452
rect 14756 11398 14782 11450
rect 14782 11398 14812 11450
rect 14836 11398 14846 11450
rect 14846 11398 14892 11450
rect 14916 11398 14962 11450
rect 14962 11398 14972 11450
rect 14996 11398 15026 11450
rect 15026 11398 15052 11450
rect 14756 11396 14812 11398
rect 14836 11396 14892 11398
rect 14916 11396 14972 11398
rect 14996 11396 15052 11398
rect 14756 10362 14812 10364
rect 14836 10362 14892 10364
rect 14916 10362 14972 10364
rect 14996 10362 15052 10364
rect 14756 10310 14782 10362
rect 14782 10310 14812 10362
rect 14836 10310 14846 10362
rect 14846 10310 14892 10362
rect 14916 10310 14962 10362
rect 14962 10310 14972 10362
rect 14996 10310 15026 10362
rect 15026 10310 15052 10362
rect 14756 10308 14812 10310
rect 14836 10308 14892 10310
rect 14916 10308 14972 10310
rect 14996 10308 15052 10310
rect 14756 9274 14812 9276
rect 14836 9274 14892 9276
rect 14916 9274 14972 9276
rect 14996 9274 15052 9276
rect 14756 9222 14782 9274
rect 14782 9222 14812 9274
rect 14836 9222 14846 9274
rect 14846 9222 14892 9274
rect 14916 9222 14962 9274
rect 14962 9222 14972 9274
rect 14996 9222 15026 9274
rect 15026 9222 15052 9274
rect 14756 9220 14812 9222
rect 14836 9220 14892 9222
rect 14916 9220 14972 9222
rect 14996 9220 15052 9222
rect 14756 8186 14812 8188
rect 14836 8186 14892 8188
rect 14916 8186 14972 8188
rect 14996 8186 15052 8188
rect 14756 8134 14782 8186
rect 14782 8134 14812 8186
rect 14836 8134 14846 8186
rect 14846 8134 14892 8186
rect 14916 8134 14962 8186
rect 14962 8134 14972 8186
rect 14996 8134 15026 8186
rect 15026 8134 15052 8186
rect 14756 8132 14812 8134
rect 14836 8132 14892 8134
rect 14916 8132 14972 8134
rect 14996 8132 15052 8134
rect 18206 21786 18262 21788
rect 18286 21786 18342 21788
rect 18366 21786 18422 21788
rect 18446 21786 18502 21788
rect 18206 21734 18232 21786
rect 18232 21734 18262 21786
rect 18286 21734 18296 21786
rect 18296 21734 18342 21786
rect 18366 21734 18412 21786
rect 18412 21734 18422 21786
rect 18446 21734 18476 21786
rect 18476 21734 18502 21786
rect 18206 21732 18262 21734
rect 18286 21732 18342 21734
rect 18366 21732 18422 21734
rect 18446 21732 18502 21734
rect 18206 20698 18262 20700
rect 18286 20698 18342 20700
rect 18366 20698 18422 20700
rect 18446 20698 18502 20700
rect 18206 20646 18232 20698
rect 18232 20646 18262 20698
rect 18286 20646 18296 20698
rect 18296 20646 18342 20698
rect 18366 20646 18412 20698
rect 18412 20646 18422 20698
rect 18446 20646 18476 20698
rect 18476 20646 18502 20698
rect 18206 20644 18262 20646
rect 18286 20644 18342 20646
rect 18366 20644 18422 20646
rect 18446 20644 18502 20646
rect 18206 19610 18262 19612
rect 18286 19610 18342 19612
rect 18366 19610 18422 19612
rect 18446 19610 18502 19612
rect 18206 19558 18232 19610
rect 18232 19558 18262 19610
rect 18286 19558 18296 19610
rect 18296 19558 18342 19610
rect 18366 19558 18412 19610
rect 18412 19558 18422 19610
rect 18446 19558 18476 19610
rect 18476 19558 18502 19610
rect 18206 19556 18262 19558
rect 18286 19556 18342 19558
rect 18366 19556 18422 19558
rect 18446 19556 18502 19558
rect 18602 19116 18604 19136
rect 18604 19116 18656 19136
rect 18656 19116 18658 19136
rect 18602 19080 18658 19116
rect 18206 18522 18262 18524
rect 18286 18522 18342 18524
rect 18366 18522 18422 18524
rect 18446 18522 18502 18524
rect 18206 18470 18232 18522
rect 18232 18470 18262 18522
rect 18286 18470 18296 18522
rect 18296 18470 18342 18522
rect 18366 18470 18412 18522
rect 18412 18470 18422 18522
rect 18446 18470 18476 18522
rect 18476 18470 18502 18522
rect 18206 18468 18262 18470
rect 18286 18468 18342 18470
rect 18366 18468 18422 18470
rect 18446 18468 18502 18470
rect 18206 17434 18262 17436
rect 18286 17434 18342 17436
rect 18366 17434 18422 17436
rect 18446 17434 18502 17436
rect 18206 17382 18232 17434
rect 18232 17382 18262 17434
rect 18286 17382 18296 17434
rect 18296 17382 18342 17434
rect 18366 17382 18412 17434
rect 18412 17382 18422 17434
rect 18446 17382 18476 17434
rect 18476 17382 18502 17434
rect 18206 17380 18262 17382
rect 18286 17380 18342 17382
rect 18366 17380 18422 17382
rect 18446 17380 18502 17382
rect 18206 16346 18262 16348
rect 18286 16346 18342 16348
rect 18366 16346 18422 16348
rect 18446 16346 18502 16348
rect 18206 16294 18232 16346
rect 18232 16294 18262 16346
rect 18286 16294 18296 16346
rect 18296 16294 18342 16346
rect 18366 16294 18412 16346
rect 18412 16294 18422 16346
rect 18446 16294 18476 16346
rect 18476 16294 18502 16346
rect 18206 16292 18262 16294
rect 18286 16292 18342 16294
rect 18366 16292 18422 16294
rect 18446 16292 18502 16294
rect 18206 15258 18262 15260
rect 18286 15258 18342 15260
rect 18366 15258 18422 15260
rect 18446 15258 18502 15260
rect 18206 15206 18232 15258
rect 18232 15206 18262 15258
rect 18286 15206 18296 15258
rect 18296 15206 18342 15258
rect 18366 15206 18412 15258
rect 18412 15206 18422 15258
rect 18446 15206 18476 15258
rect 18476 15206 18502 15258
rect 18206 15204 18262 15206
rect 18286 15204 18342 15206
rect 18366 15204 18422 15206
rect 18446 15204 18502 15206
rect 20626 20440 20682 20496
rect 20626 17720 20682 17776
rect 19246 14456 19302 14512
rect 18206 14170 18262 14172
rect 18286 14170 18342 14172
rect 18366 14170 18422 14172
rect 18446 14170 18502 14172
rect 18206 14118 18232 14170
rect 18232 14118 18262 14170
rect 18286 14118 18296 14170
rect 18296 14118 18342 14170
rect 18366 14118 18412 14170
rect 18412 14118 18422 14170
rect 18446 14118 18476 14170
rect 18476 14118 18502 14170
rect 18206 14116 18262 14118
rect 18286 14116 18342 14118
rect 18366 14116 18422 14118
rect 18446 14116 18502 14118
rect 18206 13082 18262 13084
rect 18286 13082 18342 13084
rect 18366 13082 18422 13084
rect 18446 13082 18502 13084
rect 18206 13030 18232 13082
rect 18232 13030 18262 13082
rect 18286 13030 18296 13082
rect 18296 13030 18342 13082
rect 18366 13030 18412 13082
rect 18412 13030 18422 13082
rect 18446 13030 18476 13082
rect 18476 13030 18502 13082
rect 18206 13028 18262 13030
rect 18286 13028 18342 13030
rect 18366 13028 18422 13030
rect 18446 13028 18502 13030
rect 21086 15680 21142 15736
rect 21086 12960 21142 13016
rect 18206 11994 18262 11996
rect 18286 11994 18342 11996
rect 18366 11994 18422 11996
rect 18446 11994 18502 11996
rect 18206 11942 18232 11994
rect 18232 11942 18262 11994
rect 18286 11942 18296 11994
rect 18296 11942 18342 11994
rect 18366 11942 18412 11994
rect 18412 11942 18422 11994
rect 18446 11942 18476 11994
rect 18476 11942 18502 11994
rect 18206 11940 18262 11942
rect 18286 11940 18342 11942
rect 18366 11940 18422 11942
rect 18446 11940 18502 11942
rect 18206 10906 18262 10908
rect 18286 10906 18342 10908
rect 18366 10906 18422 10908
rect 18446 10906 18502 10908
rect 18206 10854 18232 10906
rect 18232 10854 18262 10906
rect 18286 10854 18296 10906
rect 18296 10854 18342 10906
rect 18366 10854 18412 10906
rect 18412 10854 18422 10906
rect 18446 10854 18476 10906
rect 18476 10854 18502 10906
rect 18206 10852 18262 10854
rect 18286 10852 18342 10854
rect 18366 10852 18422 10854
rect 18446 10852 18502 10854
rect 21086 10240 21142 10296
rect 18206 9818 18262 9820
rect 18286 9818 18342 9820
rect 18366 9818 18422 9820
rect 18446 9818 18502 9820
rect 18206 9766 18232 9818
rect 18232 9766 18262 9818
rect 18286 9766 18296 9818
rect 18296 9766 18342 9818
rect 18366 9766 18412 9818
rect 18412 9766 18422 9818
rect 18446 9766 18476 9818
rect 18476 9766 18502 9818
rect 18206 9764 18262 9766
rect 18286 9764 18342 9766
rect 18366 9764 18422 9766
rect 18446 9764 18502 9766
rect 18206 8730 18262 8732
rect 18286 8730 18342 8732
rect 18366 8730 18422 8732
rect 18446 8730 18502 8732
rect 18206 8678 18232 8730
rect 18232 8678 18262 8730
rect 18286 8678 18296 8730
rect 18296 8678 18342 8730
rect 18366 8678 18412 8730
rect 18412 8678 18422 8730
rect 18446 8678 18476 8730
rect 18476 8678 18502 8730
rect 18206 8676 18262 8678
rect 18286 8676 18342 8678
rect 18366 8676 18422 8678
rect 18446 8676 18502 8678
rect 21086 8200 21142 8256
rect 14756 7098 14812 7100
rect 14836 7098 14892 7100
rect 14916 7098 14972 7100
rect 14996 7098 15052 7100
rect 14756 7046 14782 7098
rect 14782 7046 14812 7098
rect 14836 7046 14846 7098
rect 14846 7046 14892 7098
rect 14916 7046 14962 7098
rect 14962 7046 14972 7098
rect 14996 7046 15026 7098
rect 15026 7046 15052 7098
rect 14756 7044 14812 7046
rect 14836 7044 14892 7046
rect 14916 7044 14972 7046
rect 14996 7044 15052 7046
rect 14756 6010 14812 6012
rect 14836 6010 14892 6012
rect 14916 6010 14972 6012
rect 14996 6010 15052 6012
rect 14756 5958 14782 6010
rect 14782 5958 14812 6010
rect 14836 5958 14846 6010
rect 14846 5958 14892 6010
rect 14916 5958 14962 6010
rect 14962 5958 14972 6010
rect 14996 5958 15026 6010
rect 15026 5958 15052 6010
rect 14756 5956 14812 5958
rect 14836 5956 14892 5958
rect 14916 5956 14972 5958
rect 14996 5956 15052 5958
rect 14756 4922 14812 4924
rect 14836 4922 14892 4924
rect 14916 4922 14972 4924
rect 14996 4922 15052 4924
rect 14756 4870 14782 4922
rect 14782 4870 14812 4922
rect 14836 4870 14846 4922
rect 14846 4870 14892 4922
rect 14916 4870 14962 4922
rect 14962 4870 14972 4922
rect 14996 4870 15026 4922
rect 15026 4870 15052 4922
rect 14756 4868 14812 4870
rect 14836 4868 14892 4870
rect 14916 4868 14972 4870
rect 14996 4868 15052 4870
rect 4406 2202 4462 2204
rect 4486 2202 4542 2204
rect 4566 2202 4622 2204
rect 4646 2202 4702 2204
rect 4406 2150 4432 2202
rect 4432 2150 4462 2202
rect 4486 2150 4496 2202
rect 4496 2150 4542 2202
rect 4566 2150 4612 2202
rect 4612 2150 4622 2202
rect 4646 2150 4676 2202
rect 4676 2150 4702 2202
rect 4406 2148 4462 2150
rect 4486 2148 4542 2150
rect 4566 2148 4622 2150
rect 4646 2148 4702 2150
rect 11306 2202 11362 2204
rect 11386 2202 11442 2204
rect 11466 2202 11522 2204
rect 11546 2202 11602 2204
rect 11306 2150 11332 2202
rect 11332 2150 11362 2202
rect 11386 2150 11396 2202
rect 11396 2150 11442 2202
rect 11466 2150 11512 2202
rect 11512 2150 11522 2202
rect 11546 2150 11576 2202
rect 11576 2150 11602 2202
rect 11306 2148 11362 2150
rect 11386 2148 11442 2150
rect 11466 2148 11522 2150
rect 11546 2148 11602 2150
rect 14756 3834 14812 3836
rect 14836 3834 14892 3836
rect 14916 3834 14972 3836
rect 14996 3834 15052 3836
rect 14756 3782 14782 3834
rect 14782 3782 14812 3834
rect 14836 3782 14846 3834
rect 14846 3782 14892 3834
rect 14916 3782 14962 3834
rect 14962 3782 14972 3834
rect 14996 3782 15026 3834
rect 15026 3782 15052 3834
rect 14756 3780 14812 3782
rect 14836 3780 14892 3782
rect 14916 3780 14972 3782
rect 14996 3780 15052 3782
rect 14756 2746 14812 2748
rect 14836 2746 14892 2748
rect 14916 2746 14972 2748
rect 14996 2746 15052 2748
rect 14756 2694 14782 2746
rect 14782 2694 14812 2746
rect 14836 2694 14846 2746
rect 14846 2694 14892 2746
rect 14916 2694 14962 2746
rect 14962 2694 14972 2746
rect 14996 2694 15026 2746
rect 15026 2694 15052 2746
rect 14756 2692 14812 2694
rect 14836 2692 14892 2694
rect 14916 2692 14972 2694
rect 14996 2692 15052 2694
rect 18206 7642 18262 7644
rect 18286 7642 18342 7644
rect 18366 7642 18422 7644
rect 18446 7642 18502 7644
rect 18206 7590 18232 7642
rect 18232 7590 18262 7642
rect 18286 7590 18296 7642
rect 18296 7590 18342 7642
rect 18366 7590 18412 7642
rect 18412 7590 18422 7642
rect 18446 7590 18476 7642
rect 18476 7590 18502 7642
rect 18206 7588 18262 7590
rect 18286 7588 18342 7590
rect 18366 7588 18422 7590
rect 18446 7588 18502 7590
rect 18206 6554 18262 6556
rect 18286 6554 18342 6556
rect 18366 6554 18422 6556
rect 18446 6554 18502 6556
rect 18206 6502 18232 6554
rect 18232 6502 18262 6554
rect 18286 6502 18296 6554
rect 18296 6502 18342 6554
rect 18366 6502 18412 6554
rect 18412 6502 18422 6554
rect 18446 6502 18476 6554
rect 18476 6502 18502 6554
rect 18206 6500 18262 6502
rect 18286 6500 18342 6502
rect 18366 6500 18422 6502
rect 18446 6500 18502 6502
rect 18206 5466 18262 5468
rect 18286 5466 18342 5468
rect 18366 5466 18422 5468
rect 18446 5466 18502 5468
rect 18206 5414 18232 5466
rect 18232 5414 18262 5466
rect 18286 5414 18296 5466
rect 18296 5414 18342 5466
rect 18366 5414 18412 5466
rect 18412 5414 18422 5466
rect 18446 5414 18476 5466
rect 18476 5414 18502 5466
rect 18206 5412 18262 5414
rect 18286 5412 18342 5414
rect 18366 5412 18422 5414
rect 18446 5412 18502 5414
rect 18206 4378 18262 4380
rect 18286 4378 18342 4380
rect 18366 4378 18422 4380
rect 18446 4378 18502 4380
rect 18206 4326 18232 4378
rect 18232 4326 18262 4378
rect 18286 4326 18296 4378
rect 18296 4326 18342 4378
rect 18366 4326 18412 4378
rect 18412 4326 18422 4378
rect 18446 4326 18476 4378
rect 18476 4326 18502 4378
rect 18206 4324 18262 4326
rect 18286 4324 18342 4326
rect 18366 4324 18422 4326
rect 18446 4324 18502 4326
rect 18206 3290 18262 3292
rect 18286 3290 18342 3292
rect 18366 3290 18422 3292
rect 18446 3290 18502 3292
rect 18206 3238 18232 3290
rect 18232 3238 18262 3290
rect 18286 3238 18296 3290
rect 18296 3238 18342 3290
rect 18366 3238 18412 3290
rect 18412 3238 18422 3290
rect 18446 3238 18476 3290
rect 18476 3238 18502 3290
rect 18206 3236 18262 3238
rect 18286 3236 18342 3238
rect 18366 3236 18422 3238
rect 18446 3236 18502 3238
rect 20074 2760 20130 2816
rect 21086 5480 21142 5536
rect 18206 2202 18262 2204
rect 18286 2202 18342 2204
rect 18366 2202 18422 2204
rect 18446 2202 18502 2204
rect 18206 2150 18232 2202
rect 18232 2150 18262 2202
rect 18286 2150 18296 2202
rect 18296 2150 18342 2202
rect 18366 2150 18412 2202
rect 18412 2150 18422 2202
rect 18446 2150 18476 2202
rect 18476 2150 18502 2202
rect 18206 2148 18262 2150
rect 18286 2148 18342 2150
rect 18366 2148 18422 2150
rect 18446 2148 18502 2150
<< metal3 >>
rect 0 23218 800 23248
rect 1485 23218 1551 23221
rect 0 23216 1551 23218
rect 0 23160 1490 23216
rect 1546 23160 1551 23216
rect 0 23158 1551 23160
rect 0 23128 800 23158
rect 1485 23155 1551 23158
rect 21081 23218 21147 23221
rect 22179 23218 22979 23248
rect 21081 23216 22979 23218
rect 21081 23160 21086 23216
rect 21142 23160 22979 23216
rect 21081 23158 22979 23160
rect 21081 23155 21147 23158
rect 22179 23128 22979 23158
rect 4394 22880 4714 22881
rect 4394 22816 4402 22880
rect 4466 22816 4482 22880
rect 4546 22816 4562 22880
rect 4626 22816 4642 22880
rect 4706 22816 4714 22880
rect 4394 22815 4714 22816
rect 11294 22880 11614 22881
rect 11294 22816 11302 22880
rect 11366 22816 11382 22880
rect 11446 22816 11462 22880
rect 11526 22816 11542 22880
rect 11606 22816 11614 22880
rect 11294 22815 11614 22816
rect 18194 22880 18514 22881
rect 18194 22816 18202 22880
rect 18266 22816 18282 22880
rect 18346 22816 18362 22880
rect 18426 22816 18442 22880
rect 18506 22816 18514 22880
rect 18194 22815 18514 22816
rect 7844 22336 8164 22337
rect 7844 22272 7852 22336
rect 7916 22272 7932 22336
rect 7996 22272 8012 22336
rect 8076 22272 8092 22336
rect 8156 22272 8164 22336
rect 7844 22271 8164 22272
rect 14744 22336 15064 22337
rect 14744 22272 14752 22336
rect 14816 22272 14832 22336
rect 14896 22272 14912 22336
rect 14976 22272 14992 22336
rect 15056 22272 15064 22336
rect 14744 22271 15064 22272
rect 4394 21792 4714 21793
rect 4394 21728 4402 21792
rect 4466 21728 4482 21792
rect 4546 21728 4562 21792
rect 4626 21728 4642 21792
rect 4706 21728 4714 21792
rect 4394 21727 4714 21728
rect 11294 21792 11614 21793
rect 11294 21728 11302 21792
rect 11366 21728 11382 21792
rect 11446 21728 11462 21792
rect 11526 21728 11542 21792
rect 11606 21728 11614 21792
rect 11294 21727 11614 21728
rect 18194 21792 18514 21793
rect 18194 21728 18202 21792
rect 18266 21728 18282 21792
rect 18346 21728 18362 21792
rect 18426 21728 18442 21792
rect 18506 21728 18514 21792
rect 18194 21727 18514 21728
rect 7844 21248 8164 21249
rect 7844 21184 7852 21248
rect 7916 21184 7932 21248
rect 7996 21184 8012 21248
rect 8076 21184 8092 21248
rect 8156 21184 8164 21248
rect 7844 21183 8164 21184
rect 14744 21248 15064 21249
rect 14744 21184 14752 21248
rect 14816 21184 14832 21248
rect 14896 21184 14912 21248
rect 14976 21184 14992 21248
rect 15056 21184 15064 21248
rect 14744 21183 15064 21184
rect 4394 20704 4714 20705
rect 4394 20640 4402 20704
rect 4466 20640 4482 20704
rect 4546 20640 4562 20704
rect 4626 20640 4642 20704
rect 4706 20640 4714 20704
rect 4394 20639 4714 20640
rect 11294 20704 11614 20705
rect 11294 20640 11302 20704
rect 11366 20640 11382 20704
rect 11446 20640 11462 20704
rect 11526 20640 11542 20704
rect 11606 20640 11614 20704
rect 11294 20639 11614 20640
rect 18194 20704 18514 20705
rect 18194 20640 18202 20704
rect 18266 20640 18282 20704
rect 18346 20640 18362 20704
rect 18426 20640 18442 20704
rect 18506 20640 18514 20704
rect 18194 20639 18514 20640
rect 0 20498 800 20528
rect 1393 20498 1459 20501
rect 0 20496 1459 20498
rect 0 20440 1398 20496
rect 1454 20440 1459 20496
rect 0 20438 1459 20440
rect 0 20408 800 20438
rect 1393 20435 1459 20438
rect 20621 20498 20687 20501
rect 22179 20498 22979 20528
rect 20621 20496 22979 20498
rect 20621 20440 20626 20496
rect 20682 20440 22979 20496
rect 20621 20438 22979 20440
rect 20621 20435 20687 20438
rect 22179 20408 22979 20438
rect 7844 20160 8164 20161
rect 7844 20096 7852 20160
rect 7916 20096 7932 20160
rect 7996 20096 8012 20160
rect 8076 20096 8092 20160
rect 8156 20096 8164 20160
rect 7844 20095 8164 20096
rect 14744 20160 15064 20161
rect 14744 20096 14752 20160
rect 14816 20096 14832 20160
rect 14896 20096 14912 20160
rect 14976 20096 14992 20160
rect 15056 20096 15064 20160
rect 14744 20095 15064 20096
rect 4394 19616 4714 19617
rect 4394 19552 4402 19616
rect 4466 19552 4482 19616
rect 4546 19552 4562 19616
rect 4626 19552 4642 19616
rect 4706 19552 4714 19616
rect 4394 19551 4714 19552
rect 11294 19616 11614 19617
rect 11294 19552 11302 19616
rect 11366 19552 11382 19616
rect 11446 19552 11462 19616
rect 11526 19552 11542 19616
rect 11606 19552 11614 19616
rect 11294 19551 11614 19552
rect 18194 19616 18514 19617
rect 18194 19552 18202 19616
rect 18266 19552 18282 19616
rect 18346 19552 18362 19616
rect 18426 19552 18442 19616
rect 18506 19552 18514 19616
rect 18194 19551 18514 19552
rect 12617 19410 12683 19413
rect 17677 19410 17743 19413
rect 12617 19408 17743 19410
rect 12617 19352 12622 19408
rect 12678 19352 17682 19408
rect 17738 19352 17743 19408
rect 12617 19350 17743 19352
rect 12617 19347 12683 19350
rect 17677 19347 17743 19350
rect 14549 19274 14615 19277
rect 15193 19274 15259 19277
rect 15653 19274 15719 19277
rect 14549 19272 15719 19274
rect 14549 19216 14554 19272
rect 14610 19216 15198 19272
rect 15254 19216 15658 19272
rect 15714 19216 15719 19272
rect 14549 19214 15719 19216
rect 14549 19211 14615 19214
rect 15193 19211 15259 19214
rect 15653 19211 15719 19214
rect 15745 19138 15811 19141
rect 18597 19138 18663 19141
rect 15745 19136 18663 19138
rect 15745 19080 15750 19136
rect 15806 19080 18602 19136
rect 18658 19080 18663 19136
rect 15745 19078 18663 19080
rect 15745 19075 15811 19078
rect 18597 19075 18663 19078
rect 7844 19072 8164 19073
rect 7844 19008 7852 19072
rect 7916 19008 7932 19072
rect 7996 19008 8012 19072
rect 8076 19008 8092 19072
rect 8156 19008 8164 19072
rect 7844 19007 8164 19008
rect 14744 19072 15064 19073
rect 14744 19008 14752 19072
rect 14816 19008 14832 19072
rect 14896 19008 14912 19072
rect 14976 19008 14992 19072
rect 15056 19008 15064 19072
rect 14744 19007 15064 19008
rect 4394 18528 4714 18529
rect 4394 18464 4402 18528
rect 4466 18464 4482 18528
rect 4546 18464 4562 18528
rect 4626 18464 4642 18528
rect 4706 18464 4714 18528
rect 4394 18463 4714 18464
rect 11294 18528 11614 18529
rect 11294 18464 11302 18528
rect 11366 18464 11382 18528
rect 11446 18464 11462 18528
rect 11526 18464 11542 18528
rect 11606 18464 11614 18528
rect 11294 18463 11614 18464
rect 18194 18528 18514 18529
rect 18194 18464 18202 18528
rect 18266 18464 18282 18528
rect 18346 18464 18362 18528
rect 18426 18464 18442 18528
rect 18506 18464 18514 18528
rect 18194 18463 18514 18464
rect 7844 17984 8164 17985
rect 7844 17920 7852 17984
rect 7916 17920 7932 17984
rect 7996 17920 8012 17984
rect 8076 17920 8092 17984
rect 8156 17920 8164 17984
rect 7844 17919 8164 17920
rect 14744 17984 15064 17985
rect 14744 17920 14752 17984
rect 14816 17920 14832 17984
rect 14896 17920 14912 17984
rect 14976 17920 14992 17984
rect 15056 17920 15064 17984
rect 14744 17919 15064 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 20621 17778 20687 17781
rect 22179 17778 22979 17808
rect 20621 17776 22979 17778
rect 20621 17720 20626 17776
rect 20682 17720 22979 17776
rect 20621 17718 22979 17720
rect 20621 17715 20687 17718
rect 22179 17688 22979 17718
rect 4394 17440 4714 17441
rect 4394 17376 4402 17440
rect 4466 17376 4482 17440
rect 4546 17376 4562 17440
rect 4626 17376 4642 17440
rect 4706 17376 4714 17440
rect 4394 17375 4714 17376
rect 11294 17440 11614 17441
rect 11294 17376 11302 17440
rect 11366 17376 11382 17440
rect 11446 17376 11462 17440
rect 11526 17376 11542 17440
rect 11606 17376 11614 17440
rect 11294 17375 11614 17376
rect 18194 17440 18514 17441
rect 18194 17376 18202 17440
rect 18266 17376 18282 17440
rect 18346 17376 18362 17440
rect 18426 17376 18442 17440
rect 18506 17376 18514 17440
rect 18194 17375 18514 17376
rect 7844 16896 8164 16897
rect 7844 16832 7852 16896
rect 7916 16832 7932 16896
rect 7996 16832 8012 16896
rect 8076 16832 8092 16896
rect 8156 16832 8164 16896
rect 7844 16831 8164 16832
rect 14744 16896 15064 16897
rect 14744 16832 14752 16896
rect 14816 16832 14832 16896
rect 14896 16832 14912 16896
rect 14976 16832 14992 16896
rect 15056 16832 15064 16896
rect 14744 16831 15064 16832
rect 4394 16352 4714 16353
rect 4394 16288 4402 16352
rect 4466 16288 4482 16352
rect 4546 16288 4562 16352
rect 4626 16288 4642 16352
rect 4706 16288 4714 16352
rect 4394 16287 4714 16288
rect 11294 16352 11614 16353
rect 11294 16288 11302 16352
rect 11366 16288 11382 16352
rect 11446 16288 11462 16352
rect 11526 16288 11542 16352
rect 11606 16288 11614 16352
rect 11294 16287 11614 16288
rect 18194 16352 18514 16353
rect 18194 16288 18202 16352
rect 18266 16288 18282 16352
rect 18346 16288 18362 16352
rect 18426 16288 18442 16352
rect 18506 16288 18514 16352
rect 18194 16287 18514 16288
rect 7844 15808 8164 15809
rect 0 15738 800 15768
rect 7844 15744 7852 15808
rect 7916 15744 7932 15808
rect 7996 15744 8012 15808
rect 8076 15744 8092 15808
rect 8156 15744 8164 15808
rect 7844 15743 8164 15744
rect 14744 15808 15064 15809
rect 14744 15744 14752 15808
rect 14816 15744 14832 15808
rect 14896 15744 14912 15808
rect 14976 15744 14992 15808
rect 15056 15744 15064 15808
rect 14744 15743 15064 15744
rect 1393 15738 1459 15741
rect 0 15736 1459 15738
rect 0 15680 1398 15736
rect 1454 15680 1459 15736
rect 0 15678 1459 15680
rect 0 15648 800 15678
rect 1393 15675 1459 15678
rect 21081 15738 21147 15741
rect 22179 15738 22979 15768
rect 21081 15736 22979 15738
rect 21081 15680 21086 15736
rect 21142 15680 22979 15736
rect 21081 15678 22979 15680
rect 21081 15675 21147 15678
rect 22179 15648 22979 15678
rect 4394 15264 4714 15265
rect 4394 15200 4402 15264
rect 4466 15200 4482 15264
rect 4546 15200 4562 15264
rect 4626 15200 4642 15264
rect 4706 15200 4714 15264
rect 4394 15199 4714 15200
rect 11294 15264 11614 15265
rect 11294 15200 11302 15264
rect 11366 15200 11382 15264
rect 11446 15200 11462 15264
rect 11526 15200 11542 15264
rect 11606 15200 11614 15264
rect 11294 15199 11614 15200
rect 18194 15264 18514 15265
rect 18194 15200 18202 15264
rect 18266 15200 18282 15264
rect 18346 15200 18362 15264
rect 18426 15200 18442 15264
rect 18506 15200 18514 15264
rect 18194 15199 18514 15200
rect 14641 15058 14707 15061
rect 15285 15058 15351 15061
rect 14641 15056 15351 15058
rect 14641 15000 14646 15056
rect 14702 15000 15290 15056
rect 15346 15000 15351 15056
rect 14641 14998 15351 15000
rect 14641 14995 14707 14998
rect 15285 14995 15351 14998
rect 7844 14720 8164 14721
rect 7844 14656 7852 14720
rect 7916 14656 7932 14720
rect 7996 14656 8012 14720
rect 8076 14656 8092 14720
rect 8156 14656 8164 14720
rect 7844 14655 8164 14656
rect 14744 14720 15064 14721
rect 14744 14656 14752 14720
rect 14816 14656 14832 14720
rect 14896 14656 14912 14720
rect 14976 14656 14992 14720
rect 15056 14656 15064 14720
rect 14744 14655 15064 14656
rect 15285 14514 15351 14517
rect 19241 14514 19307 14517
rect 15285 14512 19307 14514
rect 15285 14456 15290 14512
rect 15346 14456 19246 14512
rect 19302 14456 19307 14512
rect 15285 14454 19307 14456
rect 15285 14451 15351 14454
rect 19241 14451 19307 14454
rect 4394 14176 4714 14177
rect 4394 14112 4402 14176
rect 4466 14112 4482 14176
rect 4546 14112 4562 14176
rect 4626 14112 4642 14176
rect 4706 14112 4714 14176
rect 4394 14111 4714 14112
rect 11294 14176 11614 14177
rect 11294 14112 11302 14176
rect 11366 14112 11382 14176
rect 11446 14112 11462 14176
rect 11526 14112 11542 14176
rect 11606 14112 11614 14176
rect 11294 14111 11614 14112
rect 18194 14176 18514 14177
rect 18194 14112 18202 14176
rect 18266 14112 18282 14176
rect 18346 14112 18362 14176
rect 18426 14112 18442 14176
rect 18506 14112 18514 14176
rect 18194 14111 18514 14112
rect 7844 13632 8164 13633
rect 7844 13568 7852 13632
rect 7916 13568 7932 13632
rect 7996 13568 8012 13632
rect 8076 13568 8092 13632
rect 8156 13568 8164 13632
rect 7844 13567 8164 13568
rect 14744 13632 15064 13633
rect 14744 13568 14752 13632
rect 14816 13568 14832 13632
rect 14896 13568 14912 13632
rect 14976 13568 14992 13632
rect 15056 13568 15064 13632
rect 14744 13567 15064 13568
rect 4394 13088 4714 13089
rect 0 13018 800 13048
rect 4394 13024 4402 13088
rect 4466 13024 4482 13088
rect 4546 13024 4562 13088
rect 4626 13024 4642 13088
rect 4706 13024 4714 13088
rect 4394 13023 4714 13024
rect 11294 13088 11614 13089
rect 11294 13024 11302 13088
rect 11366 13024 11382 13088
rect 11446 13024 11462 13088
rect 11526 13024 11542 13088
rect 11606 13024 11614 13088
rect 11294 13023 11614 13024
rect 18194 13088 18514 13089
rect 18194 13024 18202 13088
rect 18266 13024 18282 13088
rect 18346 13024 18362 13088
rect 18426 13024 18442 13088
rect 18506 13024 18514 13088
rect 18194 13023 18514 13024
rect 1485 13018 1551 13021
rect 0 13016 1551 13018
rect 0 12960 1490 13016
rect 1546 12960 1551 13016
rect 0 12958 1551 12960
rect 0 12928 800 12958
rect 1485 12955 1551 12958
rect 21081 13018 21147 13021
rect 22179 13018 22979 13048
rect 21081 13016 22979 13018
rect 21081 12960 21086 13016
rect 21142 12960 22979 13016
rect 21081 12958 22979 12960
rect 21081 12955 21147 12958
rect 22179 12928 22979 12958
rect 7844 12544 8164 12545
rect 7844 12480 7852 12544
rect 7916 12480 7932 12544
rect 7996 12480 8012 12544
rect 8076 12480 8092 12544
rect 8156 12480 8164 12544
rect 7844 12479 8164 12480
rect 14744 12544 15064 12545
rect 14744 12480 14752 12544
rect 14816 12480 14832 12544
rect 14896 12480 14912 12544
rect 14976 12480 14992 12544
rect 15056 12480 15064 12544
rect 14744 12479 15064 12480
rect 4394 12000 4714 12001
rect 4394 11936 4402 12000
rect 4466 11936 4482 12000
rect 4546 11936 4562 12000
rect 4626 11936 4642 12000
rect 4706 11936 4714 12000
rect 4394 11935 4714 11936
rect 11294 12000 11614 12001
rect 11294 11936 11302 12000
rect 11366 11936 11382 12000
rect 11446 11936 11462 12000
rect 11526 11936 11542 12000
rect 11606 11936 11614 12000
rect 11294 11935 11614 11936
rect 18194 12000 18514 12001
rect 18194 11936 18202 12000
rect 18266 11936 18282 12000
rect 18346 11936 18362 12000
rect 18426 11936 18442 12000
rect 18506 11936 18514 12000
rect 18194 11935 18514 11936
rect 7844 11456 8164 11457
rect 7844 11392 7852 11456
rect 7916 11392 7932 11456
rect 7996 11392 8012 11456
rect 8076 11392 8092 11456
rect 8156 11392 8164 11456
rect 7844 11391 8164 11392
rect 14744 11456 15064 11457
rect 14744 11392 14752 11456
rect 14816 11392 14832 11456
rect 14896 11392 14912 11456
rect 14976 11392 14992 11456
rect 15056 11392 15064 11456
rect 14744 11391 15064 11392
rect 4394 10912 4714 10913
rect 4394 10848 4402 10912
rect 4466 10848 4482 10912
rect 4546 10848 4562 10912
rect 4626 10848 4642 10912
rect 4706 10848 4714 10912
rect 4394 10847 4714 10848
rect 11294 10912 11614 10913
rect 11294 10848 11302 10912
rect 11366 10848 11382 10912
rect 11446 10848 11462 10912
rect 11526 10848 11542 10912
rect 11606 10848 11614 10912
rect 11294 10847 11614 10848
rect 18194 10912 18514 10913
rect 18194 10848 18202 10912
rect 18266 10848 18282 10912
rect 18346 10848 18362 10912
rect 18426 10848 18442 10912
rect 18506 10848 18514 10912
rect 18194 10847 18514 10848
rect 7844 10368 8164 10369
rect 0 10298 800 10328
rect 7844 10304 7852 10368
rect 7916 10304 7932 10368
rect 7996 10304 8012 10368
rect 8076 10304 8092 10368
rect 8156 10304 8164 10368
rect 7844 10303 8164 10304
rect 14744 10368 15064 10369
rect 14744 10304 14752 10368
rect 14816 10304 14832 10368
rect 14896 10304 14912 10368
rect 14976 10304 14992 10368
rect 15056 10304 15064 10368
rect 14744 10303 15064 10304
rect 1485 10298 1551 10301
rect 0 10296 1551 10298
rect 0 10240 1490 10296
rect 1546 10240 1551 10296
rect 0 10238 1551 10240
rect 0 10208 800 10238
rect 1485 10235 1551 10238
rect 21081 10298 21147 10301
rect 22179 10298 22979 10328
rect 21081 10296 22979 10298
rect 21081 10240 21086 10296
rect 21142 10240 22979 10296
rect 21081 10238 22979 10240
rect 21081 10235 21147 10238
rect 22179 10208 22979 10238
rect 4394 9824 4714 9825
rect 4394 9760 4402 9824
rect 4466 9760 4482 9824
rect 4546 9760 4562 9824
rect 4626 9760 4642 9824
rect 4706 9760 4714 9824
rect 4394 9759 4714 9760
rect 11294 9824 11614 9825
rect 11294 9760 11302 9824
rect 11366 9760 11382 9824
rect 11446 9760 11462 9824
rect 11526 9760 11542 9824
rect 11606 9760 11614 9824
rect 11294 9759 11614 9760
rect 18194 9824 18514 9825
rect 18194 9760 18202 9824
rect 18266 9760 18282 9824
rect 18346 9760 18362 9824
rect 18426 9760 18442 9824
rect 18506 9760 18514 9824
rect 18194 9759 18514 9760
rect 7844 9280 8164 9281
rect 7844 9216 7852 9280
rect 7916 9216 7932 9280
rect 7996 9216 8012 9280
rect 8076 9216 8092 9280
rect 8156 9216 8164 9280
rect 7844 9215 8164 9216
rect 14744 9280 15064 9281
rect 14744 9216 14752 9280
rect 14816 9216 14832 9280
rect 14896 9216 14912 9280
rect 14976 9216 14992 9280
rect 15056 9216 15064 9280
rect 14744 9215 15064 9216
rect 4394 8736 4714 8737
rect 4394 8672 4402 8736
rect 4466 8672 4482 8736
rect 4546 8672 4562 8736
rect 4626 8672 4642 8736
rect 4706 8672 4714 8736
rect 4394 8671 4714 8672
rect 11294 8736 11614 8737
rect 11294 8672 11302 8736
rect 11366 8672 11382 8736
rect 11446 8672 11462 8736
rect 11526 8672 11542 8736
rect 11606 8672 11614 8736
rect 11294 8671 11614 8672
rect 18194 8736 18514 8737
rect 18194 8672 18202 8736
rect 18266 8672 18282 8736
rect 18346 8672 18362 8736
rect 18426 8672 18442 8736
rect 18506 8672 18514 8736
rect 18194 8671 18514 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 21081 8258 21147 8261
rect 22179 8258 22979 8288
rect 21081 8256 22979 8258
rect 21081 8200 21086 8256
rect 21142 8200 22979 8256
rect 21081 8198 22979 8200
rect 21081 8195 21147 8198
rect 7844 8192 8164 8193
rect 7844 8128 7852 8192
rect 7916 8128 7932 8192
rect 7996 8128 8012 8192
rect 8076 8128 8092 8192
rect 8156 8128 8164 8192
rect 7844 8127 8164 8128
rect 14744 8192 15064 8193
rect 14744 8128 14752 8192
rect 14816 8128 14832 8192
rect 14896 8128 14912 8192
rect 14976 8128 14992 8192
rect 15056 8128 15064 8192
rect 22179 8168 22979 8198
rect 14744 8127 15064 8128
rect 4394 7648 4714 7649
rect 4394 7584 4402 7648
rect 4466 7584 4482 7648
rect 4546 7584 4562 7648
rect 4626 7584 4642 7648
rect 4706 7584 4714 7648
rect 4394 7583 4714 7584
rect 11294 7648 11614 7649
rect 11294 7584 11302 7648
rect 11366 7584 11382 7648
rect 11446 7584 11462 7648
rect 11526 7584 11542 7648
rect 11606 7584 11614 7648
rect 11294 7583 11614 7584
rect 18194 7648 18514 7649
rect 18194 7584 18202 7648
rect 18266 7584 18282 7648
rect 18346 7584 18362 7648
rect 18426 7584 18442 7648
rect 18506 7584 18514 7648
rect 18194 7583 18514 7584
rect 7844 7104 8164 7105
rect 7844 7040 7852 7104
rect 7916 7040 7932 7104
rect 7996 7040 8012 7104
rect 8076 7040 8092 7104
rect 8156 7040 8164 7104
rect 7844 7039 8164 7040
rect 14744 7104 15064 7105
rect 14744 7040 14752 7104
rect 14816 7040 14832 7104
rect 14896 7040 14912 7104
rect 14976 7040 14992 7104
rect 15056 7040 15064 7104
rect 14744 7039 15064 7040
rect 4394 6560 4714 6561
rect 4394 6496 4402 6560
rect 4466 6496 4482 6560
rect 4546 6496 4562 6560
rect 4626 6496 4642 6560
rect 4706 6496 4714 6560
rect 4394 6495 4714 6496
rect 11294 6560 11614 6561
rect 11294 6496 11302 6560
rect 11366 6496 11382 6560
rect 11446 6496 11462 6560
rect 11526 6496 11542 6560
rect 11606 6496 11614 6560
rect 11294 6495 11614 6496
rect 18194 6560 18514 6561
rect 18194 6496 18202 6560
rect 18266 6496 18282 6560
rect 18346 6496 18362 6560
rect 18426 6496 18442 6560
rect 18506 6496 18514 6560
rect 18194 6495 18514 6496
rect 7844 6016 8164 6017
rect 7844 5952 7852 6016
rect 7916 5952 7932 6016
rect 7996 5952 8012 6016
rect 8076 5952 8092 6016
rect 8156 5952 8164 6016
rect 7844 5951 8164 5952
rect 14744 6016 15064 6017
rect 14744 5952 14752 6016
rect 14816 5952 14832 6016
rect 14896 5952 14912 6016
rect 14976 5952 14992 6016
rect 15056 5952 15064 6016
rect 14744 5951 15064 5952
rect 0 5538 800 5568
rect 1485 5538 1551 5541
rect 0 5536 1551 5538
rect 0 5480 1490 5536
rect 1546 5480 1551 5536
rect 0 5478 1551 5480
rect 0 5448 800 5478
rect 1485 5475 1551 5478
rect 21081 5538 21147 5541
rect 22179 5538 22979 5568
rect 21081 5536 22979 5538
rect 21081 5480 21086 5536
rect 21142 5480 22979 5536
rect 21081 5478 22979 5480
rect 21081 5475 21147 5478
rect 4394 5472 4714 5473
rect 4394 5408 4402 5472
rect 4466 5408 4482 5472
rect 4546 5408 4562 5472
rect 4626 5408 4642 5472
rect 4706 5408 4714 5472
rect 4394 5407 4714 5408
rect 11294 5472 11614 5473
rect 11294 5408 11302 5472
rect 11366 5408 11382 5472
rect 11446 5408 11462 5472
rect 11526 5408 11542 5472
rect 11606 5408 11614 5472
rect 11294 5407 11614 5408
rect 18194 5472 18514 5473
rect 18194 5408 18202 5472
rect 18266 5408 18282 5472
rect 18346 5408 18362 5472
rect 18426 5408 18442 5472
rect 18506 5408 18514 5472
rect 22179 5448 22979 5478
rect 18194 5407 18514 5408
rect 7844 4928 8164 4929
rect 7844 4864 7852 4928
rect 7916 4864 7932 4928
rect 7996 4864 8012 4928
rect 8076 4864 8092 4928
rect 8156 4864 8164 4928
rect 7844 4863 8164 4864
rect 14744 4928 15064 4929
rect 14744 4864 14752 4928
rect 14816 4864 14832 4928
rect 14896 4864 14912 4928
rect 14976 4864 14992 4928
rect 15056 4864 15064 4928
rect 14744 4863 15064 4864
rect 4394 4384 4714 4385
rect 4394 4320 4402 4384
rect 4466 4320 4482 4384
rect 4546 4320 4562 4384
rect 4626 4320 4642 4384
rect 4706 4320 4714 4384
rect 4394 4319 4714 4320
rect 11294 4384 11614 4385
rect 11294 4320 11302 4384
rect 11366 4320 11382 4384
rect 11446 4320 11462 4384
rect 11526 4320 11542 4384
rect 11606 4320 11614 4384
rect 11294 4319 11614 4320
rect 18194 4384 18514 4385
rect 18194 4320 18202 4384
rect 18266 4320 18282 4384
rect 18346 4320 18362 4384
rect 18426 4320 18442 4384
rect 18506 4320 18514 4384
rect 18194 4319 18514 4320
rect 7844 3840 8164 3841
rect 7844 3776 7852 3840
rect 7916 3776 7932 3840
rect 7996 3776 8012 3840
rect 8076 3776 8092 3840
rect 8156 3776 8164 3840
rect 7844 3775 8164 3776
rect 14744 3840 15064 3841
rect 14744 3776 14752 3840
rect 14816 3776 14832 3840
rect 14896 3776 14912 3840
rect 14976 3776 14992 3840
rect 15056 3776 15064 3840
rect 14744 3775 15064 3776
rect 4394 3296 4714 3297
rect 4394 3232 4402 3296
rect 4466 3232 4482 3296
rect 4546 3232 4562 3296
rect 4626 3232 4642 3296
rect 4706 3232 4714 3296
rect 4394 3231 4714 3232
rect 11294 3296 11614 3297
rect 11294 3232 11302 3296
rect 11366 3232 11382 3296
rect 11446 3232 11462 3296
rect 11526 3232 11542 3296
rect 11606 3232 11614 3296
rect 11294 3231 11614 3232
rect 18194 3296 18514 3297
rect 18194 3232 18202 3296
rect 18266 3232 18282 3296
rect 18346 3232 18362 3296
rect 18426 3232 18442 3296
rect 18506 3232 18514 3296
rect 18194 3231 18514 3232
rect 0 2818 800 2848
rect 1393 2818 1459 2821
rect 0 2816 1459 2818
rect 0 2760 1398 2816
rect 1454 2760 1459 2816
rect 0 2758 1459 2760
rect 0 2728 800 2758
rect 1393 2755 1459 2758
rect 20069 2818 20135 2821
rect 22179 2818 22979 2848
rect 20069 2816 22979 2818
rect 20069 2760 20074 2816
rect 20130 2760 22979 2816
rect 20069 2758 22979 2760
rect 20069 2755 20135 2758
rect 7844 2752 8164 2753
rect 7844 2688 7852 2752
rect 7916 2688 7932 2752
rect 7996 2688 8012 2752
rect 8076 2688 8092 2752
rect 8156 2688 8164 2752
rect 7844 2687 8164 2688
rect 14744 2752 15064 2753
rect 14744 2688 14752 2752
rect 14816 2688 14832 2752
rect 14896 2688 14912 2752
rect 14976 2688 14992 2752
rect 15056 2688 15064 2752
rect 22179 2728 22979 2758
rect 14744 2687 15064 2688
rect 4394 2208 4714 2209
rect 4394 2144 4402 2208
rect 4466 2144 4482 2208
rect 4546 2144 4562 2208
rect 4626 2144 4642 2208
rect 4706 2144 4714 2208
rect 4394 2143 4714 2144
rect 11294 2208 11614 2209
rect 11294 2144 11302 2208
rect 11366 2144 11382 2208
rect 11446 2144 11462 2208
rect 11526 2144 11542 2208
rect 11606 2144 11614 2208
rect 11294 2143 11614 2144
rect 18194 2208 18514 2209
rect 18194 2144 18202 2208
rect 18266 2144 18282 2208
rect 18346 2144 18362 2208
rect 18426 2144 18442 2208
rect 18506 2144 18514 2208
rect 18194 2143 18514 2144
<< via3 >>
rect 4402 22876 4466 22880
rect 4402 22820 4406 22876
rect 4406 22820 4462 22876
rect 4462 22820 4466 22876
rect 4402 22816 4466 22820
rect 4482 22876 4546 22880
rect 4482 22820 4486 22876
rect 4486 22820 4542 22876
rect 4542 22820 4546 22876
rect 4482 22816 4546 22820
rect 4562 22876 4626 22880
rect 4562 22820 4566 22876
rect 4566 22820 4622 22876
rect 4622 22820 4626 22876
rect 4562 22816 4626 22820
rect 4642 22876 4706 22880
rect 4642 22820 4646 22876
rect 4646 22820 4702 22876
rect 4702 22820 4706 22876
rect 4642 22816 4706 22820
rect 11302 22876 11366 22880
rect 11302 22820 11306 22876
rect 11306 22820 11362 22876
rect 11362 22820 11366 22876
rect 11302 22816 11366 22820
rect 11382 22876 11446 22880
rect 11382 22820 11386 22876
rect 11386 22820 11442 22876
rect 11442 22820 11446 22876
rect 11382 22816 11446 22820
rect 11462 22876 11526 22880
rect 11462 22820 11466 22876
rect 11466 22820 11522 22876
rect 11522 22820 11526 22876
rect 11462 22816 11526 22820
rect 11542 22876 11606 22880
rect 11542 22820 11546 22876
rect 11546 22820 11602 22876
rect 11602 22820 11606 22876
rect 11542 22816 11606 22820
rect 18202 22876 18266 22880
rect 18202 22820 18206 22876
rect 18206 22820 18262 22876
rect 18262 22820 18266 22876
rect 18202 22816 18266 22820
rect 18282 22876 18346 22880
rect 18282 22820 18286 22876
rect 18286 22820 18342 22876
rect 18342 22820 18346 22876
rect 18282 22816 18346 22820
rect 18362 22876 18426 22880
rect 18362 22820 18366 22876
rect 18366 22820 18422 22876
rect 18422 22820 18426 22876
rect 18362 22816 18426 22820
rect 18442 22876 18506 22880
rect 18442 22820 18446 22876
rect 18446 22820 18502 22876
rect 18502 22820 18506 22876
rect 18442 22816 18506 22820
rect 7852 22332 7916 22336
rect 7852 22276 7856 22332
rect 7856 22276 7912 22332
rect 7912 22276 7916 22332
rect 7852 22272 7916 22276
rect 7932 22332 7996 22336
rect 7932 22276 7936 22332
rect 7936 22276 7992 22332
rect 7992 22276 7996 22332
rect 7932 22272 7996 22276
rect 8012 22332 8076 22336
rect 8012 22276 8016 22332
rect 8016 22276 8072 22332
rect 8072 22276 8076 22332
rect 8012 22272 8076 22276
rect 8092 22332 8156 22336
rect 8092 22276 8096 22332
rect 8096 22276 8152 22332
rect 8152 22276 8156 22332
rect 8092 22272 8156 22276
rect 14752 22332 14816 22336
rect 14752 22276 14756 22332
rect 14756 22276 14812 22332
rect 14812 22276 14816 22332
rect 14752 22272 14816 22276
rect 14832 22332 14896 22336
rect 14832 22276 14836 22332
rect 14836 22276 14892 22332
rect 14892 22276 14896 22332
rect 14832 22272 14896 22276
rect 14912 22332 14976 22336
rect 14912 22276 14916 22332
rect 14916 22276 14972 22332
rect 14972 22276 14976 22332
rect 14912 22272 14976 22276
rect 14992 22332 15056 22336
rect 14992 22276 14996 22332
rect 14996 22276 15052 22332
rect 15052 22276 15056 22332
rect 14992 22272 15056 22276
rect 4402 21788 4466 21792
rect 4402 21732 4406 21788
rect 4406 21732 4462 21788
rect 4462 21732 4466 21788
rect 4402 21728 4466 21732
rect 4482 21788 4546 21792
rect 4482 21732 4486 21788
rect 4486 21732 4542 21788
rect 4542 21732 4546 21788
rect 4482 21728 4546 21732
rect 4562 21788 4626 21792
rect 4562 21732 4566 21788
rect 4566 21732 4622 21788
rect 4622 21732 4626 21788
rect 4562 21728 4626 21732
rect 4642 21788 4706 21792
rect 4642 21732 4646 21788
rect 4646 21732 4702 21788
rect 4702 21732 4706 21788
rect 4642 21728 4706 21732
rect 11302 21788 11366 21792
rect 11302 21732 11306 21788
rect 11306 21732 11362 21788
rect 11362 21732 11366 21788
rect 11302 21728 11366 21732
rect 11382 21788 11446 21792
rect 11382 21732 11386 21788
rect 11386 21732 11442 21788
rect 11442 21732 11446 21788
rect 11382 21728 11446 21732
rect 11462 21788 11526 21792
rect 11462 21732 11466 21788
rect 11466 21732 11522 21788
rect 11522 21732 11526 21788
rect 11462 21728 11526 21732
rect 11542 21788 11606 21792
rect 11542 21732 11546 21788
rect 11546 21732 11602 21788
rect 11602 21732 11606 21788
rect 11542 21728 11606 21732
rect 18202 21788 18266 21792
rect 18202 21732 18206 21788
rect 18206 21732 18262 21788
rect 18262 21732 18266 21788
rect 18202 21728 18266 21732
rect 18282 21788 18346 21792
rect 18282 21732 18286 21788
rect 18286 21732 18342 21788
rect 18342 21732 18346 21788
rect 18282 21728 18346 21732
rect 18362 21788 18426 21792
rect 18362 21732 18366 21788
rect 18366 21732 18422 21788
rect 18422 21732 18426 21788
rect 18362 21728 18426 21732
rect 18442 21788 18506 21792
rect 18442 21732 18446 21788
rect 18446 21732 18502 21788
rect 18502 21732 18506 21788
rect 18442 21728 18506 21732
rect 7852 21244 7916 21248
rect 7852 21188 7856 21244
rect 7856 21188 7912 21244
rect 7912 21188 7916 21244
rect 7852 21184 7916 21188
rect 7932 21244 7996 21248
rect 7932 21188 7936 21244
rect 7936 21188 7992 21244
rect 7992 21188 7996 21244
rect 7932 21184 7996 21188
rect 8012 21244 8076 21248
rect 8012 21188 8016 21244
rect 8016 21188 8072 21244
rect 8072 21188 8076 21244
rect 8012 21184 8076 21188
rect 8092 21244 8156 21248
rect 8092 21188 8096 21244
rect 8096 21188 8152 21244
rect 8152 21188 8156 21244
rect 8092 21184 8156 21188
rect 14752 21244 14816 21248
rect 14752 21188 14756 21244
rect 14756 21188 14812 21244
rect 14812 21188 14816 21244
rect 14752 21184 14816 21188
rect 14832 21244 14896 21248
rect 14832 21188 14836 21244
rect 14836 21188 14892 21244
rect 14892 21188 14896 21244
rect 14832 21184 14896 21188
rect 14912 21244 14976 21248
rect 14912 21188 14916 21244
rect 14916 21188 14972 21244
rect 14972 21188 14976 21244
rect 14912 21184 14976 21188
rect 14992 21244 15056 21248
rect 14992 21188 14996 21244
rect 14996 21188 15052 21244
rect 15052 21188 15056 21244
rect 14992 21184 15056 21188
rect 4402 20700 4466 20704
rect 4402 20644 4406 20700
rect 4406 20644 4462 20700
rect 4462 20644 4466 20700
rect 4402 20640 4466 20644
rect 4482 20700 4546 20704
rect 4482 20644 4486 20700
rect 4486 20644 4542 20700
rect 4542 20644 4546 20700
rect 4482 20640 4546 20644
rect 4562 20700 4626 20704
rect 4562 20644 4566 20700
rect 4566 20644 4622 20700
rect 4622 20644 4626 20700
rect 4562 20640 4626 20644
rect 4642 20700 4706 20704
rect 4642 20644 4646 20700
rect 4646 20644 4702 20700
rect 4702 20644 4706 20700
rect 4642 20640 4706 20644
rect 11302 20700 11366 20704
rect 11302 20644 11306 20700
rect 11306 20644 11362 20700
rect 11362 20644 11366 20700
rect 11302 20640 11366 20644
rect 11382 20700 11446 20704
rect 11382 20644 11386 20700
rect 11386 20644 11442 20700
rect 11442 20644 11446 20700
rect 11382 20640 11446 20644
rect 11462 20700 11526 20704
rect 11462 20644 11466 20700
rect 11466 20644 11522 20700
rect 11522 20644 11526 20700
rect 11462 20640 11526 20644
rect 11542 20700 11606 20704
rect 11542 20644 11546 20700
rect 11546 20644 11602 20700
rect 11602 20644 11606 20700
rect 11542 20640 11606 20644
rect 18202 20700 18266 20704
rect 18202 20644 18206 20700
rect 18206 20644 18262 20700
rect 18262 20644 18266 20700
rect 18202 20640 18266 20644
rect 18282 20700 18346 20704
rect 18282 20644 18286 20700
rect 18286 20644 18342 20700
rect 18342 20644 18346 20700
rect 18282 20640 18346 20644
rect 18362 20700 18426 20704
rect 18362 20644 18366 20700
rect 18366 20644 18422 20700
rect 18422 20644 18426 20700
rect 18362 20640 18426 20644
rect 18442 20700 18506 20704
rect 18442 20644 18446 20700
rect 18446 20644 18502 20700
rect 18502 20644 18506 20700
rect 18442 20640 18506 20644
rect 7852 20156 7916 20160
rect 7852 20100 7856 20156
rect 7856 20100 7912 20156
rect 7912 20100 7916 20156
rect 7852 20096 7916 20100
rect 7932 20156 7996 20160
rect 7932 20100 7936 20156
rect 7936 20100 7992 20156
rect 7992 20100 7996 20156
rect 7932 20096 7996 20100
rect 8012 20156 8076 20160
rect 8012 20100 8016 20156
rect 8016 20100 8072 20156
rect 8072 20100 8076 20156
rect 8012 20096 8076 20100
rect 8092 20156 8156 20160
rect 8092 20100 8096 20156
rect 8096 20100 8152 20156
rect 8152 20100 8156 20156
rect 8092 20096 8156 20100
rect 14752 20156 14816 20160
rect 14752 20100 14756 20156
rect 14756 20100 14812 20156
rect 14812 20100 14816 20156
rect 14752 20096 14816 20100
rect 14832 20156 14896 20160
rect 14832 20100 14836 20156
rect 14836 20100 14892 20156
rect 14892 20100 14896 20156
rect 14832 20096 14896 20100
rect 14912 20156 14976 20160
rect 14912 20100 14916 20156
rect 14916 20100 14972 20156
rect 14972 20100 14976 20156
rect 14912 20096 14976 20100
rect 14992 20156 15056 20160
rect 14992 20100 14996 20156
rect 14996 20100 15052 20156
rect 15052 20100 15056 20156
rect 14992 20096 15056 20100
rect 4402 19612 4466 19616
rect 4402 19556 4406 19612
rect 4406 19556 4462 19612
rect 4462 19556 4466 19612
rect 4402 19552 4466 19556
rect 4482 19612 4546 19616
rect 4482 19556 4486 19612
rect 4486 19556 4542 19612
rect 4542 19556 4546 19612
rect 4482 19552 4546 19556
rect 4562 19612 4626 19616
rect 4562 19556 4566 19612
rect 4566 19556 4622 19612
rect 4622 19556 4626 19612
rect 4562 19552 4626 19556
rect 4642 19612 4706 19616
rect 4642 19556 4646 19612
rect 4646 19556 4702 19612
rect 4702 19556 4706 19612
rect 4642 19552 4706 19556
rect 11302 19612 11366 19616
rect 11302 19556 11306 19612
rect 11306 19556 11362 19612
rect 11362 19556 11366 19612
rect 11302 19552 11366 19556
rect 11382 19612 11446 19616
rect 11382 19556 11386 19612
rect 11386 19556 11442 19612
rect 11442 19556 11446 19612
rect 11382 19552 11446 19556
rect 11462 19612 11526 19616
rect 11462 19556 11466 19612
rect 11466 19556 11522 19612
rect 11522 19556 11526 19612
rect 11462 19552 11526 19556
rect 11542 19612 11606 19616
rect 11542 19556 11546 19612
rect 11546 19556 11602 19612
rect 11602 19556 11606 19612
rect 11542 19552 11606 19556
rect 18202 19612 18266 19616
rect 18202 19556 18206 19612
rect 18206 19556 18262 19612
rect 18262 19556 18266 19612
rect 18202 19552 18266 19556
rect 18282 19612 18346 19616
rect 18282 19556 18286 19612
rect 18286 19556 18342 19612
rect 18342 19556 18346 19612
rect 18282 19552 18346 19556
rect 18362 19612 18426 19616
rect 18362 19556 18366 19612
rect 18366 19556 18422 19612
rect 18422 19556 18426 19612
rect 18362 19552 18426 19556
rect 18442 19612 18506 19616
rect 18442 19556 18446 19612
rect 18446 19556 18502 19612
rect 18502 19556 18506 19612
rect 18442 19552 18506 19556
rect 7852 19068 7916 19072
rect 7852 19012 7856 19068
rect 7856 19012 7912 19068
rect 7912 19012 7916 19068
rect 7852 19008 7916 19012
rect 7932 19068 7996 19072
rect 7932 19012 7936 19068
rect 7936 19012 7992 19068
rect 7992 19012 7996 19068
rect 7932 19008 7996 19012
rect 8012 19068 8076 19072
rect 8012 19012 8016 19068
rect 8016 19012 8072 19068
rect 8072 19012 8076 19068
rect 8012 19008 8076 19012
rect 8092 19068 8156 19072
rect 8092 19012 8096 19068
rect 8096 19012 8152 19068
rect 8152 19012 8156 19068
rect 8092 19008 8156 19012
rect 14752 19068 14816 19072
rect 14752 19012 14756 19068
rect 14756 19012 14812 19068
rect 14812 19012 14816 19068
rect 14752 19008 14816 19012
rect 14832 19068 14896 19072
rect 14832 19012 14836 19068
rect 14836 19012 14892 19068
rect 14892 19012 14896 19068
rect 14832 19008 14896 19012
rect 14912 19068 14976 19072
rect 14912 19012 14916 19068
rect 14916 19012 14972 19068
rect 14972 19012 14976 19068
rect 14912 19008 14976 19012
rect 14992 19068 15056 19072
rect 14992 19012 14996 19068
rect 14996 19012 15052 19068
rect 15052 19012 15056 19068
rect 14992 19008 15056 19012
rect 4402 18524 4466 18528
rect 4402 18468 4406 18524
rect 4406 18468 4462 18524
rect 4462 18468 4466 18524
rect 4402 18464 4466 18468
rect 4482 18524 4546 18528
rect 4482 18468 4486 18524
rect 4486 18468 4542 18524
rect 4542 18468 4546 18524
rect 4482 18464 4546 18468
rect 4562 18524 4626 18528
rect 4562 18468 4566 18524
rect 4566 18468 4622 18524
rect 4622 18468 4626 18524
rect 4562 18464 4626 18468
rect 4642 18524 4706 18528
rect 4642 18468 4646 18524
rect 4646 18468 4702 18524
rect 4702 18468 4706 18524
rect 4642 18464 4706 18468
rect 11302 18524 11366 18528
rect 11302 18468 11306 18524
rect 11306 18468 11362 18524
rect 11362 18468 11366 18524
rect 11302 18464 11366 18468
rect 11382 18524 11446 18528
rect 11382 18468 11386 18524
rect 11386 18468 11442 18524
rect 11442 18468 11446 18524
rect 11382 18464 11446 18468
rect 11462 18524 11526 18528
rect 11462 18468 11466 18524
rect 11466 18468 11522 18524
rect 11522 18468 11526 18524
rect 11462 18464 11526 18468
rect 11542 18524 11606 18528
rect 11542 18468 11546 18524
rect 11546 18468 11602 18524
rect 11602 18468 11606 18524
rect 11542 18464 11606 18468
rect 18202 18524 18266 18528
rect 18202 18468 18206 18524
rect 18206 18468 18262 18524
rect 18262 18468 18266 18524
rect 18202 18464 18266 18468
rect 18282 18524 18346 18528
rect 18282 18468 18286 18524
rect 18286 18468 18342 18524
rect 18342 18468 18346 18524
rect 18282 18464 18346 18468
rect 18362 18524 18426 18528
rect 18362 18468 18366 18524
rect 18366 18468 18422 18524
rect 18422 18468 18426 18524
rect 18362 18464 18426 18468
rect 18442 18524 18506 18528
rect 18442 18468 18446 18524
rect 18446 18468 18502 18524
rect 18502 18468 18506 18524
rect 18442 18464 18506 18468
rect 7852 17980 7916 17984
rect 7852 17924 7856 17980
rect 7856 17924 7912 17980
rect 7912 17924 7916 17980
rect 7852 17920 7916 17924
rect 7932 17980 7996 17984
rect 7932 17924 7936 17980
rect 7936 17924 7992 17980
rect 7992 17924 7996 17980
rect 7932 17920 7996 17924
rect 8012 17980 8076 17984
rect 8012 17924 8016 17980
rect 8016 17924 8072 17980
rect 8072 17924 8076 17980
rect 8012 17920 8076 17924
rect 8092 17980 8156 17984
rect 8092 17924 8096 17980
rect 8096 17924 8152 17980
rect 8152 17924 8156 17980
rect 8092 17920 8156 17924
rect 14752 17980 14816 17984
rect 14752 17924 14756 17980
rect 14756 17924 14812 17980
rect 14812 17924 14816 17980
rect 14752 17920 14816 17924
rect 14832 17980 14896 17984
rect 14832 17924 14836 17980
rect 14836 17924 14892 17980
rect 14892 17924 14896 17980
rect 14832 17920 14896 17924
rect 14912 17980 14976 17984
rect 14912 17924 14916 17980
rect 14916 17924 14972 17980
rect 14972 17924 14976 17980
rect 14912 17920 14976 17924
rect 14992 17980 15056 17984
rect 14992 17924 14996 17980
rect 14996 17924 15052 17980
rect 15052 17924 15056 17980
rect 14992 17920 15056 17924
rect 4402 17436 4466 17440
rect 4402 17380 4406 17436
rect 4406 17380 4462 17436
rect 4462 17380 4466 17436
rect 4402 17376 4466 17380
rect 4482 17436 4546 17440
rect 4482 17380 4486 17436
rect 4486 17380 4542 17436
rect 4542 17380 4546 17436
rect 4482 17376 4546 17380
rect 4562 17436 4626 17440
rect 4562 17380 4566 17436
rect 4566 17380 4622 17436
rect 4622 17380 4626 17436
rect 4562 17376 4626 17380
rect 4642 17436 4706 17440
rect 4642 17380 4646 17436
rect 4646 17380 4702 17436
rect 4702 17380 4706 17436
rect 4642 17376 4706 17380
rect 11302 17436 11366 17440
rect 11302 17380 11306 17436
rect 11306 17380 11362 17436
rect 11362 17380 11366 17436
rect 11302 17376 11366 17380
rect 11382 17436 11446 17440
rect 11382 17380 11386 17436
rect 11386 17380 11442 17436
rect 11442 17380 11446 17436
rect 11382 17376 11446 17380
rect 11462 17436 11526 17440
rect 11462 17380 11466 17436
rect 11466 17380 11522 17436
rect 11522 17380 11526 17436
rect 11462 17376 11526 17380
rect 11542 17436 11606 17440
rect 11542 17380 11546 17436
rect 11546 17380 11602 17436
rect 11602 17380 11606 17436
rect 11542 17376 11606 17380
rect 18202 17436 18266 17440
rect 18202 17380 18206 17436
rect 18206 17380 18262 17436
rect 18262 17380 18266 17436
rect 18202 17376 18266 17380
rect 18282 17436 18346 17440
rect 18282 17380 18286 17436
rect 18286 17380 18342 17436
rect 18342 17380 18346 17436
rect 18282 17376 18346 17380
rect 18362 17436 18426 17440
rect 18362 17380 18366 17436
rect 18366 17380 18422 17436
rect 18422 17380 18426 17436
rect 18362 17376 18426 17380
rect 18442 17436 18506 17440
rect 18442 17380 18446 17436
rect 18446 17380 18502 17436
rect 18502 17380 18506 17436
rect 18442 17376 18506 17380
rect 7852 16892 7916 16896
rect 7852 16836 7856 16892
rect 7856 16836 7912 16892
rect 7912 16836 7916 16892
rect 7852 16832 7916 16836
rect 7932 16892 7996 16896
rect 7932 16836 7936 16892
rect 7936 16836 7992 16892
rect 7992 16836 7996 16892
rect 7932 16832 7996 16836
rect 8012 16892 8076 16896
rect 8012 16836 8016 16892
rect 8016 16836 8072 16892
rect 8072 16836 8076 16892
rect 8012 16832 8076 16836
rect 8092 16892 8156 16896
rect 8092 16836 8096 16892
rect 8096 16836 8152 16892
rect 8152 16836 8156 16892
rect 8092 16832 8156 16836
rect 14752 16892 14816 16896
rect 14752 16836 14756 16892
rect 14756 16836 14812 16892
rect 14812 16836 14816 16892
rect 14752 16832 14816 16836
rect 14832 16892 14896 16896
rect 14832 16836 14836 16892
rect 14836 16836 14892 16892
rect 14892 16836 14896 16892
rect 14832 16832 14896 16836
rect 14912 16892 14976 16896
rect 14912 16836 14916 16892
rect 14916 16836 14972 16892
rect 14972 16836 14976 16892
rect 14912 16832 14976 16836
rect 14992 16892 15056 16896
rect 14992 16836 14996 16892
rect 14996 16836 15052 16892
rect 15052 16836 15056 16892
rect 14992 16832 15056 16836
rect 4402 16348 4466 16352
rect 4402 16292 4406 16348
rect 4406 16292 4462 16348
rect 4462 16292 4466 16348
rect 4402 16288 4466 16292
rect 4482 16348 4546 16352
rect 4482 16292 4486 16348
rect 4486 16292 4542 16348
rect 4542 16292 4546 16348
rect 4482 16288 4546 16292
rect 4562 16348 4626 16352
rect 4562 16292 4566 16348
rect 4566 16292 4622 16348
rect 4622 16292 4626 16348
rect 4562 16288 4626 16292
rect 4642 16348 4706 16352
rect 4642 16292 4646 16348
rect 4646 16292 4702 16348
rect 4702 16292 4706 16348
rect 4642 16288 4706 16292
rect 11302 16348 11366 16352
rect 11302 16292 11306 16348
rect 11306 16292 11362 16348
rect 11362 16292 11366 16348
rect 11302 16288 11366 16292
rect 11382 16348 11446 16352
rect 11382 16292 11386 16348
rect 11386 16292 11442 16348
rect 11442 16292 11446 16348
rect 11382 16288 11446 16292
rect 11462 16348 11526 16352
rect 11462 16292 11466 16348
rect 11466 16292 11522 16348
rect 11522 16292 11526 16348
rect 11462 16288 11526 16292
rect 11542 16348 11606 16352
rect 11542 16292 11546 16348
rect 11546 16292 11602 16348
rect 11602 16292 11606 16348
rect 11542 16288 11606 16292
rect 18202 16348 18266 16352
rect 18202 16292 18206 16348
rect 18206 16292 18262 16348
rect 18262 16292 18266 16348
rect 18202 16288 18266 16292
rect 18282 16348 18346 16352
rect 18282 16292 18286 16348
rect 18286 16292 18342 16348
rect 18342 16292 18346 16348
rect 18282 16288 18346 16292
rect 18362 16348 18426 16352
rect 18362 16292 18366 16348
rect 18366 16292 18422 16348
rect 18422 16292 18426 16348
rect 18362 16288 18426 16292
rect 18442 16348 18506 16352
rect 18442 16292 18446 16348
rect 18446 16292 18502 16348
rect 18502 16292 18506 16348
rect 18442 16288 18506 16292
rect 7852 15804 7916 15808
rect 7852 15748 7856 15804
rect 7856 15748 7912 15804
rect 7912 15748 7916 15804
rect 7852 15744 7916 15748
rect 7932 15804 7996 15808
rect 7932 15748 7936 15804
rect 7936 15748 7992 15804
rect 7992 15748 7996 15804
rect 7932 15744 7996 15748
rect 8012 15804 8076 15808
rect 8012 15748 8016 15804
rect 8016 15748 8072 15804
rect 8072 15748 8076 15804
rect 8012 15744 8076 15748
rect 8092 15804 8156 15808
rect 8092 15748 8096 15804
rect 8096 15748 8152 15804
rect 8152 15748 8156 15804
rect 8092 15744 8156 15748
rect 14752 15804 14816 15808
rect 14752 15748 14756 15804
rect 14756 15748 14812 15804
rect 14812 15748 14816 15804
rect 14752 15744 14816 15748
rect 14832 15804 14896 15808
rect 14832 15748 14836 15804
rect 14836 15748 14892 15804
rect 14892 15748 14896 15804
rect 14832 15744 14896 15748
rect 14912 15804 14976 15808
rect 14912 15748 14916 15804
rect 14916 15748 14972 15804
rect 14972 15748 14976 15804
rect 14912 15744 14976 15748
rect 14992 15804 15056 15808
rect 14992 15748 14996 15804
rect 14996 15748 15052 15804
rect 15052 15748 15056 15804
rect 14992 15744 15056 15748
rect 4402 15260 4466 15264
rect 4402 15204 4406 15260
rect 4406 15204 4462 15260
rect 4462 15204 4466 15260
rect 4402 15200 4466 15204
rect 4482 15260 4546 15264
rect 4482 15204 4486 15260
rect 4486 15204 4542 15260
rect 4542 15204 4546 15260
rect 4482 15200 4546 15204
rect 4562 15260 4626 15264
rect 4562 15204 4566 15260
rect 4566 15204 4622 15260
rect 4622 15204 4626 15260
rect 4562 15200 4626 15204
rect 4642 15260 4706 15264
rect 4642 15204 4646 15260
rect 4646 15204 4702 15260
rect 4702 15204 4706 15260
rect 4642 15200 4706 15204
rect 11302 15260 11366 15264
rect 11302 15204 11306 15260
rect 11306 15204 11362 15260
rect 11362 15204 11366 15260
rect 11302 15200 11366 15204
rect 11382 15260 11446 15264
rect 11382 15204 11386 15260
rect 11386 15204 11442 15260
rect 11442 15204 11446 15260
rect 11382 15200 11446 15204
rect 11462 15260 11526 15264
rect 11462 15204 11466 15260
rect 11466 15204 11522 15260
rect 11522 15204 11526 15260
rect 11462 15200 11526 15204
rect 11542 15260 11606 15264
rect 11542 15204 11546 15260
rect 11546 15204 11602 15260
rect 11602 15204 11606 15260
rect 11542 15200 11606 15204
rect 18202 15260 18266 15264
rect 18202 15204 18206 15260
rect 18206 15204 18262 15260
rect 18262 15204 18266 15260
rect 18202 15200 18266 15204
rect 18282 15260 18346 15264
rect 18282 15204 18286 15260
rect 18286 15204 18342 15260
rect 18342 15204 18346 15260
rect 18282 15200 18346 15204
rect 18362 15260 18426 15264
rect 18362 15204 18366 15260
rect 18366 15204 18422 15260
rect 18422 15204 18426 15260
rect 18362 15200 18426 15204
rect 18442 15260 18506 15264
rect 18442 15204 18446 15260
rect 18446 15204 18502 15260
rect 18502 15204 18506 15260
rect 18442 15200 18506 15204
rect 7852 14716 7916 14720
rect 7852 14660 7856 14716
rect 7856 14660 7912 14716
rect 7912 14660 7916 14716
rect 7852 14656 7916 14660
rect 7932 14716 7996 14720
rect 7932 14660 7936 14716
rect 7936 14660 7992 14716
rect 7992 14660 7996 14716
rect 7932 14656 7996 14660
rect 8012 14716 8076 14720
rect 8012 14660 8016 14716
rect 8016 14660 8072 14716
rect 8072 14660 8076 14716
rect 8012 14656 8076 14660
rect 8092 14716 8156 14720
rect 8092 14660 8096 14716
rect 8096 14660 8152 14716
rect 8152 14660 8156 14716
rect 8092 14656 8156 14660
rect 14752 14716 14816 14720
rect 14752 14660 14756 14716
rect 14756 14660 14812 14716
rect 14812 14660 14816 14716
rect 14752 14656 14816 14660
rect 14832 14716 14896 14720
rect 14832 14660 14836 14716
rect 14836 14660 14892 14716
rect 14892 14660 14896 14716
rect 14832 14656 14896 14660
rect 14912 14716 14976 14720
rect 14912 14660 14916 14716
rect 14916 14660 14972 14716
rect 14972 14660 14976 14716
rect 14912 14656 14976 14660
rect 14992 14716 15056 14720
rect 14992 14660 14996 14716
rect 14996 14660 15052 14716
rect 15052 14660 15056 14716
rect 14992 14656 15056 14660
rect 4402 14172 4466 14176
rect 4402 14116 4406 14172
rect 4406 14116 4462 14172
rect 4462 14116 4466 14172
rect 4402 14112 4466 14116
rect 4482 14172 4546 14176
rect 4482 14116 4486 14172
rect 4486 14116 4542 14172
rect 4542 14116 4546 14172
rect 4482 14112 4546 14116
rect 4562 14172 4626 14176
rect 4562 14116 4566 14172
rect 4566 14116 4622 14172
rect 4622 14116 4626 14172
rect 4562 14112 4626 14116
rect 4642 14172 4706 14176
rect 4642 14116 4646 14172
rect 4646 14116 4702 14172
rect 4702 14116 4706 14172
rect 4642 14112 4706 14116
rect 11302 14172 11366 14176
rect 11302 14116 11306 14172
rect 11306 14116 11362 14172
rect 11362 14116 11366 14172
rect 11302 14112 11366 14116
rect 11382 14172 11446 14176
rect 11382 14116 11386 14172
rect 11386 14116 11442 14172
rect 11442 14116 11446 14172
rect 11382 14112 11446 14116
rect 11462 14172 11526 14176
rect 11462 14116 11466 14172
rect 11466 14116 11522 14172
rect 11522 14116 11526 14172
rect 11462 14112 11526 14116
rect 11542 14172 11606 14176
rect 11542 14116 11546 14172
rect 11546 14116 11602 14172
rect 11602 14116 11606 14172
rect 11542 14112 11606 14116
rect 18202 14172 18266 14176
rect 18202 14116 18206 14172
rect 18206 14116 18262 14172
rect 18262 14116 18266 14172
rect 18202 14112 18266 14116
rect 18282 14172 18346 14176
rect 18282 14116 18286 14172
rect 18286 14116 18342 14172
rect 18342 14116 18346 14172
rect 18282 14112 18346 14116
rect 18362 14172 18426 14176
rect 18362 14116 18366 14172
rect 18366 14116 18422 14172
rect 18422 14116 18426 14172
rect 18362 14112 18426 14116
rect 18442 14172 18506 14176
rect 18442 14116 18446 14172
rect 18446 14116 18502 14172
rect 18502 14116 18506 14172
rect 18442 14112 18506 14116
rect 7852 13628 7916 13632
rect 7852 13572 7856 13628
rect 7856 13572 7912 13628
rect 7912 13572 7916 13628
rect 7852 13568 7916 13572
rect 7932 13628 7996 13632
rect 7932 13572 7936 13628
rect 7936 13572 7992 13628
rect 7992 13572 7996 13628
rect 7932 13568 7996 13572
rect 8012 13628 8076 13632
rect 8012 13572 8016 13628
rect 8016 13572 8072 13628
rect 8072 13572 8076 13628
rect 8012 13568 8076 13572
rect 8092 13628 8156 13632
rect 8092 13572 8096 13628
rect 8096 13572 8152 13628
rect 8152 13572 8156 13628
rect 8092 13568 8156 13572
rect 14752 13628 14816 13632
rect 14752 13572 14756 13628
rect 14756 13572 14812 13628
rect 14812 13572 14816 13628
rect 14752 13568 14816 13572
rect 14832 13628 14896 13632
rect 14832 13572 14836 13628
rect 14836 13572 14892 13628
rect 14892 13572 14896 13628
rect 14832 13568 14896 13572
rect 14912 13628 14976 13632
rect 14912 13572 14916 13628
rect 14916 13572 14972 13628
rect 14972 13572 14976 13628
rect 14912 13568 14976 13572
rect 14992 13628 15056 13632
rect 14992 13572 14996 13628
rect 14996 13572 15052 13628
rect 15052 13572 15056 13628
rect 14992 13568 15056 13572
rect 4402 13084 4466 13088
rect 4402 13028 4406 13084
rect 4406 13028 4462 13084
rect 4462 13028 4466 13084
rect 4402 13024 4466 13028
rect 4482 13084 4546 13088
rect 4482 13028 4486 13084
rect 4486 13028 4542 13084
rect 4542 13028 4546 13084
rect 4482 13024 4546 13028
rect 4562 13084 4626 13088
rect 4562 13028 4566 13084
rect 4566 13028 4622 13084
rect 4622 13028 4626 13084
rect 4562 13024 4626 13028
rect 4642 13084 4706 13088
rect 4642 13028 4646 13084
rect 4646 13028 4702 13084
rect 4702 13028 4706 13084
rect 4642 13024 4706 13028
rect 11302 13084 11366 13088
rect 11302 13028 11306 13084
rect 11306 13028 11362 13084
rect 11362 13028 11366 13084
rect 11302 13024 11366 13028
rect 11382 13084 11446 13088
rect 11382 13028 11386 13084
rect 11386 13028 11442 13084
rect 11442 13028 11446 13084
rect 11382 13024 11446 13028
rect 11462 13084 11526 13088
rect 11462 13028 11466 13084
rect 11466 13028 11522 13084
rect 11522 13028 11526 13084
rect 11462 13024 11526 13028
rect 11542 13084 11606 13088
rect 11542 13028 11546 13084
rect 11546 13028 11602 13084
rect 11602 13028 11606 13084
rect 11542 13024 11606 13028
rect 18202 13084 18266 13088
rect 18202 13028 18206 13084
rect 18206 13028 18262 13084
rect 18262 13028 18266 13084
rect 18202 13024 18266 13028
rect 18282 13084 18346 13088
rect 18282 13028 18286 13084
rect 18286 13028 18342 13084
rect 18342 13028 18346 13084
rect 18282 13024 18346 13028
rect 18362 13084 18426 13088
rect 18362 13028 18366 13084
rect 18366 13028 18422 13084
rect 18422 13028 18426 13084
rect 18362 13024 18426 13028
rect 18442 13084 18506 13088
rect 18442 13028 18446 13084
rect 18446 13028 18502 13084
rect 18502 13028 18506 13084
rect 18442 13024 18506 13028
rect 7852 12540 7916 12544
rect 7852 12484 7856 12540
rect 7856 12484 7912 12540
rect 7912 12484 7916 12540
rect 7852 12480 7916 12484
rect 7932 12540 7996 12544
rect 7932 12484 7936 12540
rect 7936 12484 7992 12540
rect 7992 12484 7996 12540
rect 7932 12480 7996 12484
rect 8012 12540 8076 12544
rect 8012 12484 8016 12540
rect 8016 12484 8072 12540
rect 8072 12484 8076 12540
rect 8012 12480 8076 12484
rect 8092 12540 8156 12544
rect 8092 12484 8096 12540
rect 8096 12484 8152 12540
rect 8152 12484 8156 12540
rect 8092 12480 8156 12484
rect 14752 12540 14816 12544
rect 14752 12484 14756 12540
rect 14756 12484 14812 12540
rect 14812 12484 14816 12540
rect 14752 12480 14816 12484
rect 14832 12540 14896 12544
rect 14832 12484 14836 12540
rect 14836 12484 14892 12540
rect 14892 12484 14896 12540
rect 14832 12480 14896 12484
rect 14912 12540 14976 12544
rect 14912 12484 14916 12540
rect 14916 12484 14972 12540
rect 14972 12484 14976 12540
rect 14912 12480 14976 12484
rect 14992 12540 15056 12544
rect 14992 12484 14996 12540
rect 14996 12484 15052 12540
rect 15052 12484 15056 12540
rect 14992 12480 15056 12484
rect 4402 11996 4466 12000
rect 4402 11940 4406 11996
rect 4406 11940 4462 11996
rect 4462 11940 4466 11996
rect 4402 11936 4466 11940
rect 4482 11996 4546 12000
rect 4482 11940 4486 11996
rect 4486 11940 4542 11996
rect 4542 11940 4546 11996
rect 4482 11936 4546 11940
rect 4562 11996 4626 12000
rect 4562 11940 4566 11996
rect 4566 11940 4622 11996
rect 4622 11940 4626 11996
rect 4562 11936 4626 11940
rect 4642 11996 4706 12000
rect 4642 11940 4646 11996
rect 4646 11940 4702 11996
rect 4702 11940 4706 11996
rect 4642 11936 4706 11940
rect 11302 11996 11366 12000
rect 11302 11940 11306 11996
rect 11306 11940 11362 11996
rect 11362 11940 11366 11996
rect 11302 11936 11366 11940
rect 11382 11996 11446 12000
rect 11382 11940 11386 11996
rect 11386 11940 11442 11996
rect 11442 11940 11446 11996
rect 11382 11936 11446 11940
rect 11462 11996 11526 12000
rect 11462 11940 11466 11996
rect 11466 11940 11522 11996
rect 11522 11940 11526 11996
rect 11462 11936 11526 11940
rect 11542 11996 11606 12000
rect 11542 11940 11546 11996
rect 11546 11940 11602 11996
rect 11602 11940 11606 11996
rect 11542 11936 11606 11940
rect 18202 11996 18266 12000
rect 18202 11940 18206 11996
rect 18206 11940 18262 11996
rect 18262 11940 18266 11996
rect 18202 11936 18266 11940
rect 18282 11996 18346 12000
rect 18282 11940 18286 11996
rect 18286 11940 18342 11996
rect 18342 11940 18346 11996
rect 18282 11936 18346 11940
rect 18362 11996 18426 12000
rect 18362 11940 18366 11996
rect 18366 11940 18422 11996
rect 18422 11940 18426 11996
rect 18362 11936 18426 11940
rect 18442 11996 18506 12000
rect 18442 11940 18446 11996
rect 18446 11940 18502 11996
rect 18502 11940 18506 11996
rect 18442 11936 18506 11940
rect 7852 11452 7916 11456
rect 7852 11396 7856 11452
rect 7856 11396 7912 11452
rect 7912 11396 7916 11452
rect 7852 11392 7916 11396
rect 7932 11452 7996 11456
rect 7932 11396 7936 11452
rect 7936 11396 7992 11452
rect 7992 11396 7996 11452
rect 7932 11392 7996 11396
rect 8012 11452 8076 11456
rect 8012 11396 8016 11452
rect 8016 11396 8072 11452
rect 8072 11396 8076 11452
rect 8012 11392 8076 11396
rect 8092 11452 8156 11456
rect 8092 11396 8096 11452
rect 8096 11396 8152 11452
rect 8152 11396 8156 11452
rect 8092 11392 8156 11396
rect 14752 11452 14816 11456
rect 14752 11396 14756 11452
rect 14756 11396 14812 11452
rect 14812 11396 14816 11452
rect 14752 11392 14816 11396
rect 14832 11452 14896 11456
rect 14832 11396 14836 11452
rect 14836 11396 14892 11452
rect 14892 11396 14896 11452
rect 14832 11392 14896 11396
rect 14912 11452 14976 11456
rect 14912 11396 14916 11452
rect 14916 11396 14972 11452
rect 14972 11396 14976 11452
rect 14912 11392 14976 11396
rect 14992 11452 15056 11456
rect 14992 11396 14996 11452
rect 14996 11396 15052 11452
rect 15052 11396 15056 11452
rect 14992 11392 15056 11396
rect 4402 10908 4466 10912
rect 4402 10852 4406 10908
rect 4406 10852 4462 10908
rect 4462 10852 4466 10908
rect 4402 10848 4466 10852
rect 4482 10908 4546 10912
rect 4482 10852 4486 10908
rect 4486 10852 4542 10908
rect 4542 10852 4546 10908
rect 4482 10848 4546 10852
rect 4562 10908 4626 10912
rect 4562 10852 4566 10908
rect 4566 10852 4622 10908
rect 4622 10852 4626 10908
rect 4562 10848 4626 10852
rect 4642 10908 4706 10912
rect 4642 10852 4646 10908
rect 4646 10852 4702 10908
rect 4702 10852 4706 10908
rect 4642 10848 4706 10852
rect 11302 10908 11366 10912
rect 11302 10852 11306 10908
rect 11306 10852 11362 10908
rect 11362 10852 11366 10908
rect 11302 10848 11366 10852
rect 11382 10908 11446 10912
rect 11382 10852 11386 10908
rect 11386 10852 11442 10908
rect 11442 10852 11446 10908
rect 11382 10848 11446 10852
rect 11462 10908 11526 10912
rect 11462 10852 11466 10908
rect 11466 10852 11522 10908
rect 11522 10852 11526 10908
rect 11462 10848 11526 10852
rect 11542 10908 11606 10912
rect 11542 10852 11546 10908
rect 11546 10852 11602 10908
rect 11602 10852 11606 10908
rect 11542 10848 11606 10852
rect 18202 10908 18266 10912
rect 18202 10852 18206 10908
rect 18206 10852 18262 10908
rect 18262 10852 18266 10908
rect 18202 10848 18266 10852
rect 18282 10908 18346 10912
rect 18282 10852 18286 10908
rect 18286 10852 18342 10908
rect 18342 10852 18346 10908
rect 18282 10848 18346 10852
rect 18362 10908 18426 10912
rect 18362 10852 18366 10908
rect 18366 10852 18422 10908
rect 18422 10852 18426 10908
rect 18362 10848 18426 10852
rect 18442 10908 18506 10912
rect 18442 10852 18446 10908
rect 18446 10852 18502 10908
rect 18502 10852 18506 10908
rect 18442 10848 18506 10852
rect 7852 10364 7916 10368
rect 7852 10308 7856 10364
rect 7856 10308 7912 10364
rect 7912 10308 7916 10364
rect 7852 10304 7916 10308
rect 7932 10364 7996 10368
rect 7932 10308 7936 10364
rect 7936 10308 7992 10364
rect 7992 10308 7996 10364
rect 7932 10304 7996 10308
rect 8012 10364 8076 10368
rect 8012 10308 8016 10364
rect 8016 10308 8072 10364
rect 8072 10308 8076 10364
rect 8012 10304 8076 10308
rect 8092 10364 8156 10368
rect 8092 10308 8096 10364
rect 8096 10308 8152 10364
rect 8152 10308 8156 10364
rect 8092 10304 8156 10308
rect 14752 10364 14816 10368
rect 14752 10308 14756 10364
rect 14756 10308 14812 10364
rect 14812 10308 14816 10364
rect 14752 10304 14816 10308
rect 14832 10364 14896 10368
rect 14832 10308 14836 10364
rect 14836 10308 14892 10364
rect 14892 10308 14896 10364
rect 14832 10304 14896 10308
rect 14912 10364 14976 10368
rect 14912 10308 14916 10364
rect 14916 10308 14972 10364
rect 14972 10308 14976 10364
rect 14912 10304 14976 10308
rect 14992 10364 15056 10368
rect 14992 10308 14996 10364
rect 14996 10308 15052 10364
rect 15052 10308 15056 10364
rect 14992 10304 15056 10308
rect 4402 9820 4466 9824
rect 4402 9764 4406 9820
rect 4406 9764 4462 9820
rect 4462 9764 4466 9820
rect 4402 9760 4466 9764
rect 4482 9820 4546 9824
rect 4482 9764 4486 9820
rect 4486 9764 4542 9820
rect 4542 9764 4546 9820
rect 4482 9760 4546 9764
rect 4562 9820 4626 9824
rect 4562 9764 4566 9820
rect 4566 9764 4622 9820
rect 4622 9764 4626 9820
rect 4562 9760 4626 9764
rect 4642 9820 4706 9824
rect 4642 9764 4646 9820
rect 4646 9764 4702 9820
rect 4702 9764 4706 9820
rect 4642 9760 4706 9764
rect 11302 9820 11366 9824
rect 11302 9764 11306 9820
rect 11306 9764 11362 9820
rect 11362 9764 11366 9820
rect 11302 9760 11366 9764
rect 11382 9820 11446 9824
rect 11382 9764 11386 9820
rect 11386 9764 11442 9820
rect 11442 9764 11446 9820
rect 11382 9760 11446 9764
rect 11462 9820 11526 9824
rect 11462 9764 11466 9820
rect 11466 9764 11522 9820
rect 11522 9764 11526 9820
rect 11462 9760 11526 9764
rect 11542 9820 11606 9824
rect 11542 9764 11546 9820
rect 11546 9764 11602 9820
rect 11602 9764 11606 9820
rect 11542 9760 11606 9764
rect 18202 9820 18266 9824
rect 18202 9764 18206 9820
rect 18206 9764 18262 9820
rect 18262 9764 18266 9820
rect 18202 9760 18266 9764
rect 18282 9820 18346 9824
rect 18282 9764 18286 9820
rect 18286 9764 18342 9820
rect 18342 9764 18346 9820
rect 18282 9760 18346 9764
rect 18362 9820 18426 9824
rect 18362 9764 18366 9820
rect 18366 9764 18422 9820
rect 18422 9764 18426 9820
rect 18362 9760 18426 9764
rect 18442 9820 18506 9824
rect 18442 9764 18446 9820
rect 18446 9764 18502 9820
rect 18502 9764 18506 9820
rect 18442 9760 18506 9764
rect 7852 9276 7916 9280
rect 7852 9220 7856 9276
rect 7856 9220 7912 9276
rect 7912 9220 7916 9276
rect 7852 9216 7916 9220
rect 7932 9276 7996 9280
rect 7932 9220 7936 9276
rect 7936 9220 7992 9276
rect 7992 9220 7996 9276
rect 7932 9216 7996 9220
rect 8012 9276 8076 9280
rect 8012 9220 8016 9276
rect 8016 9220 8072 9276
rect 8072 9220 8076 9276
rect 8012 9216 8076 9220
rect 8092 9276 8156 9280
rect 8092 9220 8096 9276
rect 8096 9220 8152 9276
rect 8152 9220 8156 9276
rect 8092 9216 8156 9220
rect 14752 9276 14816 9280
rect 14752 9220 14756 9276
rect 14756 9220 14812 9276
rect 14812 9220 14816 9276
rect 14752 9216 14816 9220
rect 14832 9276 14896 9280
rect 14832 9220 14836 9276
rect 14836 9220 14892 9276
rect 14892 9220 14896 9276
rect 14832 9216 14896 9220
rect 14912 9276 14976 9280
rect 14912 9220 14916 9276
rect 14916 9220 14972 9276
rect 14972 9220 14976 9276
rect 14912 9216 14976 9220
rect 14992 9276 15056 9280
rect 14992 9220 14996 9276
rect 14996 9220 15052 9276
rect 15052 9220 15056 9276
rect 14992 9216 15056 9220
rect 4402 8732 4466 8736
rect 4402 8676 4406 8732
rect 4406 8676 4462 8732
rect 4462 8676 4466 8732
rect 4402 8672 4466 8676
rect 4482 8732 4546 8736
rect 4482 8676 4486 8732
rect 4486 8676 4542 8732
rect 4542 8676 4546 8732
rect 4482 8672 4546 8676
rect 4562 8732 4626 8736
rect 4562 8676 4566 8732
rect 4566 8676 4622 8732
rect 4622 8676 4626 8732
rect 4562 8672 4626 8676
rect 4642 8732 4706 8736
rect 4642 8676 4646 8732
rect 4646 8676 4702 8732
rect 4702 8676 4706 8732
rect 4642 8672 4706 8676
rect 11302 8732 11366 8736
rect 11302 8676 11306 8732
rect 11306 8676 11362 8732
rect 11362 8676 11366 8732
rect 11302 8672 11366 8676
rect 11382 8732 11446 8736
rect 11382 8676 11386 8732
rect 11386 8676 11442 8732
rect 11442 8676 11446 8732
rect 11382 8672 11446 8676
rect 11462 8732 11526 8736
rect 11462 8676 11466 8732
rect 11466 8676 11522 8732
rect 11522 8676 11526 8732
rect 11462 8672 11526 8676
rect 11542 8732 11606 8736
rect 11542 8676 11546 8732
rect 11546 8676 11602 8732
rect 11602 8676 11606 8732
rect 11542 8672 11606 8676
rect 18202 8732 18266 8736
rect 18202 8676 18206 8732
rect 18206 8676 18262 8732
rect 18262 8676 18266 8732
rect 18202 8672 18266 8676
rect 18282 8732 18346 8736
rect 18282 8676 18286 8732
rect 18286 8676 18342 8732
rect 18342 8676 18346 8732
rect 18282 8672 18346 8676
rect 18362 8732 18426 8736
rect 18362 8676 18366 8732
rect 18366 8676 18422 8732
rect 18422 8676 18426 8732
rect 18362 8672 18426 8676
rect 18442 8732 18506 8736
rect 18442 8676 18446 8732
rect 18446 8676 18502 8732
rect 18502 8676 18506 8732
rect 18442 8672 18506 8676
rect 7852 8188 7916 8192
rect 7852 8132 7856 8188
rect 7856 8132 7912 8188
rect 7912 8132 7916 8188
rect 7852 8128 7916 8132
rect 7932 8188 7996 8192
rect 7932 8132 7936 8188
rect 7936 8132 7992 8188
rect 7992 8132 7996 8188
rect 7932 8128 7996 8132
rect 8012 8188 8076 8192
rect 8012 8132 8016 8188
rect 8016 8132 8072 8188
rect 8072 8132 8076 8188
rect 8012 8128 8076 8132
rect 8092 8188 8156 8192
rect 8092 8132 8096 8188
rect 8096 8132 8152 8188
rect 8152 8132 8156 8188
rect 8092 8128 8156 8132
rect 14752 8188 14816 8192
rect 14752 8132 14756 8188
rect 14756 8132 14812 8188
rect 14812 8132 14816 8188
rect 14752 8128 14816 8132
rect 14832 8188 14896 8192
rect 14832 8132 14836 8188
rect 14836 8132 14892 8188
rect 14892 8132 14896 8188
rect 14832 8128 14896 8132
rect 14912 8188 14976 8192
rect 14912 8132 14916 8188
rect 14916 8132 14972 8188
rect 14972 8132 14976 8188
rect 14912 8128 14976 8132
rect 14992 8188 15056 8192
rect 14992 8132 14996 8188
rect 14996 8132 15052 8188
rect 15052 8132 15056 8188
rect 14992 8128 15056 8132
rect 4402 7644 4466 7648
rect 4402 7588 4406 7644
rect 4406 7588 4462 7644
rect 4462 7588 4466 7644
rect 4402 7584 4466 7588
rect 4482 7644 4546 7648
rect 4482 7588 4486 7644
rect 4486 7588 4542 7644
rect 4542 7588 4546 7644
rect 4482 7584 4546 7588
rect 4562 7644 4626 7648
rect 4562 7588 4566 7644
rect 4566 7588 4622 7644
rect 4622 7588 4626 7644
rect 4562 7584 4626 7588
rect 4642 7644 4706 7648
rect 4642 7588 4646 7644
rect 4646 7588 4702 7644
rect 4702 7588 4706 7644
rect 4642 7584 4706 7588
rect 11302 7644 11366 7648
rect 11302 7588 11306 7644
rect 11306 7588 11362 7644
rect 11362 7588 11366 7644
rect 11302 7584 11366 7588
rect 11382 7644 11446 7648
rect 11382 7588 11386 7644
rect 11386 7588 11442 7644
rect 11442 7588 11446 7644
rect 11382 7584 11446 7588
rect 11462 7644 11526 7648
rect 11462 7588 11466 7644
rect 11466 7588 11522 7644
rect 11522 7588 11526 7644
rect 11462 7584 11526 7588
rect 11542 7644 11606 7648
rect 11542 7588 11546 7644
rect 11546 7588 11602 7644
rect 11602 7588 11606 7644
rect 11542 7584 11606 7588
rect 18202 7644 18266 7648
rect 18202 7588 18206 7644
rect 18206 7588 18262 7644
rect 18262 7588 18266 7644
rect 18202 7584 18266 7588
rect 18282 7644 18346 7648
rect 18282 7588 18286 7644
rect 18286 7588 18342 7644
rect 18342 7588 18346 7644
rect 18282 7584 18346 7588
rect 18362 7644 18426 7648
rect 18362 7588 18366 7644
rect 18366 7588 18422 7644
rect 18422 7588 18426 7644
rect 18362 7584 18426 7588
rect 18442 7644 18506 7648
rect 18442 7588 18446 7644
rect 18446 7588 18502 7644
rect 18502 7588 18506 7644
rect 18442 7584 18506 7588
rect 7852 7100 7916 7104
rect 7852 7044 7856 7100
rect 7856 7044 7912 7100
rect 7912 7044 7916 7100
rect 7852 7040 7916 7044
rect 7932 7100 7996 7104
rect 7932 7044 7936 7100
rect 7936 7044 7992 7100
rect 7992 7044 7996 7100
rect 7932 7040 7996 7044
rect 8012 7100 8076 7104
rect 8012 7044 8016 7100
rect 8016 7044 8072 7100
rect 8072 7044 8076 7100
rect 8012 7040 8076 7044
rect 8092 7100 8156 7104
rect 8092 7044 8096 7100
rect 8096 7044 8152 7100
rect 8152 7044 8156 7100
rect 8092 7040 8156 7044
rect 14752 7100 14816 7104
rect 14752 7044 14756 7100
rect 14756 7044 14812 7100
rect 14812 7044 14816 7100
rect 14752 7040 14816 7044
rect 14832 7100 14896 7104
rect 14832 7044 14836 7100
rect 14836 7044 14892 7100
rect 14892 7044 14896 7100
rect 14832 7040 14896 7044
rect 14912 7100 14976 7104
rect 14912 7044 14916 7100
rect 14916 7044 14972 7100
rect 14972 7044 14976 7100
rect 14912 7040 14976 7044
rect 14992 7100 15056 7104
rect 14992 7044 14996 7100
rect 14996 7044 15052 7100
rect 15052 7044 15056 7100
rect 14992 7040 15056 7044
rect 4402 6556 4466 6560
rect 4402 6500 4406 6556
rect 4406 6500 4462 6556
rect 4462 6500 4466 6556
rect 4402 6496 4466 6500
rect 4482 6556 4546 6560
rect 4482 6500 4486 6556
rect 4486 6500 4542 6556
rect 4542 6500 4546 6556
rect 4482 6496 4546 6500
rect 4562 6556 4626 6560
rect 4562 6500 4566 6556
rect 4566 6500 4622 6556
rect 4622 6500 4626 6556
rect 4562 6496 4626 6500
rect 4642 6556 4706 6560
rect 4642 6500 4646 6556
rect 4646 6500 4702 6556
rect 4702 6500 4706 6556
rect 4642 6496 4706 6500
rect 11302 6556 11366 6560
rect 11302 6500 11306 6556
rect 11306 6500 11362 6556
rect 11362 6500 11366 6556
rect 11302 6496 11366 6500
rect 11382 6556 11446 6560
rect 11382 6500 11386 6556
rect 11386 6500 11442 6556
rect 11442 6500 11446 6556
rect 11382 6496 11446 6500
rect 11462 6556 11526 6560
rect 11462 6500 11466 6556
rect 11466 6500 11522 6556
rect 11522 6500 11526 6556
rect 11462 6496 11526 6500
rect 11542 6556 11606 6560
rect 11542 6500 11546 6556
rect 11546 6500 11602 6556
rect 11602 6500 11606 6556
rect 11542 6496 11606 6500
rect 18202 6556 18266 6560
rect 18202 6500 18206 6556
rect 18206 6500 18262 6556
rect 18262 6500 18266 6556
rect 18202 6496 18266 6500
rect 18282 6556 18346 6560
rect 18282 6500 18286 6556
rect 18286 6500 18342 6556
rect 18342 6500 18346 6556
rect 18282 6496 18346 6500
rect 18362 6556 18426 6560
rect 18362 6500 18366 6556
rect 18366 6500 18422 6556
rect 18422 6500 18426 6556
rect 18362 6496 18426 6500
rect 18442 6556 18506 6560
rect 18442 6500 18446 6556
rect 18446 6500 18502 6556
rect 18502 6500 18506 6556
rect 18442 6496 18506 6500
rect 7852 6012 7916 6016
rect 7852 5956 7856 6012
rect 7856 5956 7912 6012
rect 7912 5956 7916 6012
rect 7852 5952 7916 5956
rect 7932 6012 7996 6016
rect 7932 5956 7936 6012
rect 7936 5956 7992 6012
rect 7992 5956 7996 6012
rect 7932 5952 7996 5956
rect 8012 6012 8076 6016
rect 8012 5956 8016 6012
rect 8016 5956 8072 6012
rect 8072 5956 8076 6012
rect 8012 5952 8076 5956
rect 8092 6012 8156 6016
rect 8092 5956 8096 6012
rect 8096 5956 8152 6012
rect 8152 5956 8156 6012
rect 8092 5952 8156 5956
rect 14752 6012 14816 6016
rect 14752 5956 14756 6012
rect 14756 5956 14812 6012
rect 14812 5956 14816 6012
rect 14752 5952 14816 5956
rect 14832 6012 14896 6016
rect 14832 5956 14836 6012
rect 14836 5956 14892 6012
rect 14892 5956 14896 6012
rect 14832 5952 14896 5956
rect 14912 6012 14976 6016
rect 14912 5956 14916 6012
rect 14916 5956 14972 6012
rect 14972 5956 14976 6012
rect 14912 5952 14976 5956
rect 14992 6012 15056 6016
rect 14992 5956 14996 6012
rect 14996 5956 15052 6012
rect 15052 5956 15056 6012
rect 14992 5952 15056 5956
rect 4402 5468 4466 5472
rect 4402 5412 4406 5468
rect 4406 5412 4462 5468
rect 4462 5412 4466 5468
rect 4402 5408 4466 5412
rect 4482 5468 4546 5472
rect 4482 5412 4486 5468
rect 4486 5412 4542 5468
rect 4542 5412 4546 5468
rect 4482 5408 4546 5412
rect 4562 5468 4626 5472
rect 4562 5412 4566 5468
rect 4566 5412 4622 5468
rect 4622 5412 4626 5468
rect 4562 5408 4626 5412
rect 4642 5468 4706 5472
rect 4642 5412 4646 5468
rect 4646 5412 4702 5468
rect 4702 5412 4706 5468
rect 4642 5408 4706 5412
rect 11302 5468 11366 5472
rect 11302 5412 11306 5468
rect 11306 5412 11362 5468
rect 11362 5412 11366 5468
rect 11302 5408 11366 5412
rect 11382 5468 11446 5472
rect 11382 5412 11386 5468
rect 11386 5412 11442 5468
rect 11442 5412 11446 5468
rect 11382 5408 11446 5412
rect 11462 5468 11526 5472
rect 11462 5412 11466 5468
rect 11466 5412 11522 5468
rect 11522 5412 11526 5468
rect 11462 5408 11526 5412
rect 11542 5468 11606 5472
rect 11542 5412 11546 5468
rect 11546 5412 11602 5468
rect 11602 5412 11606 5468
rect 11542 5408 11606 5412
rect 18202 5468 18266 5472
rect 18202 5412 18206 5468
rect 18206 5412 18262 5468
rect 18262 5412 18266 5468
rect 18202 5408 18266 5412
rect 18282 5468 18346 5472
rect 18282 5412 18286 5468
rect 18286 5412 18342 5468
rect 18342 5412 18346 5468
rect 18282 5408 18346 5412
rect 18362 5468 18426 5472
rect 18362 5412 18366 5468
rect 18366 5412 18422 5468
rect 18422 5412 18426 5468
rect 18362 5408 18426 5412
rect 18442 5468 18506 5472
rect 18442 5412 18446 5468
rect 18446 5412 18502 5468
rect 18502 5412 18506 5468
rect 18442 5408 18506 5412
rect 7852 4924 7916 4928
rect 7852 4868 7856 4924
rect 7856 4868 7912 4924
rect 7912 4868 7916 4924
rect 7852 4864 7916 4868
rect 7932 4924 7996 4928
rect 7932 4868 7936 4924
rect 7936 4868 7992 4924
rect 7992 4868 7996 4924
rect 7932 4864 7996 4868
rect 8012 4924 8076 4928
rect 8012 4868 8016 4924
rect 8016 4868 8072 4924
rect 8072 4868 8076 4924
rect 8012 4864 8076 4868
rect 8092 4924 8156 4928
rect 8092 4868 8096 4924
rect 8096 4868 8152 4924
rect 8152 4868 8156 4924
rect 8092 4864 8156 4868
rect 14752 4924 14816 4928
rect 14752 4868 14756 4924
rect 14756 4868 14812 4924
rect 14812 4868 14816 4924
rect 14752 4864 14816 4868
rect 14832 4924 14896 4928
rect 14832 4868 14836 4924
rect 14836 4868 14892 4924
rect 14892 4868 14896 4924
rect 14832 4864 14896 4868
rect 14912 4924 14976 4928
rect 14912 4868 14916 4924
rect 14916 4868 14972 4924
rect 14972 4868 14976 4924
rect 14912 4864 14976 4868
rect 14992 4924 15056 4928
rect 14992 4868 14996 4924
rect 14996 4868 15052 4924
rect 15052 4868 15056 4924
rect 14992 4864 15056 4868
rect 4402 4380 4466 4384
rect 4402 4324 4406 4380
rect 4406 4324 4462 4380
rect 4462 4324 4466 4380
rect 4402 4320 4466 4324
rect 4482 4380 4546 4384
rect 4482 4324 4486 4380
rect 4486 4324 4542 4380
rect 4542 4324 4546 4380
rect 4482 4320 4546 4324
rect 4562 4380 4626 4384
rect 4562 4324 4566 4380
rect 4566 4324 4622 4380
rect 4622 4324 4626 4380
rect 4562 4320 4626 4324
rect 4642 4380 4706 4384
rect 4642 4324 4646 4380
rect 4646 4324 4702 4380
rect 4702 4324 4706 4380
rect 4642 4320 4706 4324
rect 11302 4380 11366 4384
rect 11302 4324 11306 4380
rect 11306 4324 11362 4380
rect 11362 4324 11366 4380
rect 11302 4320 11366 4324
rect 11382 4380 11446 4384
rect 11382 4324 11386 4380
rect 11386 4324 11442 4380
rect 11442 4324 11446 4380
rect 11382 4320 11446 4324
rect 11462 4380 11526 4384
rect 11462 4324 11466 4380
rect 11466 4324 11522 4380
rect 11522 4324 11526 4380
rect 11462 4320 11526 4324
rect 11542 4380 11606 4384
rect 11542 4324 11546 4380
rect 11546 4324 11602 4380
rect 11602 4324 11606 4380
rect 11542 4320 11606 4324
rect 18202 4380 18266 4384
rect 18202 4324 18206 4380
rect 18206 4324 18262 4380
rect 18262 4324 18266 4380
rect 18202 4320 18266 4324
rect 18282 4380 18346 4384
rect 18282 4324 18286 4380
rect 18286 4324 18342 4380
rect 18342 4324 18346 4380
rect 18282 4320 18346 4324
rect 18362 4380 18426 4384
rect 18362 4324 18366 4380
rect 18366 4324 18422 4380
rect 18422 4324 18426 4380
rect 18362 4320 18426 4324
rect 18442 4380 18506 4384
rect 18442 4324 18446 4380
rect 18446 4324 18502 4380
rect 18502 4324 18506 4380
rect 18442 4320 18506 4324
rect 7852 3836 7916 3840
rect 7852 3780 7856 3836
rect 7856 3780 7912 3836
rect 7912 3780 7916 3836
rect 7852 3776 7916 3780
rect 7932 3836 7996 3840
rect 7932 3780 7936 3836
rect 7936 3780 7992 3836
rect 7992 3780 7996 3836
rect 7932 3776 7996 3780
rect 8012 3836 8076 3840
rect 8012 3780 8016 3836
rect 8016 3780 8072 3836
rect 8072 3780 8076 3836
rect 8012 3776 8076 3780
rect 8092 3836 8156 3840
rect 8092 3780 8096 3836
rect 8096 3780 8152 3836
rect 8152 3780 8156 3836
rect 8092 3776 8156 3780
rect 14752 3836 14816 3840
rect 14752 3780 14756 3836
rect 14756 3780 14812 3836
rect 14812 3780 14816 3836
rect 14752 3776 14816 3780
rect 14832 3836 14896 3840
rect 14832 3780 14836 3836
rect 14836 3780 14892 3836
rect 14892 3780 14896 3836
rect 14832 3776 14896 3780
rect 14912 3836 14976 3840
rect 14912 3780 14916 3836
rect 14916 3780 14972 3836
rect 14972 3780 14976 3836
rect 14912 3776 14976 3780
rect 14992 3836 15056 3840
rect 14992 3780 14996 3836
rect 14996 3780 15052 3836
rect 15052 3780 15056 3836
rect 14992 3776 15056 3780
rect 4402 3292 4466 3296
rect 4402 3236 4406 3292
rect 4406 3236 4462 3292
rect 4462 3236 4466 3292
rect 4402 3232 4466 3236
rect 4482 3292 4546 3296
rect 4482 3236 4486 3292
rect 4486 3236 4542 3292
rect 4542 3236 4546 3292
rect 4482 3232 4546 3236
rect 4562 3292 4626 3296
rect 4562 3236 4566 3292
rect 4566 3236 4622 3292
rect 4622 3236 4626 3292
rect 4562 3232 4626 3236
rect 4642 3292 4706 3296
rect 4642 3236 4646 3292
rect 4646 3236 4702 3292
rect 4702 3236 4706 3292
rect 4642 3232 4706 3236
rect 11302 3292 11366 3296
rect 11302 3236 11306 3292
rect 11306 3236 11362 3292
rect 11362 3236 11366 3292
rect 11302 3232 11366 3236
rect 11382 3292 11446 3296
rect 11382 3236 11386 3292
rect 11386 3236 11442 3292
rect 11442 3236 11446 3292
rect 11382 3232 11446 3236
rect 11462 3292 11526 3296
rect 11462 3236 11466 3292
rect 11466 3236 11522 3292
rect 11522 3236 11526 3292
rect 11462 3232 11526 3236
rect 11542 3292 11606 3296
rect 11542 3236 11546 3292
rect 11546 3236 11602 3292
rect 11602 3236 11606 3292
rect 11542 3232 11606 3236
rect 18202 3292 18266 3296
rect 18202 3236 18206 3292
rect 18206 3236 18262 3292
rect 18262 3236 18266 3292
rect 18202 3232 18266 3236
rect 18282 3292 18346 3296
rect 18282 3236 18286 3292
rect 18286 3236 18342 3292
rect 18342 3236 18346 3292
rect 18282 3232 18346 3236
rect 18362 3292 18426 3296
rect 18362 3236 18366 3292
rect 18366 3236 18422 3292
rect 18422 3236 18426 3292
rect 18362 3232 18426 3236
rect 18442 3292 18506 3296
rect 18442 3236 18446 3292
rect 18446 3236 18502 3292
rect 18502 3236 18506 3292
rect 18442 3232 18506 3236
rect 7852 2748 7916 2752
rect 7852 2692 7856 2748
rect 7856 2692 7912 2748
rect 7912 2692 7916 2748
rect 7852 2688 7916 2692
rect 7932 2748 7996 2752
rect 7932 2692 7936 2748
rect 7936 2692 7992 2748
rect 7992 2692 7996 2748
rect 7932 2688 7996 2692
rect 8012 2748 8076 2752
rect 8012 2692 8016 2748
rect 8016 2692 8072 2748
rect 8072 2692 8076 2748
rect 8012 2688 8076 2692
rect 8092 2748 8156 2752
rect 8092 2692 8096 2748
rect 8096 2692 8152 2748
rect 8152 2692 8156 2748
rect 8092 2688 8156 2692
rect 14752 2748 14816 2752
rect 14752 2692 14756 2748
rect 14756 2692 14812 2748
rect 14812 2692 14816 2748
rect 14752 2688 14816 2692
rect 14832 2748 14896 2752
rect 14832 2692 14836 2748
rect 14836 2692 14892 2748
rect 14892 2692 14896 2748
rect 14832 2688 14896 2692
rect 14912 2748 14976 2752
rect 14912 2692 14916 2748
rect 14916 2692 14972 2748
rect 14972 2692 14976 2748
rect 14912 2688 14976 2692
rect 14992 2748 15056 2752
rect 14992 2692 14996 2748
rect 14996 2692 15052 2748
rect 15052 2692 15056 2748
rect 14992 2688 15056 2692
rect 4402 2204 4466 2208
rect 4402 2148 4406 2204
rect 4406 2148 4462 2204
rect 4462 2148 4466 2204
rect 4402 2144 4466 2148
rect 4482 2204 4546 2208
rect 4482 2148 4486 2204
rect 4486 2148 4542 2204
rect 4542 2148 4546 2204
rect 4482 2144 4546 2148
rect 4562 2204 4626 2208
rect 4562 2148 4566 2204
rect 4566 2148 4622 2204
rect 4622 2148 4626 2204
rect 4562 2144 4626 2148
rect 4642 2204 4706 2208
rect 4642 2148 4646 2204
rect 4646 2148 4702 2204
rect 4702 2148 4706 2204
rect 4642 2144 4706 2148
rect 11302 2204 11366 2208
rect 11302 2148 11306 2204
rect 11306 2148 11362 2204
rect 11362 2148 11366 2204
rect 11302 2144 11366 2148
rect 11382 2204 11446 2208
rect 11382 2148 11386 2204
rect 11386 2148 11442 2204
rect 11442 2148 11446 2204
rect 11382 2144 11446 2148
rect 11462 2204 11526 2208
rect 11462 2148 11466 2204
rect 11466 2148 11522 2204
rect 11522 2148 11526 2204
rect 11462 2144 11526 2148
rect 11542 2204 11606 2208
rect 11542 2148 11546 2204
rect 11546 2148 11602 2204
rect 11602 2148 11606 2204
rect 11542 2144 11606 2148
rect 18202 2204 18266 2208
rect 18202 2148 18206 2204
rect 18206 2148 18262 2204
rect 18262 2148 18266 2204
rect 18202 2144 18266 2148
rect 18282 2204 18346 2208
rect 18282 2148 18286 2204
rect 18286 2148 18342 2204
rect 18342 2148 18346 2204
rect 18282 2144 18346 2148
rect 18362 2204 18426 2208
rect 18362 2148 18366 2204
rect 18366 2148 18422 2204
rect 18422 2148 18426 2204
rect 18362 2144 18426 2148
rect 18442 2204 18506 2208
rect 18442 2148 18446 2204
rect 18446 2148 18502 2204
rect 18502 2148 18506 2204
rect 18442 2144 18506 2148
<< metal4 >>
rect 4394 22880 4714 22896
rect 4394 22816 4402 22880
rect 4466 22816 4482 22880
rect 4546 22816 4562 22880
rect 4626 22816 4642 22880
rect 4706 22816 4714 22880
rect 4394 21792 4714 22816
rect 4394 21728 4402 21792
rect 4466 21728 4482 21792
rect 4546 21728 4562 21792
rect 4626 21728 4642 21792
rect 4706 21728 4714 21792
rect 4394 20704 4714 21728
rect 4394 20640 4402 20704
rect 4466 20640 4482 20704
rect 4546 20640 4562 20704
rect 4626 20640 4642 20704
rect 4706 20640 4714 20704
rect 4394 19616 4714 20640
rect 4394 19552 4402 19616
rect 4466 19552 4482 19616
rect 4546 19552 4562 19616
rect 4626 19552 4642 19616
rect 4706 19552 4714 19616
rect 4394 19472 4714 19552
rect 4394 19236 4436 19472
rect 4672 19236 4714 19472
rect 4394 18528 4714 19236
rect 4394 18464 4402 18528
rect 4466 18464 4482 18528
rect 4546 18464 4562 18528
rect 4626 18464 4642 18528
rect 4706 18464 4714 18528
rect 4394 17440 4714 18464
rect 4394 17376 4402 17440
rect 4466 17376 4482 17440
rect 4546 17376 4562 17440
rect 4626 17376 4642 17440
rect 4706 17376 4714 17440
rect 4394 16352 4714 17376
rect 4394 16288 4402 16352
rect 4466 16288 4482 16352
rect 4546 16288 4562 16352
rect 4626 16288 4642 16352
rect 4706 16288 4714 16352
rect 4394 15264 4714 16288
rect 4394 15200 4402 15264
rect 4466 15200 4482 15264
rect 4546 15200 4562 15264
rect 4626 15200 4642 15264
rect 4706 15200 4714 15264
rect 4394 14176 4714 15200
rect 4394 14112 4402 14176
rect 4466 14112 4482 14176
rect 4546 14112 4562 14176
rect 4626 14112 4642 14176
rect 4706 14112 4714 14176
rect 4394 13088 4714 14112
rect 4394 13024 4402 13088
rect 4466 13024 4482 13088
rect 4546 13024 4562 13088
rect 4626 13024 4642 13088
rect 4706 13024 4714 13088
rect 4394 12582 4714 13024
rect 4394 12346 4436 12582
rect 4672 12346 4714 12582
rect 4394 12000 4714 12346
rect 4394 11936 4402 12000
rect 4466 11936 4482 12000
rect 4546 11936 4562 12000
rect 4626 11936 4642 12000
rect 4706 11936 4714 12000
rect 4394 10912 4714 11936
rect 4394 10848 4402 10912
rect 4466 10848 4482 10912
rect 4546 10848 4562 10912
rect 4626 10848 4642 10912
rect 4706 10848 4714 10912
rect 4394 9824 4714 10848
rect 4394 9760 4402 9824
rect 4466 9760 4482 9824
rect 4546 9760 4562 9824
rect 4626 9760 4642 9824
rect 4706 9760 4714 9824
rect 4394 8736 4714 9760
rect 4394 8672 4402 8736
rect 4466 8672 4482 8736
rect 4546 8672 4562 8736
rect 4626 8672 4642 8736
rect 4706 8672 4714 8736
rect 4394 7648 4714 8672
rect 4394 7584 4402 7648
rect 4466 7584 4482 7648
rect 4546 7584 4562 7648
rect 4626 7584 4642 7648
rect 4706 7584 4714 7648
rect 4394 6560 4714 7584
rect 4394 6496 4402 6560
rect 4466 6496 4482 6560
rect 4546 6496 4562 6560
rect 4626 6496 4642 6560
rect 4706 6496 4714 6560
rect 4394 5691 4714 6496
rect 4394 5472 4436 5691
rect 4672 5472 4714 5691
rect 4394 5408 4402 5472
rect 4466 5408 4482 5455
rect 4546 5408 4562 5455
rect 4626 5408 4642 5455
rect 4706 5408 4714 5472
rect 4394 4384 4714 5408
rect 4394 4320 4402 4384
rect 4466 4320 4482 4384
rect 4546 4320 4562 4384
rect 4626 4320 4642 4384
rect 4706 4320 4714 4384
rect 4394 3296 4714 4320
rect 4394 3232 4402 3296
rect 4466 3232 4482 3296
rect 4546 3232 4562 3296
rect 4626 3232 4642 3296
rect 4706 3232 4714 3296
rect 4394 2208 4714 3232
rect 4394 2144 4402 2208
rect 4466 2144 4482 2208
rect 4546 2144 4562 2208
rect 4626 2144 4642 2208
rect 4706 2144 4714 2208
rect 4394 2128 4714 2144
rect 7844 22336 8164 22896
rect 7844 22272 7852 22336
rect 7916 22272 7932 22336
rect 7996 22272 8012 22336
rect 8076 22272 8092 22336
rect 8156 22272 8164 22336
rect 7844 21248 8164 22272
rect 7844 21184 7852 21248
rect 7916 21184 7932 21248
rect 7996 21184 8012 21248
rect 8076 21184 8092 21248
rect 8156 21184 8164 21248
rect 7844 20160 8164 21184
rect 7844 20096 7852 20160
rect 7916 20096 7932 20160
rect 7996 20096 8012 20160
rect 8076 20096 8092 20160
rect 8156 20096 8164 20160
rect 7844 19072 8164 20096
rect 7844 19008 7852 19072
rect 7916 19008 7932 19072
rect 7996 19008 8012 19072
rect 8076 19008 8092 19072
rect 8156 19008 8164 19072
rect 7844 17984 8164 19008
rect 7844 17920 7852 17984
rect 7916 17920 7932 17984
rect 7996 17920 8012 17984
rect 8076 17920 8092 17984
rect 8156 17920 8164 17984
rect 7844 16896 8164 17920
rect 7844 16832 7852 16896
rect 7916 16832 7932 16896
rect 7996 16832 8012 16896
rect 8076 16832 8092 16896
rect 8156 16832 8164 16896
rect 7844 16027 8164 16832
rect 7844 15808 7886 16027
rect 8122 15808 8164 16027
rect 7844 15744 7852 15808
rect 7916 15744 7932 15791
rect 7996 15744 8012 15791
rect 8076 15744 8092 15791
rect 8156 15744 8164 15808
rect 7844 14720 8164 15744
rect 7844 14656 7852 14720
rect 7916 14656 7932 14720
rect 7996 14656 8012 14720
rect 8076 14656 8092 14720
rect 8156 14656 8164 14720
rect 7844 13632 8164 14656
rect 7844 13568 7852 13632
rect 7916 13568 7932 13632
rect 7996 13568 8012 13632
rect 8076 13568 8092 13632
rect 8156 13568 8164 13632
rect 7844 12544 8164 13568
rect 7844 12480 7852 12544
rect 7916 12480 7932 12544
rect 7996 12480 8012 12544
rect 8076 12480 8092 12544
rect 8156 12480 8164 12544
rect 7844 11456 8164 12480
rect 7844 11392 7852 11456
rect 7916 11392 7932 11456
rect 7996 11392 8012 11456
rect 8076 11392 8092 11456
rect 8156 11392 8164 11456
rect 7844 10368 8164 11392
rect 7844 10304 7852 10368
rect 7916 10304 7932 10368
rect 7996 10304 8012 10368
rect 8076 10304 8092 10368
rect 8156 10304 8164 10368
rect 7844 9280 8164 10304
rect 7844 9216 7852 9280
rect 7916 9216 7932 9280
rect 7996 9216 8012 9280
rect 8076 9216 8092 9280
rect 8156 9216 8164 9280
rect 7844 9136 8164 9216
rect 7844 8900 7886 9136
rect 8122 8900 8164 9136
rect 7844 8192 8164 8900
rect 7844 8128 7852 8192
rect 7916 8128 7932 8192
rect 7996 8128 8012 8192
rect 8076 8128 8092 8192
rect 8156 8128 8164 8192
rect 7844 7104 8164 8128
rect 7844 7040 7852 7104
rect 7916 7040 7932 7104
rect 7996 7040 8012 7104
rect 8076 7040 8092 7104
rect 8156 7040 8164 7104
rect 7844 6016 8164 7040
rect 7844 5952 7852 6016
rect 7916 5952 7932 6016
rect 7996 5952 8012 6016
rect 8076 5952 8092 6016
rect 8156 5952 8164 6016
rect 7844 4928 8164 5952
rect 7844 4864 7852 4928
rect 7916 4864 7932 4928
rect 7996 4864 8012 4928
rect 8076 4864 8092 4928
rect 8156 4864 8164 4928
rect 7844 3840 8164 4864
rect 7844 3776 7852 3840
rect 7916 3776 7932 3840
rect 7996 3776 8012 3840
rect 8076 3776 8092 3840
rect 8156 3776 8164 3840
rect 7844 2752 8164 3776
rect 7844 2688 7852 2752
rect 7916 2688 7932 2752
rect 7996 2688 8012 2752
rect 8076 2688 8092 2752
rect 8156 2688 8164 2752
rect 7844 2128 8164 2688
rect 11294 22880 11614 22896
rect 11294 22816 11302 22880
rect 11366 22816 11382 22880
rect 11446 22816 11462 22880
rect 11526 22816 11542 22880
rect 11606 22816 11614 22880
rect 11294 21792 11614 22816
rect 11294 21728 11302 21792
rect 11366 21728 11382 21792
rect 11446 21728 11462 21792
rect 11526 21728 11542 21792
rect 11606 21728 11614 21792
rect 11294 20704 11614 21728
rect 11294 20640 11302 20704
rect 11366 20640 11382 20704
rect 11446 20640 11462 20704
rect 11526 20640 11542 20704
rect 11606 20640 11614 20704
rect 11294 19616 11614 20640
rect 11294 19552 11302 19616
rect 11366 19552 11382 19616
rect 11446 19552 11462 19616
rect 11526 19552 11542 19616
rect 11606 19552 11614 19616
rect 11294 19472 11614 19552
rect 11294 19236 11336 19472
rect 11572 19236 11614 19472
rect 11294 18528 11614 19236
rect 11294 18464 11302 18528
rect 11366 18464 11382 18528
rect 11446 18464 11462 18528
rect 11526 18464 11542 18528
rect 11606 18464 11614 18528
rect 11294 17440 11614 18464
rect 11294 17376 11302 17440
rect 11366 17376 11382 17440
rect 11446 17376 11462 17440
rect 11526 17376 11542 17440
rect 11606 17376 11614 17440
rect 11294 16352 11614 17376
rect 11294 16288 11302 16352
rect 11366 16288 11382 16352
rect 11446 16288 11462 16352
rect 11526 16288 11542 16352
rect 11606 16288 11614 16352
rect 11294 15264 11614 16288
rect 11294 15200 11302 15264
rect 11366 15200 11382 15264
rect 11446 15200 11462 15264
rect 11526 15200 11542 15264
rect 11606 15200 11614 15264
rect 11294 14176 11614 15200
rect 11294 14112 11302 14176
rect 11366 14112 11382 14176
rect 11446 14112 11462 14176
rect 11526 14112 11542 14176
rect 11606 14112 11614 14176
rect 11294 13088 11614 14112
rect 11294 13024 11302 13088
rect 11366 13024 11382 13088
rect 11446 13024 11462 13088
rect 11526 13024 11542 13088
rect 11606 13024 11614 13088
rect 11294 12582 11614 13024
rect 11294 12346 11336 12582
rect 11572 12346 11614 12582
rect 11294 12000 11614 12346
rect 11294 11936 11302 12000
rect 11366 11936 11382 12000
rect 11446 11936 11462 12000
rect 11526 11936 11542 12000
rect 11606 11936 11614 12000
rect 11294 10912 11614 11936
rect 11294 10848 11302 10912
rect 11366 10848 11382 10912
rect 11446 10848 11462 10912
rect 11526 10848 11542 10912
rect 11606 10848 11614 10912
rect 11294 9824 11614 10848
rect 11294 9760 11302 9824
rect 11366 9760 11382 9824
rect 11446 9760 11462 9824
rect 11526 9760 11542 9824
rect 11606 9760 11614 9824
rect 11294 8736 11614 9760
rect 11294 8672 11302 8736
rect 11366 8672 11382 8736
rect 11446 8672 11462 8736
rect 11526 8672 11542 8736
rect 11606 8672 11614 8736
rect 11294 7648 11614 8672
rect 11294 7584 11302 7648
rect 11366 7584 11382 7648
rect 11446 7584 11462 7648
rect 11526 7584 11542 7648
rect 11606 7584 11614 7648
rect 11294 6560 11614 7584
rect 11294 6496 11302 6560
rect 11366 6496 11382 6560
rect 11446 6496 11462 6560
rect 11526 6496 11542 6560
rect 11606 6496 11614 6560
rect 11294 5691 11614 6496
rect 11294 5472 11336 5691
rect 11572 5472 11614 5691
rect 11294 5408 11302 5472
rect 11366 5408 11382 5455
rect 11446 5408 11462 5455
rect 11526 5408 11542 5455
rect 11606 5408 11614 5472
rect 11294 4384 11614 5408
rect 11294 4320 11302 4384
rect 11366 4320 11382 4384
rect 11446 4320 11462 4384
rect 11526 4320 11542 4384
rect 11606 4320 11614 4384
rect 11294 3296 11614 4320
rect 11294 3232 11302 3296
rect 11366 3232 11382 3296
rect 11446 3232 11462 3296
rect 11526 3232 11542 3296
rect 11606 3232 11614 3296
rect 11294 2208 11614 3232
rect 11294 2144 11302 2208
rect 11366 2144 11382 2208
rect 11446 2144 11462 2208
rect 11526 2144 11542 2208
rect 11606 2144 11614 2208
rect 11294 2128 11614 2144
rect 14744 22336 15064 22896
rect 14744 22272 14752 22336
rect 14816 22272 14832 22336
rect 14896 22272 14912 22336
rect 14976 22272 14992 22336
rect 15056 22272 15064 22336
rect 14744 21248 15064 22272
rect 14744 21184 14752 21248
rect 14816 21184 14832 21248
rect 14896 21184 14912 21248
rect 14976 21184 14992 21248
rect 15056 21184 15064 21248
rect 14744 20160 15064 21184
rect 14744 20096 14752 20160
rect 14816 20096 14832 20160
rect 14896 20096 14912 20160
rect 14976 20096 14992 20160
rect 15056 20096 15064 20160
rect 14744 19072 15064 20096
rect 14744 19008 14752 19072
rect 14816 19008 14832 19072
rect 14896 19008 14912 19072
rect 14976 19008 14992 19072
rect 15056 19008 15064 19072
rect 14744 17984 15064 19008
rect 14744 17920 14752 17984
rect 14816 17920 14832 17984
rect 14896 17920 14912 17984
rect 14976 17920 14992 17984
rect 15056 17920 15064 17984
rect 14744 16896 15064 17920
rect 14744 16832 14752 16896
rect 14816 16832 14832 16896
rect 14896 16832 14912 16896
rect 14976 16832 14992 16896
rect 15056 16832 15064 16896
rect 14744 16027 15064 16832
rect 14744 15808 14786 16027
rect 15022 15808 15064 16027
rect 14744 15744 14752 15808
rect 14816 15744 14832 15791
rect 14896 15744 14912 15791
rect 14976 15744 14992 15791
rect 15056 15744 15064 15808
rect 14744 14720 15064 15744
rect 14744 14656 14752 14720
rect 14816 14656 14832 14720
rect 14896 14656 14912 14720
rect 14976 14656 14992 14720
rect 15056 14656 15064 14720
rect 14744 13632 15064 14656
rect 14744 13568 14752 13632
rect 14816 13568 14832 13632
rect 14896 13568 14912 13632
rect 14976 13568 14992 13632
rect 15056 13568 15064 13632
rect 14744 12544 15064 13568
rect 14744 12480 14752 12544
rect 14816 12480 14832 12544
rect 14896 12480 14912 12544
rect 14976 12480 14992 12544
rect 15056 12480 15064 12544
rect 14744 11456 15064 12480
rect 14744 11392 14752 11456
rect 14816 11392 14832 11456
rect 14896 11392 14912 11456
rect 14976 11392 14992 11456
rect 15056 11392 15064 11456
rect 14744 10368 15064 11392
rect 14744 10304 14752 10368
rect 14816 10304 14832 10368
rect 14896 10304 14912 10368
rect 14976 10304 14992 10368
rect 15056 10304 15064 10368
rect 14744 9280 15064 10304
rect 14744 9216 14752 9280
rect 14816 9216 14832 9280
rect 14896 9216 14912 9280
rect 14976 9216 14992 9280
rect 15056 9216 15064 9280
rect 14744 9136 15064 9216
rect 14744 8900 14786 9136
rect 15022 8900 15064 9136
rect 14744 8192 15064 8900
rect 14744 8128 14752 8192
rect 14816 8128 14832 8192
rect 14896 8128 14912 8192
rect 14976 8128 14992 8192
rect 15056 8128 15064 8192
rect 14744 7104 15064 8128
rect 14744 7040 14752 7104
rect 14816 7040 14832 7104
rect 14896 7040 14912 7104
rect 14976 7040 14992 7104
rect 15056 7040 15064 7104
rect 14744 6016 15064 7040
rect 14744 5952 14752 6016
rect 14816 5952 14832 6016
rect 14896 5952 14912 6016
rect 14976 5952 14992 6016
rect 15056 5952 15064 6016
rect 14744 4928 15064 5952
rect 14744 4864 14752 4928
rect 14816 4864 14832 4928
rect 14896 4864 14912 4928
rect 14976 4864 14992 4928
rect 15056 4864 15064 4928
rect 14744 3840 15064 4864
rect 14744 3776 14752 3840
rect 14816 3776 14832 3840
rect 14896 3776 14912 3840
rect 14976 3776 14992 3840
rect 15056 3776 15064 3840
rect 14744 2752 15064 3776
rect 14744 2688 14752 2752
rect 14816 2688 14832 2752
rect 14896 2688 14912 2752
rect 14976 2688 14992 2752
rect 15056 2688 15064 2752
rect 14744 2128 15064 2688
rect 18194 22880 18514 22896
rect 18194 22816 18202 22880
rect 18266 22816 18282 22880
rect 18346 22816 18362 22880
rect 18426 22816 18442 22880
rect 18506 22816 18514 22880
rect 18194 21792 18514 22816
rect 18194 21728 18202 21792
rect 18266 21728 18282 21792
rect 18346 21728 18362 21792
rect 18426 21728 18442 21792
rect 18506 21728 18514 21792
rect 18194 20704 18514 21728
rect 18194 20640 18202 20704
rect 18266 20640 18282 20704
rect 18346 20640 18362 20704
rect 18426 20640 18442 20704
rect 18506 20640 18514 20704
rect 18194 19616 18514 20640
rect 18194 19552 18202 19616
rect 18266 19552 18282 19616
rect 18346 19552 18362 19616
rect 18426 19552 18442 19616
rect 18506 19552 18514 19616
rect 18194 19472 18514 19552
rect 18194 19236 18236 19472
rect 18472 19236 18514 19472
rect 18194 18528 18514 19236
rect 18194 18464 18202 18528
rect 18266 18464 18282 18528
rect 18346 18464 18362 18528
rect 18426 18464 18442 18528
rect 18506 18464 18514 18528
rect 18194 17440 18514 18464
rect 18194 17376 18202 17440
rect 18266 17376 18282 17440
rect 18346 17376 18362 17440
rect 18426 17376 18442 17440
rect 18506 17376 18514 17440
rect 18194 16352 18514 17376
rect 18194 16288 18202 16352
rect 18266 16288 18282 16352
rect 18346 16288 18362 16352
rect 18426 16288 18442 16352
rect 18506 16288 18514 16352
rect 18194 15264 18514 16288
rect 18194 15200 18202 15264
rect 18266 15200 18282 15264
rect 18346 15200 18362 15264
rect 18426 15200 18442 15264
rect 18506 15200 18514 15264
rect 18194 14176 18514 15200
rect 18194 14112 18202 14176
rect 18266 14112 18282 14176
rect 18346 14112 18362 14176
rect 18426 14112 18442 14176
rect 18506 14112 18514 14176
rect 18194 13088 18514 14112
rect 18194 13024 18202 13088
rect 18266 13024 18282 13088
rect 18346 13024 18362 13088
rect 18426 13024 18442 13088
rect 18506 13024 18514 13088
rect 18194 12582 18514 13024
rect 18194 12346 18236 12582
rect 18472 12346 18514 12582
rect 18194 12000 18514 12346
rect 18194 11936 18202 12000
rect 18266 11936 18282 12000
rect 18346 11936 18362 12000
rect 18426 11936 18442 12000
rect 18506 11936 18514 12000
rect 18194 10912 18514 11936
rect 18194 10848 18202 10912
rect 18266 10848 18282 10912
rect 18346 10848 18362 10912
rect 18426 10848 18442 10912
rect 18506 10848 18514 10912
rect 18194 9824 18514 10848
rect 18194 9760 18202 9824
rect 18266 9760 18282 9824
rect 18346 9760 18362 9824
rect 18426 9760 18442 9824
rect 18506 9760 18514 9824
rect 18194 8736 18514 9760
rect 18194 8672 18202 8736
rect 18266 8672 18282 8736
rect 18346 8672 18362 8736
rect 18426 8672 18442 8736
rect 18506 8672 18514 8736
rect 18194 7648 18514 8672
rect 18194 7584 18202 7648
rect 18266 7584 18282 7648
rect 18346 7584 18362 7648
rect 18426 7584 18442 7648
rect 18506 7584 18514 7648
rect 18194 6560 18514 7584
rect 18194 6496 18202 6560
rect 18266 6496 18282 6560
rect 18346 6496 18362 6560
rect 18426 6496 18442 6560
rect 18506 6496 18514 6560
rect 18194 5691 18514 6496
rect 18194 5472 18236 5691
rect 18472 5472 18514 5691
rect 18194 5408 18202 5472
rect 18266 5408 18282 5455
rect 18346 5408 18362 5455
rect 18426 5408 18442 5455
rect 18506 5408 18514 5472
rect 18194 4384 18514 5408
rect 18194 4320 18202 4384
rect 18266 4320 18282 4384
rect 18346 4320 18362 4384
rect 18426 4320 18442 4384
rect 18506 4320 18514 4384
rect 18194 3296 18514 4320
rect 18194 3232 18202 3296
rect 18266 3232 18282 3296
rect 18346 3232 18362 3296
rect 18426 3232 18442 3296
rect 18506 3232 18514 3296
rect 18194 2208 18514 3232
rect 18194 2144 18202 2208
rect 18266 2144 18282 2208
rect 18346 2144 18362 2208
rect 18426 2144 18442 2208
rect 18506 2144 18514 2208
rect 18194 2128 18514 2144
<< via4 >>
rect 4436 19236 4672 19472
rect 4436 12346 4672 12582
rect 4436 5472 4672 5691
rect 4436 5455 4466 5472
rect 4466 5455 4482 5472
rect 4482 5455 4546 5472
rect 4546 5455 4562 5472
rect 4562 5455 4626 5472
rect 4626 5455 4642 5472
rect 4642 5455 4672 5472
rect 7886 15808 8122 16027
rect 7886 15791 7916 15808
rect 7916 15791 7932 15808
rect 7932 15791 7996 15808
rect 7996 15791 8012 15808
rect 8012 15791 8076 15808
rect 8076 15791 8092 15808
rect 8092 15791 8122 15808
rect 7886 8900 8122 9136
rect 11336 19236 11572 19472
rect 11336 12346 11572 12582
rect 11336 5472 11572 5691
rect 11336 5455 11366 5472
rect 11366 5455 11382 5472
rect 11382 5455 11446 5472
rect 11446 5455 11462 5472
rect 11462 5455 11526 5472
rect 11526 5455 11542 5472
rect 11542 5455 11572 5472
rect 14786 15808 15022 16027
rect 14786 15791 14816 15808
rect 14816 15791 14832 15808
rect 14832 15791 14896 15808
rect 14896 15791 14912 15808
rect 14912 15791 14976 15808
rect 14976 15791 14992 15808
rect 14992 15791 15022 15808
rect 14786 8900 15022 9136
rect 18236 19236 18472 19472
rect 18236 12346 18472 12582
rect 18236 5472 18472 5691
rect 18236 5455 18266 5472
rect 18266 5455 18282 5472
rect 18282 5455 18346 5472
rect 18346 5455 18362 5472
rect 18362 5455 18426 5472
rect 18426 5455 18442 5472
rect 18442 5455 18472 5472
<< metal5 >>
rect 1104 19472 21804 19515
rect 1104 19236 4436 19472
rect 4672 19236 11336 19472
rect 11572 19236 18236 19472
rect 18472 19236 21804 19472
rect 1104 19194 21804 19236
rect 1104 16027 21804 16069
rect 1104 15791 7886 16027
rect 8122 15791 14786 16027
rect 15022 15791 21804 16027
rect 1104 15749 21804 15791
rect 1104 12582 21804 12624
rect 1104 12346 4436 12582
rect 4672 12346 11336 12582
rect 11572 12346 18236 12582
rect 18472 12346 21804 12582
rect 1104 12304 21804 12346
rect 1104 9136 21804 9179
rect 1104 8900 7886 9136
rect 8122 8900 14786 9136
rect 15022 8900 21804 9136
rect 1104 8858 21804 8900
rect 1104 5691 21804 5733
rect 1104 5455 4436 5691
rect 4672 5455 11336 5691
rect 11572 5455 18236 5691
rect 18472 5455 21804 5691
rect 1104 5413 21804 5455
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1618419204
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1618419204
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1619507013
transform 1 0 1840 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output83 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 2208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp 1618419204
transform 1 0 1748 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12
timestamp 1618419204
transform 1 0 2208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_11
timestamp 1618419204
transform 1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 2852 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input43 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 2576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1619507013
transform 1 0 2484 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 2760 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 3864 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37
timestamp 1618419204
transform 1 0 4508 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30
timestamp 1618419204
transform 1 0 3864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1618419204
transform -1 0 4508 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1618419204
transform -1 0 4692 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45
timestamp 1618419204
transform 1 0 5244 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1618419204
transform -1 0 5796 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1618419204
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_58
timestamp 1618419204
transform 1 0 6440 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_51
timestamp 1618419204
transform 1 0 5796 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1618419204
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1618419204
transform 1 0 6348 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51
timestamp 1618419204
transform 1 0 5796 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1618419204
transform -1 0 7084 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1618419204
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1618419204
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1618419204
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_65
timestamp 1618419204
transform 1 0 7084 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_66
timestamp 1618419204
transform 1 0 7176 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_81
timestamp 1618419204
transform 1 0 8556 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_77
timestamp 1618419204
transform 1 0 8188 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1618419204
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78
timestamp 1618419204
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1618419204
transform -1 0 8740 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 8924 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_94
timestamp 1618419204
transform 1 0 9752 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_85
timestamp 1618419204
transform 1 0 8924 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1618419204
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1618419204
transform -1 0 9844 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1618419204
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[11\].id.delayen1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 9752 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_1_98
timestamp 1618419204
transform 1 0 10120 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95
timestamp 1618419204
transform 1 0 9844 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _355_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 10212 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_1_108
timestamp 1618419204
transform 1 0 11040 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_105
timestamp 1618419204
transform 1 0 10764 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101
timestamp 1618419204
transform 1 0 10396 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1618419204
transform -1 0 10764 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1618419204
transform -1 0 11408 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_115
timestamp 1618419204
transform 1 0 11684 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117
timestamp 1618419204
transform 1 0 11868 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1618419204
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1618419204
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1618419204
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_123
timestamp 1618419204
transform 1 0 12420 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp 1618419204
transform -1 0 13340 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_125
timestamp 1618419204
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen1
timestamp 1618419204
transform 1 0 12788 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_1_133
timestamp 1618419204
transform 1 0 13340 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_132
timestamp 1618419204
transform 1 0 13248 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[9\].id.delayenb1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 13708 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1618419204
transform 1 0 13616 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_142
timestamp 1618419204
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_139
timestamp 1618419204
transform 1 0 13892 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp 1618419204
transform 1 0 14812 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_146
timestamp 1618419204
transform 1 0 14536 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1618419204
transform 1 0 14536 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1618419204
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_157
timestamp 1618419204
transform 1 0 15548 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_152
timestamp 1618419204
transform 1 0 15088 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1619507013
transform 1 0 15916 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1618419204
transform 1 0 15180 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1618419204
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_165
timestamp 1618419204
transform 1 0 16284 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_172
timestamp 1618419204
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_164
timestamp 1618419204
transform 1 0 16192 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1618419204
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 16284 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1618419204
transform 1 0 17664 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_182
timestamp 1618419204
transform 1 0 17848 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1618419204
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1618419204
transform 1 0 17572 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1618419204
transform -1 0 17664 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1618419204
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1618419204
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_196
timestamp 1618419204
transform 1 0 19136 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_190
timestamp 1618419204
transform 1 0 18584 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1618419204
transform 1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_187
timestamp 1618419204
transform 1 0 18308 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_205
timestamp 1618419204
transform 1 0 19964 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_199
timestamp 1618419204
transform 1 0 19412 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_204
timestamp 1618419204
transform 1 0 19872 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_202
timestamp 1618419204
transform 1 0 19688 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1618419204
transform -1 0 20332 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1618419204
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_216
timestamp 1618419204
transform 1 0 20976 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_209
timestamp 1618419204
transform 1 0 20332 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_212
timestamp 1618419204
transform 1 0 20608 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1618419204
transform -1 0 21068 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1618419204
transform 1 0 20700 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_221
timestamp 1618419204
transform 1 0 21436 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_217
timestamp 1618419204
transform 1 0 21068 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1618419204
transform -1 0 21804 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1618419204
transform -1 0 21804 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1618419204
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1618419204
transform -1 0 1656 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_6
timestamp 1618419204
transform 1 0 1656 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1618419204
transform 1 0 2760 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1618419204
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_26
timestamp 1618419204
transform 1 0 3496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1618419204
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_42
timestamp 1618419204
transform 1 0 4968 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_4  ringosc.dstage\[11\].id.delayen0
timestamp 1619507013
transform 1 0 7636 0 -1 3808
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1618419204
transform -1 0 6348 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_50
timestamp 1618419204
transform 1 0 5704 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_57
timestamp 1618419204
transform 1 0 6348 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_69
timestamp 1618419204
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[11\].id.delayenb1
timestamp 1618419204
transform -1 0 9936 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1618419204
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_82
timestamp 1618419204
transform 1 0 8648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1618419204
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_96
timestamp 1618419204
transform 1 0 9936 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1618419204
transform 1 0 10304 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1618419204
transform 1 0 11224 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1618419204
transform 1 0 11960 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_103
timestamp 1618419204
transform 1 0 10580 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_109
timestamp 1618419204
transform 1 0 11132 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_113
timestamp 1618419204
transform 1 0 11500 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_117
timestamp 1618419204
transform 1 0 11868 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_121
timestamp 1618419204
transform 1 0 12236 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1618419204
transform 1 0 14720 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen0
timestamp 1618419204
transform -1 0 13800 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1618419204
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_138
timestamp 1618419204
transform 1 0 13800 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_142
timestamp 1618419204
transform 1 0 14168 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_144
timestamp 1618419204
transform 1 0 14352 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_157
timestamp 1618419204
transform 1 0 15548 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_169
timestamp 1618419204
transform 1 0 16652 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_181
timestamp 1618419204
transform 1 0 17756 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_193
timestamp 1618419204
transform 1 0 18860 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1618419204
transform -1 0 21804 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1618419204
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1618419204
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_199
timestamp 1618419204
transform 1 0 19412 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_201
timestamp 1618419204
transform 1 0 19596 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_213
timestamp 1618419204
transform 1 0 20700 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_218
timestamp 1618419204
transform 1 0 21160 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1618419204
transform 1 0 3220 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1618419204
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output45
timestamp 1618419204
transform 1 0 1840 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1618419204
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1618419204
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_11
timestamp 1618419204
transform 1 0 2116 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1618419204
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1618419204
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1618419204
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1618419204
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1618419204
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_70
timestamp 1618419204
transform 1 0 7544 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_74
timestamp 1618419204
transform 1 0 7912 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb0
timestamp 1619507013
transform 1 0 8004 0 1 3808
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1618419204
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_98
timestamp 1618419204
transform 1 0 10120 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1618419204
transform -1 0 12328 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1618419204
transform -1 0 10948 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1618419204
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_102
timestamp 1618419204
transform 1 0 10488 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_107
timestamp 1618419204
transform 1 0 10948 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1618419204
transform 1 0 11500 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1618419204
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_122
timestamp 1618419204
transform 1 0 12328 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[9\].id.delayenb0
timestamp 1618419204
transform -1 0 13708 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1618419204
transform 1 0 14076 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_130
timestamp 1618419204
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_137
timestamp 1618419204
transform 1 0 13708 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_144
timestamp 1618419204
transform 1 0 14352 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1619507013
transform 1 0 16192 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1618419204
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_156
timestamp 1618419204
transform 1 0 15456 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_167
timestamp 1618419204
transform 1 0 16468 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_172
timestamp 1618419204
transform 1 0 16928 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1618419204
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1618419204
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1618419204
transform -1 0 21804 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output43
timestamp 1618419204
transform -1 0 20516 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_211
timestamp 1618419204
transform 1 0 20516 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_219
timestamp 1618419204
transform 1 0 21252 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1618419204
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1618419204
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1618419204
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_4  irb
timestamp 1619507013
transform -1 0 5980 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1618419204
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1618419204
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1618419204
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_42
timestamp 1618419204
transform 1 0 4968 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1
timestamp 1619507013
transform 1 0 6624 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_53
timestamp 1618419204
transform 1 0 5980 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_59
timestamp 1618419204
transform 1 0 6532 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_63
timestamp 1618419204
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _356_
timestamp 1618419204
transform -1 0 10948 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1618419204
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_75
timestamp 1618419204
transform 1 0 8004 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_83
timestamp 1618419204
transform 1 0 8740 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_87
timestamp 1618419204
transform 1 0 9108 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_95
timestamp 1618419204
transform 1 0 9844 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen0
timestamp 1618419204
transform 1 0 11316 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[10\].id.delayenb0
timestamp 1618419204
transform 1 0 12144 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_4_107
timestamp 1618419204
transform 1 0 10948 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_116
timestamp 1618419204
transform 1 0 11776 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  ringosc.dstage\[10\].id.delaybuf0
timestamp 1619507013
transform -1 0 13340 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1618419204
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_125
timestamp 1618419204
transform 1 0 12604 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_129
timestamp 1618419204
transform 1 0 12972 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_133
timestamp 1618419204
transform 1 0 13340 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1618419204
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144
timestamp 1618419204
transform 1 0 14352 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__nor3_2  _324_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 16744 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_156
timestamp 1618419204
transform 1 0 15456 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_170
timestamp 1618419204
transform 1 0 16744 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _325_
timestamp 1618419204
transform 1 0 17112 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_182
timestamp 1618419204
transform 1 0 17848 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_194
timestamp 1618419204
transform 1 0 18952 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1618419204
transform -1 0 21804 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1618419204
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_201
timestamp 1618419204
transform 1 0 19596 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_213
timestamp 1618419204
transform 1 0 20700 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_221
timestamp 1618419204
transform 1 0 21436 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfrbp_2  idiv4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 2484 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1618419204
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output41
timestamp 1618419204
transform 1 0 1748 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1618419204
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_10
timestamp 1618419204
transform 1 0 2024 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_14
timestamp 1618419204
transform 1 0 2392 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 5980 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_5_39
timestamp 1618419204
transform 1 0 4692 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_45
timestamp 1618419204
transform 1 0 5244 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 7176 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1618419204
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_53
timestamp 1618419204
transform 1 0 5980 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_58
timestamp 1618419204
transform 1 0 6440 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_66
timestamp 1618419204
transform 1 0 7176 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1618419204
transform -1 0 9844 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_1  ringosc.iss.delayenb1
timestamp 1618419204
transform -1 0 9200 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1618419204
transform 1 0 8280 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_82
timestamp 1618419204
transform 1 0 8648 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_88
timestamp 1618419204
transform 1 0 9200 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_95
timestamp 1618419204
transform 1 0 9844 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen1
timestamp 1618419204
transform 1 0 12052 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1618419204
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_107
timestamp 1618419204
transform 1 0 10948 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1618419204
transform 1 0 11500 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_115
timestamp 1618419204
transform 1 0 11684 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_124
timestamp 1618419204
transform 1 0 12512 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1618419204
transform 1 0 12880 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_131
timestamp 1618419204
transform 1 0 13156 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_143
timestamp 1618419204
transform 1 0 14260 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__nor3_2  _323_
timestamp 1618419204
transform -1 0 16376 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1618419204
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_155
timestamp 1618419204
transform 1 0 15364 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_166
timestamp 1618419204
transform 1 0 16376 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_170
timestamp 1618419204
transform 1 0 16744 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_172
timestamp 1618419204
transform 1 0 16928 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1619507013
transform -1 0 17572 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfrbp_1  idiv16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 20240 0 1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_6  FILLER_5_179
timestamp 1618419204
transform 1 0 17572 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1618419204
transform -1 0 21804 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1618419204
transform 1 0 20884 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_208
timestamp 1618419204
transform 1 0 20240 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_214
timestamp 1618419204
transform 1 0 20792 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_218
timestamp 1618419204
transform 1 0 21160 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrbp_2  idiv2
timestamp 1618419204
transform 1 0 2392 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1618419204
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1618419204
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1618419204
transform -1 0 1748 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_7
timestamp 1618419204
transform 1 0 1748 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_19
timestamp 1618419204
transform 1 0 2852 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1618419204
transform 1 0 1380 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_11
timestamp 1618419204
transform 1 0 2116 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1618419204
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1618419204
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1618419204
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_42
timestamp 1618419204
transform 1 0 4968 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_38
timestamp 1618419204
transform 1 0 4600 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_58
timestamp 1618419204
transform 1 0 6440 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_56
timestamp 1618419204
transform 1 0 6256 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1618419204
transform 1 0 5704 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_50
timestamp 1618419204
transform 1 0 5704 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1618419204
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.reseten0
timestamp 1619507013
transform 1 0 5888 0 -1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_7_72
timestamp 1618419204
transform 1 0 7728 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_66
timestamp 1618419204
transform 1 0 7176 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_63
timestamp 1618419204
transform 1 0 6900 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb0
timestamp 1619507013
transform 1 0 7636 0 -1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__or2_1  ringosc.iss.ctrlen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 7728 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1618419204
transform 1 0 9568 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.delayen0
timestamp 1619507013
transform 1 0 8188 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.delayen1
timestamp 1618419204
transform 1 0 9476 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1618419204
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_82
timestamp 1618419204
transform 1 0 8648 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1618419204
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_96
timestamp 1618419204
transform 1 0 9936 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_76
timestamp 1618419204
transform 1 0 8096 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_88
timestamp 1618419204
transform 1 0 9200 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1618419204
transform 1 0 10304 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_123
timestamp 1618419204
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_119
timestamp 1618419204
transform 1 0 12052 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_115
timestamp 1618419204
transform 1 0 11684 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 1618419204
transform 1 0 11500 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_115
timestamp 1618419204
transform 1 0 11684 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1618419204
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[10\].id.delayenb1
timestamp 1618419204
transform 1 0 11868 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  ringosc.dstage\[0\].id.delaybuf0
timestamp 1619507013
transform 1 0 12144 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_101
timestamp 1618419204
transform 1 0 10396 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_122
timestamp 1618419204
transform 1 0 12328 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_103
timestamp 1618419204
transform 1 0 10580 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_132
timestamp 1618419204
transform 1 0 13248 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_134
timestamp 1618419204
transform 1 0 13432 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[0\].id.delayenb1
timestamp 1618419204
transform 1 0 12788 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_7_139
timestamp 1618419204
transform 1 0 13892 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_142
timestamp 1618419204
transform 1 0 14168 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1618419204
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 1618419204
transform 1 0 13616 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1618419204
transform 1 0 14260 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_148
timestamp 1618419204
transform 1 0 14720 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_144
timestamp 1618419204
transform 1 0 14352 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1618419204
transform 1 0 14812 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_152
timestamp 1618419204
transform 1 0 15088 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_158
timestamp 1618419204
transform 1 0 15640 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _322_
timestamp 1618419204
transform -1 0 16192 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_164
timestamp 1618419204
transform 1 0 16192 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_162
timestamp 1618419204
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1618419204
transform 1 0 16100 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_7_172
timestamp 1618419204
transform 1 0 16928 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_170
timestamp 1618419204
transform 1 0 16744 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_172
timestamp 1618419204
transform 1 0 16928 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1618419204
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1618419204
transform 1 0 17296 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfrbp_1  idiv8
timestamp 1618419204
transform 1 0 17664 0 1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_12  FILLER_6_185
timestamp 1618419204
transform 1 0 18124 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp 1618419204
transform 1 0 19228 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_211
timestamp 1618419204
transform 1 0 20516 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_203
timestamp 1618419204
transform 1 0 19780 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1618419204
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_216
timestamp 1618419204
transform 1 0 20976 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_216
timestamp 1618419204
transform 1 0 20976 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1618419204
transform 1 0 20700 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1619507013
transform -1 0 20976 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1618419204
transform -1 0 21804 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1618419204
transform -1 0 21804 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_201
timestamp 1618419204
transform 1 0 19596 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1618419204
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output39
timestamp 1618419204
transform 1 0 1748 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output40
timestamp 1618419204
transform 1 0 2392 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1618419204
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_10
timestamp 1618419204
transform 1 0 2024 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_17
timestamp 1618419204
transform 1 0 2668 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _377_
timestamp 1618419204
transform -1 0 5428 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1618419204
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_30
timestamp 1618419204
transform 1 0 3864 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_47
timestamp 1618419204
transform 1 0 5428 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 6992 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_8_64
timestamp 1618419204
transform 1 0 6992 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1618419204
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 1618419204
transform 1 0 8096 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1618419204
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1618419204
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_99
timestamp 1618419204
transform 1 0 10212 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _368_
timestamp 1618419204
transform 1 0 10856 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_105
timestamp 1618419204
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_115
timestamp 1618419204
transform 1 0 11684 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1618419204
transform 1 0 13616 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen1
timestamp 1618419204
transform 1 0 12788 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1618419204
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_132
timestamp 1618419204
transform 1 0 13248 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_139
timestamp 1618419204
transform 1 0 13892 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1618419204
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_156
timestamp 1618419204
transform 1 0 15456 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_168
timestamp 1618419204
transform 1 0 16560 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_180
timestamp 1618419204
transform 1 0 17664 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_192
timestamp 1618419204
transform 1 0 18768 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1618419204
transform -1 0 21804 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1618419204
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  output42
timestamp 1619507013
transform 1 0 20700 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_201
timestamp 1618419204
transform 1 0 19596 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_216
timestamp 1618419204
transform 1 0 20976 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  ringosc.ibufp11
timestamp 1619507013
transform -1 0 3036 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1618419204
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1618419204
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_15
timestamp 1618419204
transform 1 0 2484 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_21
timestamp 1618419204
transform 1 0 3036 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_8  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 4508 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_33
timestamp 1618419204
transform 1 0 4140 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1618419204
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_53
timestamp 1618419204
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1618419204
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_70
timestamp 1618419204
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen1
timestamp 1618419204
transform 1 0 9844 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_9_82
timestamp 1618419204
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_94
timestamp 1618419204
transform 1 0 9752 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen0
timestamp 1618419204
transform 1 0 10672 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[4\].id.delayenb1
timestamp 1618419204
transform -1 0 12512 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1618419204
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_100
timestamp 1618419204
transform 1 0 10304 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_109
timestamp 1618419204
transform 1 0 11132 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1618419204
transform 1 0 11500 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_115
timestamp 1618419204
transform 1 0 11684 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_124
timestamp 1618419204
transform 1 0 12512 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen0
timestamp 1618419204
transform -1 0 14168 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[0\].id.delayenb0
timestamp 1618419204
transform -1 0 13340 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_9_133
timestamp 1618419204
transform 1 0 13340 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_142
timestamp 1618419204
transform 1 0 14168 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1618419204
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_154
timestamp 1618419204
transform 1 0 15272 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_166
timestamp 1618419204
transform 1 0 16376 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_170
timestamp 1618419204
transform 1 0 16744 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_172
timestamp 1618419204
transform 1 0 16928 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1618419204
transform -1 0 17848 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_182
timestamp 1618419204
transform 1 0 17848 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_194
timestamp 1618419204
transform 1 0 18952 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1618419204
transform -1 0 21804 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_206
timestamp 1618419204
transform 1 0 20056 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_218
timestamp 1618419204
transform 1 0 21160 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1618419204
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1618419204
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1618419204
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1618419204
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1618419204
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1618419204
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1618419204
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  ringosc.dstage\[5\].id.delaybuf0
timestamp 1619507013
transform -1 0 6348 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  repeater46
timestamp 1619507013
transform -1 0 8372 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_57
timestamp 1618419204
transform 1 0 6348 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_69
timestamp 1618419204
transform 1 0 7452 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _369_
timestamp 1618419204
transform -1 0 10304 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1618419204
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_79
timestamp 1618419204
transform 1 0 8372 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1618419204
transform 1 0 8924 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1618419204
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1618419204
transform 1 0 11776 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb0
timestamp 1619507013
transform 1 0 10764 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_10_100
timestamp 1618419204
transform 1 0 10304 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_104
timestamp 1618419204
transform 1 0 10672 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_112
timestamp 1618419204
transform 1 0 11408 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_119
timestamp 1618419204
transform 1 0 12052 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _347_
timestamp 1618419204
transform -1 0 13064 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  ringosc.dstage\[1\].id.delaybuf0
timestamp 1619507013
transform 1 0 14812 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1618419204
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_130
timestamp 1618419204
transform 1 0 13064 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_142
timestamp 1618419204
transform 1 0 14168 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_144
timestamp 1618419204
transform 1 0 14352 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_148
timestamp 1618419204
transform 1 0 14720 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp 1618419204
transform 1 0 15456 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_152
timestamp 1618419204
transform 1 0 15088 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1618419204
transform 1 0 16284 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1618419204
transform 1 0 17388 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_189
timestamp 1618419204
transform 1 0 18492 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp 1618419204
transform 1 0 19228 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1618419204
transform -1 0 21804 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1618419204
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1618419204
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1618419204
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_213
timestamp 1618419204
transform 1 0 20700 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_218
timestamp 1618419204
transform 1 0 21160 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb0
timestamp 1619507013
transform 1 0 2116 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__inv_1  ringosc.ibufp10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 3496 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1618419204
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1618419204
transform -1 0 1748 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1618419204
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_7
timestamp 1618419204
transform 1 0 1748 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_18
timestamp 1618419204
transform 1 0 2760 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_22
timestamp 1618419204
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1618419204
transform -1 0 5060 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_26
timestamp 1618419204
transform 1 0 3496 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_38
timestamp 1618419204
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_43
timestamp 1618419204
transform 1 0 5060 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1618419204
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_55
timestamp 1618419204
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1618419204
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_70
timestamp 1618419204
transform 1 0 7544 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _321_
timestamp 1619507013
transform -1 0 9936 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_82
timestamp 1618419204
transform 1 0 8648 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_96
timestamp 1618419204
transform 1 0 9936 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1618419204
transform 1 0 10948 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1618419204
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_104
timestamp 1618419204
transform 1 0 10672 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_110
timestamp 1618419204
transform 1 0 11224 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_115
timestamp 1618419204
transform 1 0 11684 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1618419204
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1618419204
transform 1 0 12604 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[1\].id.delayenb1
timestamp 1618419204
transform 1 0 14536 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_11_134
timestamp 1618419204
transform 1 0 13432 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1618419204
transform 1 0 16192 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen1
timestamp 1618419204
transform 1 0 15364 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1618419204
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_151
timestamp 1618419204
transform 1 0 14996 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_160
timestamp 1618419204
transform 1 0 15824 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_167
timestamp 1618419204
transform 1 0 16468 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_172
timestamp 1618419204
transform 1 0 16928 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1618419204
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1618419204
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1618419204
transform -1 0 21804 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1618419204
transform 1 0 20700 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_208
timestamp 1618419204
transform 1 0 20240 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_212
timestamp 1618419204
transform 1 0 20608 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_216
timestamp 1618419204
transform 1 0 20976 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _360_
timestamp 1618419204
transform 1 0 2024 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1618419204
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1618419204
transform -1 0 1656 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_6
timestamp 1618419204
transform 1 0 1656 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_19
timestamp 1618419204
transform 1 0 2852 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[5\].id.delayen1
timestamp 1618419204
transform -1 0 5704 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[5\].id.delayenb0
timestamp 1619507013
transform 1 0 4232 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1618419204
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1618419204
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_30
timestamp 1618419204
transform 1 0 3864 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_41
timestamp 1618419204
transform 1 0 4876 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _354_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 7820 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1618419204
transform 1 0 6072 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_50
timestamp 1618419204
transform 1 0 5704 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_57
timestamp 1618419204
transform 1 0 6348 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_63
timestamp 1618419204
transform 1 0 6900 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_73
timestamp 1618419204
transform 1 0 7820 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1618419204
transform 1 0 9476 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1618419204
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1618419204
transform 1 0 8924 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1618419204
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _306_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 11132 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  ringosc.dstage\[4\].id.delaybuf0
timestamp 1619507013
transform -1 0 12144 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_100
timestamp 1618419204
transform 1 0 10304 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_109
timestamp 1618419204
transform 1 0 11132 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_120
timestamp 1618419204
transform 1 0 12144 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1618419204
transform 1 0 12696 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1618419204
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_135
timestamp 1618419204
transform 1 0 13524 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_144
timestamp 1618419204
transform 1 0 14352 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen0
timestamp 1618419204
transform 1 0 15272 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1618419204
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_152
timestamp 1618419204
transform 1 0 15088 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_159
timestamp 1618419204
transform 1 0 15732 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1618419204
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1618419204
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_190
timestamp 1618419204
transform 1 0 18584 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_198
timestamp 1618419204
transform 1 0 19320 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1618419204
transform -1 0 21804 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1618419204
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1618419204
transform 1 0 20700 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1618419204
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_216
timestamp 1618419204
transform 1 0 20976 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_7
timestamp 1618419204
transform 1 0 1748 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1618419204
transform 1 0 1380 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1618419204
transform -1 0 1748 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1618419204
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1618419204
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1619507013
transform 1 0 2116 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_14_23
timestamp 1618419204
transform 1 0 3220 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_16
timestamp 1618419204
transform 1 0 2576 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1618419204
transform 1 0 2944 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1618419204
transform 1 0 2300 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_18
timestamp 1618419204
transform 1 0 2760 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1618419204
transform 1 0 5520 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1619507013
transform 1 0 4140 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[5\].id.delayenb1
timestamp 1618419204
transform -1 0 5612 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1618419204
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_30
timestamp 1618419204
transform 1 0 3864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_40
timestamp 1618419204
transform 1 0 4784 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_49
timestamp 1618419204
transform 1 0 5612 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1618419204
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_42
timestamp 1618419204
transform 1 0 4968 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 7268 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 7912 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _372_
timestamp 1618419204
transform -1 0 7544 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1618419204
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_58
timestamp 1618419204
transform 1 0 6440 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_66
timestamp 1618419204
transform 1 0 7176 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_73
timestamp 1618419204
transform 1 0 7820 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_57
timestamp 1618419204
transform 1 0 6348 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_70
timestamp 1618419204
transform 1 0 7544 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1618419204
transform 1 0 8924 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_81
timestamp 1618419204
transform 1 0 8556 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_86
timestamp 1618419204
transform 1 0 9016 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1618419204
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1618419204
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1619507013
transform -1 0 9016 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_94
timestamp 1618419204
transform 1 0 9752 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_87
timestamp 1618419204
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_92
timestamp 1618419204
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _319_
timestamp 1619507013
transform 1 0 9660 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1619507013
transform 1 0 9476 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_99
timestamp 1618419204
transform 1 0 10212 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _291_
timestamp 1618419204
transform 1 0 12052 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _312_
timestamp 1619507013
transform -1 0 10948 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1618419204
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_111
timestamp 1618419204
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1618419204
transform 1 0 11684 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_124
timestamp 1618419204
transform 1 0 12512 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_100
timestamp 1618419204
transform 1 0 10304 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_107
timestamp 1618419204
transform 1 0 10948 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_119
timestamp 1618419204
transform 1 0 12052 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen0
timestamp 1618419204
transform -1 0 13340 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[3\].id.delayenb0
timestamp 1618419204
transform 1 0 12604 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1618419204
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_133
timestamp 1618419204
transform 1 0 13340 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_145
timestamp 1618419204
transform 1 0 14444 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_130
timestamp 1618419204
transform 1 0 13064 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_142
timestamp 1618419204
transform 1 0 14168 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_144
timestamp 1618419204
transform 1 0 14352 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[1\].id.delayenb0
timestamp 1618419204
transform 1 0 15088 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  ringosc.dstage\[2\].id.delaybuf0
timestamp 1619507013
transform 1 0 15732 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1618419204
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_151
timestamp 1618419204
transform 1 0 14996 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_157
timestamp 1618419204
transform 1 0 15548 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1618419204
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1618419204
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_156
timestamp 1618419204
transform 1 0 15456 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_162
timestamp 1618419204
transform 1 0 16008 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1618419204
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1618419204
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_174
timestamp 1618419204
transform 1 0 17112 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_186
timestamp 1618419204
transform 1 0 18216 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_198
timestamp 1618419204
transform 1 0 19320 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1618419204
transform -1 0 21804 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1618419204
transform -1 0 21804 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1618419204
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1618419204
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1618419204
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_220
timestamp 1618419204
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1618419204
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_213
timestamp 1618419204
transform 1 0 20700 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_218
timestamp 1618419204
transform 1 0 21160 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen1
timestamp 1618419204
transform 1 0 1840 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[8\].id.delayenb1
timestamp 1618419204
transform -1 0 3128 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1618419204
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1618419204
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1618419204
transform 1 0 1748 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1618419204
transform 1 0 2300 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_22
timestamp 1618419204
transform 1 0 3128 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  ringosc.dstage\[6\].id.delaybuf0
timestamp 1619507013
transform -1 0 4048 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_28
timestamp 1618419204
transform 1 0 3680 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_32
timestamp 1618419204
transform 1 0 4048 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1618419204
transform 1 0 5152 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1618419204
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_56
timestamp 1618419204
transform 1 0 6256 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_58
timestamp 1618419204
transform 1 0 6440 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_70
timestamp 1618419204
transform 1 0 7544 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _300_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 8096 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _301_
timestamp 1618419204
transform 1 0 8832 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _302_
timestamp 1618419204
transform 1 0 9568 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_80
timestamp 1618419204
transform 1 0 8464 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_88
timestamp 1618419204
transform 1 0 9200 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_96
timestamp 1618419204
transform 1 0 9936 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _315_
timestamp 1619507013
transform -1 0 10764 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1618419204
transform -1 0 12696 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1618419204
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_105
timestamp 1618419204
transform 1 0 10764 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1618419204
transform 1 0 11500 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_115
timestamp 1618419204
transform 1 0 11684 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1618419204
transform -1 0 13892 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  ringosc.dstage\[3\].id.delaybuf0
timestamp 1619507013
transform -1 0 14720 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_126
timestamp 1618419204
transform 1 0 12696 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_139
timestamp 1618419204
transform 1 0 13892 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_148
timestamp 1618419204
transform 1 0 14720 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen0
timestamp 1618419204
transform -1 0 15548 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[2\].id.delayenb0
timestamp 1618419204
transform 1 0 15916 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1618419204
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_157
timestamp 1618419204
transform 1 0 15548 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_166
timestamp 1618419204
transform 1 0 16376 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_170
timestamp 1618419204
transform 1 0 16744 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_172
timestamp 1618419204
transform 1 0 16928 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1618419204
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1618419204
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1618419204
transform -1 0 21804 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1618419204
transform 1 0 20700 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_208
timestamp 1618419204
transform 1 0 20240 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_212
timestamp 1618419204
transform 1 0 20608 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_216
timestamp 1618419204
transform 1 0 20976 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  ringosc.dstage\[8\].id.delaybuf0
timestamp 1619507013
transform 1 0 2208 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1618419204
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1618419204
transform 1 0 1380 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_11
timestamp 1618419204
transform 1 0 2116 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1618419204
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _366_
timestamp 1618419204
transform 1 0 5152 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen1
timestamp 1618419204
transform -1 0 4692 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1618419204
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1618419204
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_30
timestamp 1618419204
transform 1 0 3864 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_39
timestamp 1618419204
transform 1 0 4692 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_43
timestamp 1618419204
transform 1 0 5060 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _304_
timestamp 1618419204
transform 1 0 6348 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _308_
timestamp 1618419204
transform 1 0 7360 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_16_53
timestamp 1618419204
transform 1 0 5980 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_64
timestamp 1618419204
transform 1 0 6992 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1619507013
transform 1 0 8372 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _311_
timestamp 1619507013
transform 1 0 9568 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1618419204
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_75
timestamp 1618419204
transform 1 0 8004 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_82
timestamp 1618419204
transform 1 0 8648 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1618419204
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1618419204
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _365_
timestamp 1618419204
transform 1 0 11224 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_101
timestamp 1618419204
transform 1 0 10396 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_109
timestamp 1618419204
transform 1 0 11132 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_119
timestamp 1618419204
transform 1 0 12052 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen1
timestamp 1618419204
transform 1 0 12880 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1618419204
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_127
timestamp 1618419204
transform 1 0 12788 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_133
timestamp 1618419204
transform 1 0 13340 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1618419204
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_144
timestamp 1618419204
transform 1 0 14352 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen1
timestamp 1618419204
transform 1 0 15548 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[2\].id.delayenb1
timestamp 1618419204
transform 1 0 16376 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1618419204
transform -1 0 15180 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_153
timestamp 1618419204
transform 1 0 15180 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_162
timestamp 1618419204
transform 1 0 16008 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_171
timestamp 1618419204
transform 1 0 16836 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1618419204
transform 1 0 17204 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1618419204
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_190
timestamp 1618419204
transform 1 0 18584 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_198
timestamp 1618419204
transform 1 0 19320 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1618419204
transform -1 0 21804 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1618419204
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_201
timestamp 1618419204
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_213
timestamp 1618419204
transform 1 0 20700 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_221
timestamp 1618419204
transform 1 0 21436 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1618419204
transform -1 0 2668 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1618419204
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1618419204
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1618419204
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_17
timestamp 1618419204
transform 1 0 2668 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _314_
timestamp 1619507013
transform 1 0 5428 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1618419204
transform 1 0 4324 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[6\].id.delayenb1
timestamp 1618419204
transform -1 0 3956 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_17_25
timestamp 1618419204
transform 1 0 3404 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_31
timestamp 1618419204
transform 1 0 3956 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_38
timestamp 1618419204
transform 1 0 4600 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_46
timestamp 1618419204
transform 1 0 5336 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _296_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 7268 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1618419204
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_53
timestamp 1618419204
transform 1 0 5980 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_58
timestamp 1618419204
transform 1 0 6440 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_67
timestamp 1618419204
transform 1 0 7268 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _298_
timestamp 1618419204
transform -1 0 9108 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_17_79
timestamp 1618419204
transform 1 0 8372 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_87
timestamp 1618419204
transform 1 0 9108 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_99
timestamp 1618419204
transform 1 0 10212 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _317_
timestamp 1619507013
transform -1 0 11132 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1618419204
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_109
timestamp 1618419204
transform 1 0 11132 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1618419204
transform 1 0 11500 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_115
timestamp 1618419204
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1618419204
transform 1 0 13708 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[3\].id.delayenb1
timestamp 1618419204
transform 1 0 12880 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_17_127
timestamp 1618419204
transform 1 0 12788 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_133
timestamp 1618419204
transform 1 0 13340 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_140
timestamp 1618419204
transform 1 0 13984 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _373_
timestamp 1618419204
transform -1 0 16284 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1618419204
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_152
timestamp 1618419204
transform 1 0 15088 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_165
timestamp 1618419204
transform 1 0 16284 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_172
timestamp 1618419204
transform 1 0 16928 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1618419204
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1618419204
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1618419204
transform -1 0 21804 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1619507013
transform -1 0 20976 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_208
timestamp 1618419204
transform 1 0 20240 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_212
timestamp 1618419204
transform 1 0 20608 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_216
timestamp 1618419204
transform 1 0 20976 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1618419204
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1618419204
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1618419204
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1618419204
transform 1 0 4232 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1618419204
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1618419204
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_30
timestamp 1618419204
transform 1 0 3864 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_37
timestamp 1618419204
transform 1 0 4508 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_49
timestamp 1618419204
transform 1 0 5612 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _248_
timestamp 1618419204
transform 1 0 6072 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1619507013
transform 1 0 7176 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _310_
timestamp 1619507013
transform -1 0 8280 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_18_53
timestamp 1618419204
transform 1 0 5980 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_59
timestamp 1618419204
transform 1 0 6532 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_65
timestamp 1618419204
transform 1 0 7084 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_69
timestamp 1618419204
transform 1 0 7452 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 10856 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1618419204
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_78
timestamp 1618419204
transform 1 0 8280 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_87
timestamp 1618419204
transform 1 0 9108 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_95
timestamp 1618419204
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  _290_
timestamp 1618419204
transform 1 0 11500 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 12788 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_18_106
timestamp 1618419204
transform 1 0 10856 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_112
timestamp 1618419204
transform 1 0 11408 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_118
timestamp 1618419204
transform 1 0 11960 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1618419204
transform 1 0 14720 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1618419204
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_127
timestamp 1618419204
transform 1 0 12788 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_139
timestamp 1618419204
transform 1 0 13892 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_144
timestamp 1618419204
transform 1 0 14352 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_157
timestamp 1618419204
transform 1 0 15548 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_169
timestamp 1618419204
transform 1 0 16652 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _341_
timestamp 1618419204
transform 1 0 17296 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_175
timestamp 1618419204
transform 1 0 17204 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_179
timestamp 1618419204
transform 1 0 17572 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_191
timestamp 1618419204
transform 1 0 18676 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1618419204
transform 1 0 19964 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1618419204
transform -1 0 21804 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1618419204
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1618419204
transform 1 0 20700 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_199
timestamp 1618419204
transform 1 0 19412 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_201
timestamp 1618419204
transform 1 0 19596 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_208
timestamp 1618419204
transform 1 0 20240 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_212
timestamp 1618419204
transform 1 0 20608 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_216
timestamp 1618419204
transform 1 0 20976 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1618419204
transform 1 0 1380 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_7
timestamp 1618419204
transform 1 0 1748 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1618419204
transform -1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1618419204
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1618419204
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_15
timestamp 1618419204
transform 1 0 2484 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_9
timestamp 1618419204
transform 1 0 1932 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_15
timestamp 1618419204
transform 1 0 2484 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[7\].id.delayenb0
timestamp 1618419204
transform 1 0 2024 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_20_21
timestamp 1618419204
transform 1 0 3036 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_23
timestamp 1618419204
transform 1 0 3220 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  ringosc.dstage\[7\].id.delaybuf0
timestamp 1619507013
transform -1 0 3404 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[6\].id.delayenb0
timestamp 1618419204
transform 1 0 2760 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _305_
timestamp 1618419204
transform 1 0 5612 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _364_
timestamp 1618419204
transform 1 0 4232 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen0
timestamp 1618419204
transform 1 0 3588 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1618419204
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_32
timestamp 1618419204
transform 1 0 4048 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_44
timestamp 1618419204
transform 1 0 5152 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_25
timestamp 1618419204
transform 1 0 3404 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_30
timestamp 1618419204
transform 1 0 3864 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_43
timestamp 1618419204
transform 1 0 5060 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_56
timestamp 1618419204
transform 1 0 6256 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_58
timestamp 1618419204
transform 1 0 6440 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_56
timestamp 1618419204
transform 1 0 6256 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1618419204
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_66
timestamp 1618419204
transform 1 0 7176 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _293_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 7176 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _254_
timestamp 1618419204
transform 1 0 6808 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_20_73
timestamp 1618419204
transform 1 0 7820 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_69
timestamp 1618419204
transform 1 0 7452 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1619507013
transform 1 0 7544 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1619507013
transform -1 0 8464 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _294_
timestamp 1618419204
transform 1 0 8188 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _309_
timestamp 1618419204
transform 1 0 9384 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _320_
timestamp 1618419204
transform 1 0 9844 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1618419204
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_82
timestamp 1618419204
transform 1 0 8648 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_95
timestamp 1618419204
transform 1 0 9844 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_80
timestamp 1618419204
transform 1 0 8464 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_87
timestamp 1618419204
transform 1 0 9108 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 11224 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _371_
timestamp 1618419204
transform -1 0 12972 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1618419204
transform -1 0 12696 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1618419204
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_110
timestamp 1618419204
transform 1 0 11224 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_115
timestamp 1618419204
transform 1 0 11684 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1618419204
transform 1 0 12052 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_104
timestamp 1618419204
transform 1 0 10672 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_116
timestamp 1618419204
transform 1 0 11776 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _292_
timestamp 1618419204
transform 1 0 13340 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1618419204
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_129
timestamp 1618419204
transform 1 0 12972 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_138
timestamp 1618419204
transform 1 0 13800 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_126
timestamp 1618419204
transform 1 0 12696 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_138
timestamp 1618419204
transform 1 0 13800 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_142
timestamp 1618419204
transform 1 0 14168 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_144
timestamp 1618419204
transform 1 0 14352 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_160
timestamp 1618419204
transform 1 0 15824 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_153
timestamp 1618419204
transform 1 0 15180 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1618419204
transform 1 0 15548 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _207_
timestamp 1619507013
transform -1 0 15180 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_170
timestamp 1618419204
transform 1 0 16744 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_162
timestamp 1618419204
transform 1 0 16008 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1618419204
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_172
timestamp 1618419204
transform 1 0 16928 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_150
timestamp 1618419204
transform 1 0 14904 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _386_
timestamp 1619507013
transform -1 0 18308 0 -1 13600
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _385_
timestamp 1619507013
transform 1 0 18216 0 1 12512
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1618419204
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_187
timestamp 1618419204
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_199
timestamp 1618419204
transform 1 0 19412 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_209
timestamp 1618419204
transform 1 0 20332 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1618419204
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_221
timestamp 1618419204
transform 1 0 21436 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_213
timestamp 1618419204
transform 1 0 20700 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_218
timestamp 1618419204
transform 1 0 21160 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1618419204
transform 1 0 20884 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1618419204
transform -1 0 21804 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1618419204
transform -1 0 21804 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_201
timestamp 1618419204
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1618419204
transform 1 0 1932 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen1
timestamp 1618419204
transform 1 0 3128 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1618419204
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1618419204
transform 1 0 1380 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_18
timestamp 1618419204
transform 1 0 2760 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1618419204
transform 1 0 3956 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1618419204
transform 1 0 3588 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_34
timestamp 1618419204
transform 1 0 4232 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_46
timestamp 1618419204
transform 1 0 5336 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1618419204
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_54
timestamp 1618419204
transform 1 0 6072 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1618419204
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_70
timestamp 1618419204
transform 1 0 7544 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1619507013
transform -1 0 8740 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1618419204
transform 1 0 9476 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_78
timestamp 1618419204
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_83
timestamp 1618419204
transform 1 0 8740 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1618419204
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_100
timestamp 1618419204
transform 1 0 10304 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_112
timestamp 1618419204
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_115
timestamp 1618419204
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _401_
timestamp 1619507013
transform 1 0 13984 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1618419204
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_139
timestamp 1618419204
transform 1 0 13892 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1618419204
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1618419204
transform 1 0 15824 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_168
timestamp 1618419204
transform 1 0 16560 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_172
timestamp 1618419204
transform 1 0 16928 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _285_
timestamp 1618419204
transform -1 0 17664 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _288_
timestamp 1618419204
transform 1 0 18032 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_21_180
timestamp 1618419204
transform 1 0 17664 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_189
timestamp 1618419204
transform 1 0 18492 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_197
timestamp 1618419204
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _200_
timestamp 1619507013
transform -1 0 20056 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1618419204
transform 1 0 20700 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1618419204
transform -1 0 21804 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_206
timestamp 1618419204
transform 1 0 20056 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_212
timestamp 1618419204
transform 1 0 20608 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_216
timestamp 1618419204
transform 1 0 20976 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen0
timestamp 1618419204
transform 1 0 1932 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_1  ringosc.dstage\[7\].id.delayenb1
timestamp 1618419204
transform -1 0 3220 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1618419204
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1618419204
transform 1 0 1380 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_14
timestamp 1618419204
transform 1 0 2392 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_23
timestamp 1618419204
transform 1 0 3220 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1618419204
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1618419204
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_42
timestamp 1618419204
transform 1 0 4968 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _251_
timestamp 1619507013
transform -1 0 6808 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1619507013
transform -1 0 7452 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_54
timestamp 1618419204
transform 1 0 6072 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_62
timestamp 1618419204
transform 1 0 6808 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_69
timestamp 1618419204
transform 1 0 7452 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1619507013
transform 1 0 9844 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1619507013
transform 1 0 8372 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1618419204
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_77
timestamp 1618419204
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_82
timestamp 1618419204
transform 1 0 8648 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_87
timestamp 1618419204
transform 1 0 9108 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_98
timestamp 1618419204
transform 1 0 10120 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1619507013
transform 1 0 10488 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _395_
timestamp 1619507013
transform 1 0 11132 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_22_105
timestamp 1618419204
transform 1 0 10764 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _199_
timestamp 1619507013
transform -1 0 15364 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1618419204
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_130
timestamp 1618419204
transform 1 0 13064 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_142
timestamp 1618419204
transform 1 0 14168 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_144
timestamp 1618419204
transform 1 0 14352 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1619507013
transform 1 0 16192 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _286_
timestamp 1618419204
transform -1 0 17480 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_22_155
timestamp 1618419204
transform 1 0 15364 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_163
timestamp 1618419204
transform 1 0 16100 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1618419204
transform 1 0 16468 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 18676 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_178
timestamp 1618419204
transform 1 0 17480 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_191
timestamp 1618419204
transform 1 0 18676 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 19964 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1618419204
transform -1 0 21804 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1618419204
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_199
timestamp 1618419204
transform 1 0 19412 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_201
timestamp 1618419204
transform 1 0 19596 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_213
timestamp 1618419204
transform 1 0 20700 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_221
timestamp 1618419204
transform 1 0 21436 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1618419204
transform -1 0 2852 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1618419204
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1618419204
transform -1 0 2116 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1618419204
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1618419204
transform 1 0 1748 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_11
timestamp 1618419204
transform 1 0 2116 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_15
timestamp 1618419204
transform 1 0 2484 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_19
timestamp 1618419204
transform 1 0 2852 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _262_
timestamp 1618419204
transform -1 0 5980 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _267_
timestamp 1618419204
transform 1 0 4876 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_31
timestamp 1618419204
transform 1 0 3956 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_39
timestamp 1618419204
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_44
timestamp 1618419204
transform 1 0 5152 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _252_
timestamp 1619507013
transform 1 0 7912 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _256_
timestamp 1619507013
transform -1 0 7544 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1618419204
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_53
timestamp 1618419204
transform 1 0 5980 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_58
timestamp 1618419204
transform 1 0 6440 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_70
timestamp 1618419204
transform 1 0 7544 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _258_
timestamp 1619507013
transform 1 0 8924 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _261_
timestamp 1618419204
transform -1 0 10304 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_81
timestamp 1618419204
transform 1 0 8556 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_92
timestamp 1618419204
transform 1 0 9568 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1618419204
transform 1 0 12328 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1618419204
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_100
timestamp 1618419204
transform 1 0 10304 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_112
timestamp 1618419204
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_115
timestamp 1618419204
transform 1 0 11684 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1618419204
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _212_
timestamp 1618419204
transform 1 0 14352 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1618419204
transform 1 0 12604 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_137
timestamp 1618419204
transform 1 0 13708 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_143
timestamp 1618419204
transform 1 0 14260 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1619507013
transform -1 0 16468 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _223_
timestamp 1619507013
transform 1 0 15456 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1618419204
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_152
timestamp 1618419204
transform 1 0 15088 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_160
timestamp 1618419204
transform 1 0 15824 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_167
timestamp 1618419204
transform 1 0 16468 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_172
timestamp 1618419204
transform 1 0 16928 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _210_
timestamp 1619507013
transform -1 0 18952 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _279_
timestamp 1618419204
transform -1 0 17756 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _400_
timestamp 1619507013
transform 1 0 19320 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_23_181
timestamp 1618419204
transform 1 0 17756 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_194
timestamp 1618419204
transform 1 0 18952 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1618419204
transform -1 0 21804 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_218
timestamp 1618419204
transform 1 0 21160 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1618419204
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1618419204
transform -1 0 1656 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_6
timestamp 1618419204
transform 1 0 1656 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_18
timestamp 1618419204
transform 1 0 2760 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 5060 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1618419204
transform 1 0 4416 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1618419204
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_26
timestamp 1618419204
transform 1 0 3496 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_30
timestamp 1618419204
transform 1 0 3864 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_39
timestamp 1618419204
transform 1 0 4692 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 7912 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1619507013
transform -1 0 6440 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _265_
timestamp 1618419204
transform 1 0 6808 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_51
timestamp 1618419204
transform 1 0 5796 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_58
timestamp 1618419204
transform 1 0 6440 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_70
timestamp 1618419204
transform 1 0 7544 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _394_
timestamp 1619507013
transform 1 0 9476 0 -1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1618419204
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_82
timestamp 1618419204
transform 1 0 8648 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_87
timestamp 1618419204
transform 1 0 9108 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_112
timestamp 1618419204
transform 1 0 11408 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_124
timestamp 1618419204
transform 1 0 12512 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_1  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 14720 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1618419204
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_136
timestamp 1618419204
transform 1 0 13616 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_142
timestamp 1618419204
transform 1 0 14168 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_144
timestamp 1618419204
transform 1 0 14352 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1619507013
transform -1 0 17112 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_156
timestamp 1618419204
transform 1 0 15456 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_168
timestamp 1618419204
transform 1 0 16560 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1619507013
transform -1 0 18400 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_174
timestamp 1618419204
transform 1 0 17112 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_182
timestamp 1618419204
transform 1 0 17848 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_188
timestamp 1618419204
transform 1 0 18400 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1618419204
transform -1 0 21804 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1618419204
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1618419204
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_201
timestamp 1618419204
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_213
timestamp 1618419204
transform 1 0 20700 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_218
timestamp 1618419204
transform 1 0 21160 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1619507013
transform 1 0 2576 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _393_
timestamp 1619507013
transform 1 0 3312 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1618419204
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1618419204
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 1618419204
transform 1 0 2484 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_19
timestamp 1618419204
transform 1 0 2852 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_23
timestamp 1618419204
transform 1 0 3220 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_45
timestamp 1618419204
transform 1 0 5244 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _263_
timestamp 1618419204
transform -1 0 7176 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1618419204
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_58
timestamp 1618419204
transform 1 0 6440 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_66
timestamp 1618419204
transform 1 0 7176 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _266_
timestamp 1618419204
transform -1 0 9108 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_78
timestamp 1618419204
transform 1 0 8280 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_82
timestamp 1618419204
transform 1 0 8648 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_87
timestamp 1618419204
transform 1 0 9108 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_99
timestamp 1618419204
transform 1 0 10212 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp 1618419204
transform -1 0 10764 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1618419204
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_105
timestamp 1618419204
transform 1 0 10764 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1618419204
transform 1 0 11500 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1618419204
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _219_
timestamp 1618419204
transform 1 0 13892 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _220_
timestamp 1618419204
transform 1 0 12788 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1618419204
transform 1 0 13524 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_145
timestamp 1618419204
transform 1 0 14444 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1618419204
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_157
timestamp 1618419204
transform 1 0 15548 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1618419204
transform 1 0 16652 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_172
timestamp 1618419204
transform 1 0 16928 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2ai_1  _228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 19596 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 17296 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_25_183
timestamp 1618419204
transform 1 0 17940 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_191
timestamp 1618419204
transform 1 0 18676 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1618419204
transform -1 0 21804 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1618419204
transform 1 0 20700 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_201
timestamp 1618419204
transform 1 0 19596 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_216
timestamp 1618419204
transform 1 0 20976 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1618419204
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1618419204
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1618419204
transform -1 0 2576 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1618419204
transform -1 0 1932 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1618419204
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_9
timestamp 1618419204
transform 1 0 1932 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_16
timestamp 1618419204
transform 1 0 2576 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1618419204
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1618419204
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1618419204
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_28
timestamp 1618419204
transform 1 0 3680 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1618419204
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_42
timestamp 1618419204
transform 1 0 4968 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1618419204
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_39
timestamp 1618419204
transform 1 0 4692 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_47
timestamp 1618419204
transform 1 0 5428 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_58
timestamp 1618419204
transform 1 0 6440 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_53
timestamp 1618419204
transform 1 0 5980 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1618419204
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_1  _250_
timestamp 1619507013
transform 1 0 6808 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1619507013
transform -1 0 5980 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_70
timestamp 1618419204
transform 1 0 7544 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_66
timestamp 1618419204
transform 1 0 7176 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _270_
timestamp 1618419204
transform -1 0 8280 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1619507013
transform 1 0 7268 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_70
timestamp 1618419204
transform 1 0 7544 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_54
timestamp 1618419204
transform 1 0 6072 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1619507013
transform 1 0 8648 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1618419204
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_82
timestamp 1618419204
transform 1 0 8648 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1618419204
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_99
timestamp 1618419204
transform 1 0 10212 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_78
timestamp 1618419204
transform 1 0 8280 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_85
timestamp 1618419204
transform 1 0 8924 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_97
timestamp 1618419204
transform 1 0 10028 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _221_
timestamp 1618419204
transform -1 0 12512 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 11408 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1618419204
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_111
timestamp 1618419204
transform 1 0 11316 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_120
timestamp 1618419204
transform 1 0 12144 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_109
timestamp 1618419204
transform 1 0 11132 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1618419204
transform 1 0 11500 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_115
timestamp 1618419204
transform 1 0 11684 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_124
timestamp 1618419204
transform 1 0 12512 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _198_
timestamp 1619507013
transform 1 0 14720 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _206_
timestamp 1619507013
transform -1 0 13892 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _402_
timestamp 1619507013
transform -1 0 15548 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1618419204
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_132
timestamp 1618419204
transform 1 0 13248 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_139
timestamp 1618419204
transform 1 0 13892 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_144
timestamp 1618419204
transform 1 0 14352 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_136
timestamp 1618419204
transform 1 0 13616 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _384_
timestamp 1619507013
transform 1 0 16284 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1618419204
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_155
timestamp 1618419204
transform 1 0 15364 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_163
timestamp 1618419204
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_157
timestamp 1618419204
transform 1 0 15548 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1618419204
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_172
timestamp 1618419204
transform 1 0 16928 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1619507013
transform 1 0 18860 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _227_
timestamp 1618419204
transform -1 0 18952 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _289_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 17296 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _399_
timestamp 1619507013
transform 1 0 19320 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_26_185
timestamp 1618419204
transform 1 0 18124 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_196
timestamp 1618419204
transform 1 0 19136 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_184
timestamp 1618419204
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_194
timestamp 1618419204
transform 1 0 18952 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_201
timestamp 1618419204
transform 1 0 19596 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1618419204
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1618419204
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _208_
timestamp 1619507013
transform 1 0 19964 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1618419204
transform 1 0 20792 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_218
timestamp 1618419204
transform 1 0 21160 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_221
timestamp 1618419204
transform 1 0 21436 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_217
timestamp 1618419204
transform 1 0 21068 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1618419204
transform -1 0 21804 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1618419204
transform -1 0 21804 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1618419204
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1618419204
transform -1 0 1656 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_6
timestamp 1618419204
transform 1 0 1656 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_18
timestamp 1618419204
transform 1 0 2760 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _391_
timestamp 1619507013
transform 1 0 4232 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1618419204
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_26
timestamp 1618419204
transform 1 0 3496 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_30
timestamp 1618419204
transform 1 0 3864 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _244_
timestamp 1619507013
transform 1 0 6532 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _272_
timestamp 1618419204
transform 1 0 7636 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_55
timestamp 1618419204
transform 1 0 6164 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_66
timestamp 1618419204
transform 1 0 7176 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_70
timestamp 1618419204
transform 1 0 7544 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _392_
timestamp 1619507013
transform 1 0 9476 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1618419204
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_79
timestamp 1618419204
transform 1 0 8372 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 1618419204
transform 1 0 8924 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_87
timestamp 1618419204
transform 1 0 9108 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_2  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 12880 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_112
timestamp 1618419204
transform 1 0 11408 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _213_
timestamp 1618419204
transform -1 0 15456 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1618419204
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_128
timestamp 1618419204
transform 1 0 12880 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_140
timestamp 1618419204
transform 1 0 13984 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_144
timestamp 1618419204
transform 1 0 14352 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_156
timestamp 1618419204
transform 1 0 15456 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_168
timestamp 1618419204
transform 1 0 16560 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1619507013
transform -1 0 19136 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _343_
timestamp 1618419204
transform 1 0 17388 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_176
timestamp 1618419204
transform 1 0 17296 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1618419204
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_192
timestamp 1618419204
transform 1 0 18768 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_196
timestamp 1618419204
transform 1 0 19136 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _201_
timestamp 1619507013
transform 1 0 19964 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1618419204
transform -1 0 21804 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1618419204
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_201
timestamp 1618419204
transform 1 0 19596 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_212
timestamp 1618419204
transform 1 0 20608 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_220
timestamp 1618419204
transform 1 0 21344 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1618419204
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1618419204
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1618419204
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_1  _275_
timestamp 1618419204
transform 1 0 5152 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1618419204
transform -1 0 4784 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_27
timestamp 1618419204
transform 1 0 3588 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_35
timestamp 1618419204
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_40
timestamp 1618419204
transform 1 0 4784 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _246_
timestamp 1619507013
transform 1 0 7820 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _269_
timestamp 1618419204
transform 1 0 6808 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1618419204
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1618419204
transform 1 0 5888 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_56
timestamp 1618419204
transform 1 0 6256 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_58
timestamp 1618419204
transform 1 0 6440 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_67
timestamp 1618419204
transform 1 0 7268 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _273_
timestamp 1618419204
transform -1 0 9200 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1618419204
transform -1 0 10120 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_80
timestamp 1618419204
transform 1 0 8464 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_88
timestamp 1618419204
transform 1 0 9200 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_94
timestamp 1618419204
transform 1 0 9752 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_98
timestamp 1618419204
transform 1 0 10120 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1619507013
transform 1 0 10948 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _237_
timestamp 1618419204
transform 1 0 12052 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1618419204
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_106
timestamp 1618419204
transform 1 0 10856 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_110
timestamp 1618419204
transform 1 0 11224 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_115
timestamp 1618419204
transform 1 0 11684 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_124
timestamp 1618419204
transform 1 0 12512 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _218_
timestamp 1618419204
transform 1 0 13708 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1619507013
transform -1 0 13156 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_131
timestamp 1618419204
transform 1 0 13156 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_140
timestamp 1618419204
transform 1 0 13984 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1618419204
transform -1 0 16468 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1618419204
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_152
timestamp 1618419204
transform 1 0 15088 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_167
timestamp 1618419204
transform 1 0 16468 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_172
timestamp 1618419204
transform 1 0 16928 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1619507013
transform -1 0 18400 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _231_
timestamp 1618419204
transform -1 0 19596 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp 1618419204
transform 1 0 17296 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_179
timestamp 1618419204
transform 1 0 17572 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_188
timestamp 1618419204
transform 1 0 18400 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1618419204
transform -1 0 21804 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1618419204
transform 1 0 20884 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_201
timestamp 1618419204
transform 1 0 19596 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_213
timestamp 1618419204
transform 1 0 20700 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_218
timestamp 1618419204
transform 1 0 21160 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1618419204
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1618419204
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1618419204
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _274_
timestamp 1618419204
transform -1 0 6072 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1618419204
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1618419204
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_30
timestamp 1618419204
transform 1 0 3864 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_42
timestamp 1618419204
transform 1 0 4968 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_48
timestamp 1618419204
transform 1 0 5520 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1619507013
transform 1 0 6440 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1619507013
transform 1 0 7820 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1619507013
transform -1 0 7452 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_54
timestamp 1618419204
transform 1 0 6072 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_61
timestamp 1618419204
transform 1 0 6716 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_65
timestamp 1618419204
transform 1 0 7084 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_69
timestamp 1618419204
transform 1 0 7452 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1618419204
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_76
timestamp 1618419204
transform 1 0 8096 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_84
timestamp 1618419204
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_87
timestamp 1618419204
transform 1 0 9108 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_99
timestamp 1618419204
transform 1 0 10212 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_4  _238_
timestamp 1619507013
transform 1 0 11132 0 -1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_30_107
timestamp 1618419204
transform 1 0 10948 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  _214_
timestamp 1618419204
transform -1 0 13892 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1618419204
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_126
timestamp 1618419204
transform 1 0 12696 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_139
timestamp 1618419204
transform 1 0 13892 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_144
timestamp 1618419204
transform 1 0 14352 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _387_
timestamp 1619507013
transform 1 0 15916 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_30_156
timestamp 1618419204
transform 1 0 15456 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_160
timestamp 1618419204
transform 1 0 15824 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a21boi_1  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 18584 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_182
timestamp 1618419204
transform 1 0 17848 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_196
timestamp 1618419204
transform 1 0 19136 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1618419204
transform -1 0 21804 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1618419204
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_201
timestamp 1618419204
transform 1 0 19596 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_213
timestamp 1618419204
transform 1 0 20700 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_221
timestamp 1618419204
transform 1 0 21436 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1618419204
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1619507013
transform 1 0 2392 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1618419204
transform 1 0 1380 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_11
timestamp 1618419204
transform 1 0 2116 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_17
timestamp 1618419204
transform 1 0 2668 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _338_
timestamp 1618419204
transform 1 0 4416 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_29
timestamp 1618419204
transform 1 0 3772 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_35
timestamp 1618419204
transform 1 0 4324 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_39
timestamp 1618419204
transform 1 0 4692 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_47
timestamp 1618419204
transform 1 0 5428 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1619507013
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1619507013
transform 1 0 7728 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _241_
timestamp 1618419204
transform -1 0 5980 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1618419204
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_53
timestamp 1618419204
transform 1 0 5980 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_58
timestamp 1618419204
transform 1 0 6440 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_65
timestamp 1618419204
transform 1 0 7084 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_71
timestamp 1618419204
transform 1 0 7636 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_75
timestamp 1618419204
transform 1 0 8004 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_87
timestamp 1618419204
transform 1 0 9108 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_99
timestamp 1618419204
transform 1 0 10212 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__a41o_2  _234_
timestamp 1619507013
transform 1 0 12052 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1618419204
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_111
timestamp 1618419204
transform 1 0 11316 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_115
timestamp 1618419204
transform 1 0 11684 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _216_
timestamp 1618419204
transform 1 0 13800 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_31_128
timestamp 1618419204
transform 1 0 12880 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_136
timestamp 1618419204
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_147
timestamp 1618419204
transform 1 0 14628 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1619507013
transform 1 0 14996 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _283_
timestamp 1618419204
transform 1 0 15640 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1618419204
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_154
timestamp 1618419204
transform 1 0 15272 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_167
timestamp 1618419204
transform 1 0 16468 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_172
timestamp 1618419204
transform 1 0 16928 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_4  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 18400 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _236_
timestamp 1618419204
transform -1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_184
timestamp 1618419204
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_195
timestamp 1618419204
transform 1 0 19044 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _229_
timestamp 1618419204
transform 1 0 19412 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1618419204
transform -1 0 21804 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_202
timestamp 1618419204
transform 1 0 19688 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_214
timestamp 1618419204
transform 1 0 20792 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1618419204
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1618419204
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1618419204
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _278_
timestamp 1619507013
transform 1 0 4784 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1618419204
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1618419204
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_30
timestamp 1618419204
transform 1 0 3864 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_38
timestamp 1618419204
transform 1 0 4600 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_47
timestamp 1618419204
transform 1 0 5428 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _240_
timestamp 1619507013
transform 1 0 6164 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _276_
timestamp 1618419204
transform 1 0 7176 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_32_62
timestamp 1618419204
transform 1 0 6808 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_71
timestamp 1618419204
transform 1 0 7636 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1619507013
transform 1 0 8004 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1618419204
transform 1 0 9476 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1618419204
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_78
timestamp 1618419204
transform 1 0 8280 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_87
timestamp 1618419204
transform 1 0 9108 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1618419204
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1619507013
transform -1 0 11960 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_106
timestamp 1618419204
transform 1 0 10856 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_114
timestamp 1618419204
transform 1 0 11592 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_118
timestamp 1618419204
transform 1 0 11960 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _205_
timestamp 1619507013
transform -1 0 15364 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _215_
timestamp 1618419204
transform 1 0 13156 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1618419204
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_130
timestamp 1618419204
transform 1 0 13064 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_139
timestamp 1618419204
transform 1 0 13892 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_144
timestamp 1618419204
transform 1 0 14352 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _282_
timestamp 1619507013
transform 1 0 15732 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_155
timestamp 1618419204
transform 1 0 15364 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_163
timestamp 1618419204
transform 1 0 16100 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_175
timestamp 1618419204
transform 1 0 17204 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1618419204
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp 1618419204
transform 1 0 20608 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1618419204
transform -1 0 21804 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1618419204
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_199
timestamp 1618419204
transform 1 0 19412 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_201
timestamp 1618419204
transform 1 0 19596 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_209
timestamp 1618419204
transform 1 0 20332 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_215
timestamp 1618419204
transform 1 0 20884 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_221
timestamp 1618419204
transform 1 0 21436 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _389_
timestamp 1619507013
transform 1 0 3220 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1618419204
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1618419204
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1618419204
transform -1 0 1656 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_6
timestamp 1618419204
transform 1 0 1656 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_18
timestamp 1618419204
transform 1 0 2760 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_22
timestamp 1618419204
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1618419204
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1618419204
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1619507013
transform -1 0 5704 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1618419204
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_43
timestamp 1618419204
transform 1 0 5060 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1618419204
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_30
timestamp 1618419204
transform 1 0 3864 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_42
timestamp 1618419204
transform 1 0 4968 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_50
timestamp 1618419204
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_58
timestamp 1618419204
transform 1 0 6440 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_56
timestamp 1618419204
transform 1 0 6256 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_50
timestamp 1618419204
transform 1 0 5704 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1618419204
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_1  _277_
timestamp 1618419204
transform 1 0 5796 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _242_
timestamp 1618419204
transform -1 0 7176 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_71
timestamp 1618419204
transform 1 0 7636 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_59
timestamp 1618419204
transform 1 0 6532 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_66
timestamp 1618419204
transform 1 0 7176 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _398_
timestamp 1619507013
transform 1 0 8372 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1618419204
transform 1 0 9016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1619507013
transform 1 0 8188 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_78
timestamp 1618419204
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_99
timestamp 1618419204
transform 1 0 10212 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_80
timestamp 1618419204
transform 1 0 8464 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_87
timestamp 1618419204
transform 1 0 9108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_99
timestamp 1618419204
transform 1 0 10212 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _202_
timestamp 1619507013
transform -1 0 11224 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 10580 0 -1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1618419204
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_110
timestamp 1618419204
transform 1 0 11224 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_115
timestamp 1618419204
transform 1 0 11684 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_113
timestamp 1618419204
transform 1 0 11500 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _195_
timestamp 1619507013
transform -1 0 14628 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1618419204
transform 1 0 14260 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_127
timestamp 1618419204
transform 1 0 12788 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_139
timestamp 1618419204
transform 1 0 13892 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_147
timestamp 1618419204
transform 1 0 14628 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_125
timestamp 1618419204
transform 1 0 12604 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_137
timestamp 1618419204
transform 1 0 13708 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_144
timestamp 1618419204
transform 1 0 14352 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1619507013
transform 1 0 14996 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _388_
timestamp 1619507013
transform 1 0 15180 0 -1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1618419204
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_154
timestamp 1618419204
transform 1 0 15272 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_166
timestamp 1618419204
transform 1 0 16376 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_170
timestamp 1618419204
transform 1 0 16744 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_172
timestamp 1618419204
transform 1 0 16928 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 1618419204
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _339_
timestamp 1618419204
transform 1 0 17480 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp 1618419204
transform 1 0 18124 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _383_
timestamp 1619507013
transform 1 0 19320 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1618419204
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_196
timestamp 1618419204
transform 1 0 19136 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_174
timestamp 1618419204
transform 1 0 17112 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_181
timestamp 1618419204
transform 1 0 17756 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_188
timestamp 1618419204
transform 1 0 18400 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1618419204
transform -1 0 21804 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1618419204
transform -1 0 21804 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1618419204
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1618419204
transform 1 0 19964 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1618419204
transform 1 0 20792 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1618419204
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_201
timestamp 1618419204
transform 1 0 19596 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_208
timestamp 1618419204
transform 1 0 20240 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_218
timestamp 1618419204
transform 1 0 21160 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _349_
timestamp 1618419204
transform 1 0 2484 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1618419204
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output44
timestamp 1618419204
transform 1 0 1748 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1618419204
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_10
timestamp 1618419204
transform 1 0 2024 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_14
timestamp 1618419204
transform 1 0 2392 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_18
timestamp 1618419204
transform 1 0 2760 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_24
timestamp 1618419204
transform 1 0 3312 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1619507013
transform 1 0 3404 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1619507013
transform 1 0 5060 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_28
timestamp 1618419204
transform 1 0 3680 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_40
timestamp 1618419204
transform 1 0 4784 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_46
timestamp 1618419204
transform 1 0 5336 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1618419204
transform 1 0 6808 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _396_
timestamp 1619507013
transform 1 0 7452 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1618419204
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1619507013
transform 1 0 5704 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_53
timestamp 1618419204
transform 1 0 5980 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_58
timestamp 1618419204
transform 1 0 6440 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_65
timestamp 1618419204
transform 1 0 7084 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _204_
timestamp 1618419204
transform -1 0 10120 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_35_89
timestamp 1618419204
transform 1 0 9292 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_98
timestamp 1618419204
transform 1 0 10120 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _203_
timestamp 1619507013
transform 1 0 10488 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1618419204
transform 1 0 12052 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1618419204
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_109
timestamp 1618419204
transform 1 0 11132 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 1618419204
transform 1 0 11500 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_115
timestamp 1618419204
transform 1 0 11684 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_122
timestamp 1618419204
transform 1 0 12328 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _403_
timestamp 1619507013
transform 1 0 12972 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_35_128
timestamp 1618419204
transform 1 0 12880 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_149
timestamp 1618419204
transform 1 0 14812 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1618419204
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1618419204
transform 1 0 15180 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1618419204
transform 1 0 15824 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_156
timestamp 1618419204
transform 1 0 15456 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_163
timestamp 1618419204
transform 1 0 16100 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_172
timestamp 1618419204
transform 1 0 16928 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _381_
timestamp 1619507013
transform -1 0 19136 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_35_196
timestamp 1618419204
transform 1 0 19136 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_4  _193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 21160 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1618419204
transform -1 0 21804 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_218
timestamp 1618419204
transform 1 0 21160 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1618419204
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1618419204
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1618419204
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _390_
timestamp 1619507013
transform 1 0 5152 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1618419204
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1618419204
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_30
timestamp 1618419204
transform 1 0 3864 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_42
timestamp 1618419204
transform 1 0 4968 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_64
timestamp 1618419204
transform 1 0 6992 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 1618419204
transform -1 0 8648 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1618419204
transform 1 0 9016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1619507013
transform 1 0 9476 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_76
timestamp 1618419204
transform 1 0 8096 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_82
timestamp 1618419204
transform 1 0 8648 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_87
timestamp 1618419204
transform 1 0 9108 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_94
timestamp 1618419204
transform 1 0 9752 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _397_
timestamp 1619507013
transform 1 0 10672 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_36_102
timestamp 1618419204
transform 1 0 10488 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_124
timestamp 1618419204
transform 1 0 12512 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp 1618419204
transform 1 0 14720 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1618419204
transform 1 0 14260 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1619507013
transform 1 0 13064 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_133
timestamp 1618419204
transform 1 0 13340 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1618419204
transform 1 0 14076 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_144
timestamp 1618419204
transform 1 0 14352 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1618419204
transform -1 0 16928 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_151
timestamp 1618419204
transform 1 0 14996 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_163
timestamp 1618419204
transform 1 0 16100 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_172
timestamp 1618419204
transform 1 0 16928 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _382_
timestamp 1619507013
transform 1 0 17296 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_36_196
timestamp 1618419204
transform 1 0 19136 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _345_
timestamp 1618419204
transform 1 0 19964 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1618419204
transform -1 0 21804 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1618419204
transform 1 0 19504 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input75
timestamp 1619507013
transform -1 0 21160 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_201
timestamp 1618419204
transform 1 0 19596 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_208
timestamp 1618419204
transform 1 0 20240 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_214
timestamp 1618419204
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_218
timestamp 1618419204
transform 1 0 21160 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1618419204
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1618419204
transform -1 0 3036 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1618419204
transform 1 0 2116 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1618419204
transform -1 0 1748 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_7
timestamp 1618419204
transform 1 0 1748 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_14
timestamp 1618419204
transform 1 0 2392 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_21
timestamp 1618419204
transform 1 0 3036 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1618419204
transform 1 0 3772 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1618419204
transform -1 0 4876 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_30
timestamp 1618419204
transform 1 0 3864 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_41
timestamp 1618419204
transform 1 0 4876 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_49
timestamp 1618419204
transform 1 0 5612 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1618419204
transform 1 0 6440 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1618419204
transform -1 0 8096 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1618419204
transform 1 0 5796 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_54
timestamp 1618419204
transform 1 0 6072 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_59
timestamp 1618419204
transform 1 0 6532 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_71
timestamp 1618419204
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1618419204
transform 1 0 9108 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1618419204
transform 1 0 9660 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_76
timestamp 1618419204
transform 1 0 8096 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_84
timestamp 1618419204
transform 1 0 8832 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_88
timestamp 1618419204
transform 1 0 9200 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_92
timestamp 1618419204
transform 1 0 9568 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_96
timestamp 1618419204
transform 1 0 9936 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1618419204
transform 1 0 11776 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1618419204
transform 1 0 10672 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1618419204
transform 1 0 12236 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_107
timestamp 1618419204
transform 1 0 10948 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_115
timestamp 1618419204
transform 1 0 11684 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_117
timestamp 1618419204
transform 1 0 11868 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_124
timestamp 1618419204
transform 1 0 12512 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1618419204
transform 1 0 14444 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1618419204
transform -1 0 13156 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_131
timestamp 1618419204
transform 1 0 13156 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_143
timestamp 1618419204
transform 1 0 14260 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_146
timestamp 1618419204
transform 1 0 14536 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1618419204
transform -1 0 15180 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1618419204
transform 1 0 16468 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_153
timestamp 1618419204
transform 1 0 15180 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_165
timestamp 1618419204
transform 1 0 16284 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_170
timestamp 1618419204
transform 1 0 16744 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1618419204
transform 1 0 17112 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1618419204
transform 1 0 17940 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_175
timestamp 1618419204
transform 1 0 17204 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_186
timestamp 1618419204
transform 1 0 18216 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_198
timestamp 1618419204
transform 1 0 19320 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1618419204
transform -1 0 21804 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1618419204
transform 1 0 19780 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1618419204
transform 1 0 20240 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1619507013
transform -1 0 21160 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_202
timestamp 1618419204
transform 1 0 19688 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_204
timestamp 1618419204
transform 1 0 19872 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_211
timestamp 1618419204
transform 1 0 20516 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_218
timestamp 1618419204
transform 1 0 21160 0 1 22304
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 10208 800 10328 6 clockc
port 0 nsew signal tristate
rlabel metal3 s 0 12928 800 13048 6 clockd[0]
port 1 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 clockd[1]
port 2 nsew signal tristate
rlabel metal3 s 22179 20408 22979 20528 6 clockd[2]
port 3 nsew signal tristate
rlabel metal2 s 20718 0 20774 800 6 clockd[3]
port 4 nsew signal tristate
rlabel metal3 s 0 23128 800 23248 6 clockp[0]
port 5 nsew signal tristate
rlabel metal2 s 1858 0 1914 800 6 clockp[1]
port 6 nsew signal tristate
rlabel metal2 s 15658 0 15714 800 6 dco
port 7 nsew signal input
rlabel metal3 s 22179 15648 22979 15768 6 div[0]
port 8 nsew signal input
rlabel metal2 s 19798 24323 19854 25123 6 div[1]
port 9 nsew signal input
rlabel metal2 s 7838 24323 7894 25123 6 div[2]
port 10 nsew signal input
rlabel metal2 s 478 0 534 800 6 div[3]
port 11 nsew signal input
rlabel metal2 s 14738 24323 14794 25123 6 div[4]
port 12 nsew signal input
rlabel metal2 s 16578 24323 16634 25123 6 ext_trim[0]
port 13 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 ext_trim[10]
port 14 nsew signal input
rlabel metal2 s 2778 24323 2834 25123 6 ext_trim[11]
port 15 nsew signal input
rlabel metal3 s 22179 5448 22979 5568 6 ext_trim[12]
port 16 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 ext_trim[13]
port 17 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 ext_trim[14]
port 18 nsew signal input
rlabel metal3 s 22179 17688 22979 17808 6 ext_trim[15]
port 19 nsew signal input
rlabel metal2 s 4618 24323 4674 25123 6 ext_trim[16]
port 20 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 ext_trim[17]
port 21 nsew signal input
rlabel metal2 s 5998 24323 6054 25123 6 ext_trim[18]
port 22 nsew signal input
rlabel metal3 s 22179 10208 22979 10328 6 ext_trim[19]
port 23 nsew signal input
rlabel metal2 s 12898 24323 12954 25123 6 ext_trim[1]
port 24 nsew signal input
rlabel metal2 s 11518 24323 11574 25123 6 ext_trim[20]
port 25 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 ext_trim[21]
port 26 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 ext_trim[22]
port 27 nsew signal input
rlabel metal3 s 22179 23128 22979 23248 6 ext_trim[23]
port 28 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 ext_trim[24]
port 29 nsew signal input
rlabel metal2 s 9678 24323 9734 25123 6 ext_trim[25]
port 30 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 ext_trim[2]
port 31 nsew signal input
rlabel metal3 s 22179 8168 22979 8288 6 ext_trim[3]
port 32 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 ext_trim[4]
port 33 nsew signal input
rlabel metal3 s 22179 12928 22979 13048 6 ext_trim[5]
port 34 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 ext_trim[6]
port 35 nsew signal input
rlabel metal2 s 938 24323 994 25123 6 ext_trim[7]
port 36 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 ext_trim[8]
port 37 nsew signal input
rlabel metal3 s 22179 2728 22979 2848 6 ext_trim[9]
port 38 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 extclk_sel
port 39 nsew signal input
rlabel metal2 s 17958 24323 18014 25123 6 osc
port 40 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 reset
port 41 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 sel[0]
port 42 nsew signal input
rlabel metal2 s 21638 24323 21694 25123 6 sel[1]
port 43 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 sel[2]
port 44 nsew signal input
rlabel metal4 s 18194 2128 18514 22896 6 VPWR
port 45 nsew power bidirectional
rlabel metal4 s 11294 2128 11614 22896 6 VPWR
port 46 nsew power bidirectional
rlabel metal4 s 4394 2128 4714 22896 6 VPWR
port 47 nsew power bidirectional
rlabel metal5 s 1104 19195 21804 19515 6 VPWR
port 48 nsew power bidirectional
rlabel metal5 s 1104 12304 21804 12624 6 VPWR
port 49 nsew power bidirectional
rlabel metal5 s 1104 5413 21804 5733 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 14744 2128 15064 22896 6 VGND
port 51 nsew ground bidirectional
rlabel metal4 s 7844 2128 8164 22896 6 VGND
port 52 nsew ground bidirectional
rlabel metal5 s 1104 15749 21804 16069 6 VGND
port 53 nsew ground bidirectional
rlabel metal5 s 1104 8859 21804 9179 6 VGND
port 54 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 22979 25123
<< end >>
