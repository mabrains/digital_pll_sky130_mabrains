magic
tech sky130A
magscale 1 2
timestamp 1619673532
<< locali >>
rect 19165 18411 19199 19261
rect 6929 9503 6963 9605
rect 19165 1411 19199 2465
<< viali >>
rect 1501 20009 1535 20043
rect 18613 19941 18647 19975
rect 1593 19873 1627 19907
rect 1777 19873 1811 19907
rect 2329 19873 2363 19907
rect 3893 19873 3927 19907
rect 5549 19873 5583 19907
rect 6929 19873 6963 19907
rect 8309 19873 8343 19907
rect 9873 19873 9907 19907
rect 11713 19873 11747 19907
rect 13093 19873 13127 19907
rect 14749 19873 14783 19907
rect 15853 19873 15887 19907
rect 17693 19873 17727 19907
rect 18337 19873 18371 19907
rect 7113 19737 7147 19771
rect 18153 19737 18187 19771
rect 18429 19737 18463 19771
rect 1961 19669 1995 19703
rect 2513 19669 2547 19703
rect 4077 19669 4111 19703
rect 5733 19669 5767 19703
rect 8493 19669 8527 19703
rect 9689 19669 9723 19703
rect 11529 19669 11563 19703
rect 12909 19669 12943 19703
rect 14565 19669 14599 19703
rect 15669 19669 15703 19703
rect 17509 19669 17543 19703
rect 1685 19465 1719 19499
rect 2697 19329 2731 19363
rect 4813 19329 4847 19363
rect 9229 19329 9263 19363
rect 9965 19329 9999 19363
rect 17417 19329 17451 19363
rect 1869 19261 1903 19295
rect 2421 19261 2455 19295
rect 4537 19261 4571 19295
rect 6929 19261 6963 19295
rect 9505 19261 9539 19295
rect 9689 19261 9723 19295
rect 12817 19261 12851 19295
rect 15301 19261 15335 19295
rect 16589 19261 16623 19295
rect 17785 19261 17819 19295
rect 17969 19261 18003 19295
rect 18429 19261 18463 19295
rect 18521 19261 18555 19295
rect 19165 19261 19199 19295
rect 7113 19193 7147 19227
rect 7297 19193 7331 19227
rect 13093 19193 13127 19227
rect 4169 19125 4203 19159
rect 6285 19125 6319 19159
rect 7757 19125 7791 19159
rect 11437 19125 11471 19159
rect 14565 19125 14599 19159
rect 15485 19125 15519 19159
rect 16773 19125 16807 19159
rect 3433 18921 3467 18955
rect 3893 18921 3927 18955
rect 5733 18921 5767 18955
rect 9137 18921 9171 18955
rect 10609 18921 10643 18955
rect 11253 18921 11287 18955
rect 13829 18921 13863 18955
rect 16221 18921 16255 18955
rect 4629 18853 4663 18887
rect 8033 18853 8067 18887
rect 8585 18853 8619 18887
rect 11529 18853 11563 18887
rect 14749 18853 14783 18887
rect 16589 18853 16623 18887
rect 18521 18853 18555 18887
rect 3249 18785 3283 18819
rect 4077 18785 4111 18819
rect 4169 18785 4203 18819
rect 4445 18785 4479 18819
rect 4721 18785 4755 18819
rect 5917 18785 5951 18819
rect 7849 18785 7883 18819
rect 7941 18785 7975 18819
rect 8217 18785 8251 18819
rect 8355 18785 8389 18819
rect 8493 18785 8527 18819
rect 8723 18785 8757 18819
rect 9321 18785 9355 18819
rect 10425 18785 10459 18819
rect 11437 18785 11471 18819
rect 11621 18785 11655 18819
rect 11785 18785 11819 18819
rect 12081 18785 12115 18819
rect 13645 18785 13679 18819
rect 18337 18785 18371 18819
rect 14473 18717 14507 18751
rect 16313 18717 16347 18751
rect 18705 18649 18739 18683
rect 4353 18581 4387 18615
rect 7665 18581 7699 18615
rect 8861 18581 8895 18615
rect 11989 18581 12023 18615
rect 18061 18581 18095 18615
rect 18153 18581 18187 18615
rect 8217 18377 8251 18411
rect 12817 18377 12851 18411
rect 18705 18377 18739 18411
rect 19165 18377 19199 18411
rect 6745 18241 6779 18275
rect 12633 18241 12667 18275
rect 16957 18241 16991 18275
rect 17233 18241 17267 18275
rect 4721 18173 4755 18207
rect 6469 18173 6503 18207
rect 8309 18173 8343 18207
rect 8493 18173 8527 18207
rect 8861 18173 8895 18207
rect 9045 18173 9079 18207
rect 9137 18173 9171 18207
rect 11713 18173 11747 18207
rect 11897 18173 11931 18207
rect 12081 18173 12115 18207
rect 12725 18173 12759 18207
rect 13001 18173 13035 18207
rect 13093 18173 13127 18207
rect 11989 18105 12023 18139
rect 12817 18105 12851 18139
rect 4813 18037 4847 18071
rect 12265 18037 12299 18071
rect 6653 17833 6687 17867
rect 4445 17765 4479 17799
rect 1409 17697 1443 17731
rect 4629 17697 4663 17731
rect 4721 17697 4755 17731
rect 4905 17697 4939 17731
rect 6469 17697 6503 17731
rect 11069 17697 11103 17731
rect 11253 17697 11287 17731
rect 11529 17697 11563 17731
rect 11713 17697 11747 17731
rect 11897 17697 11931 17731
rect 12081 17697 12115 17731
rect 12817 17697 12851 17731
rect 13185 17697 13219 17731
rect 13369 17697 13403 17731
rect 13461 17697 13495 17731
rect 13737 17697 13771 17731
rect 14565 17697 14599 17731
rect 11805 17629 11839 17663
rect 12173 17629 12207 17663
rect 12357 17629 12391 17663
rect 12449 17629 12483 17663
rect 13553 17629 13587 17663
rect 1593 17493 1627 17527
rect 4261 17493 4295 17527
rect 4813 17493 4847 17527
rect 11161 17493 11195 17527
rect 11345 17493 11379 17527
rect 13921 17493 13955 17527
rect 14749 17493 14783 17527
rect 4445 17289 4479 17323
rect 12081 17289 12115 17323
rect 13369 17289 13403 17323
rect 16037 17289 16071 17323
rect 3341 17221 3375 17255
rect 10333 17221 10367 17255
rect 15301 17221 15335 17255
rect 1869 17153 1903 17187
rect 3709 17153 3743 17187
rect 4905 17153 4939 17187
rect 5181 17153 5215 17187
rect 9689 17153 9723 17187
rect 9873 17153 9907 17187
rect 9965 17153 9999 17187
rect 10149 17153 10183 17187
rect 15853 17153 15887 17187
rect 1593 17085 1627 17119
rect 3617 17085 3651 17119
rect 3893 17085 3927 17119
rect 4195 17085 4229 17119
rect 4353 17085 4387 17119
rect 4629 17085 4663 17119
rect 4721 17085 4755 17119
rect 4997 17085 5031 17119
rect 5089 17085 5123 17119
rect 7389 17085 7423 17119
rect 9597 17085 9631 17119
rect 10425 17085 10459 17119
rect 10701 17085 10735 17119
rect 13277 17085 13311 17119
rect 13461 17085 13495 17119
rect 13553 17085 13587 17119
rect 16313 17085 16347 17119
rect 16589 17085 16623 17119
rect 16957 17085 16991 17119
rect 17141 17085 17175 17119
rect 3985 17017 4019 17051
rect 4077 17017 4111 17051
rect 9413 17017 9447 17051
rect 10057 17017 10091 17051
rect 10149 17017 10183 17051
rect 11713 17017 11747 17051
rect 11897 17017 11931 17051
rect 13829 17017 13863 17051
rect 16497 17017 16531 17051
rect 17049 17017 17083 17051
rect 3433 16949 3467 16983
rect 7573 16949 7607 16983
rect 10609 16949 10643 16983
rect 16221 16949 16255 16983
rect 5825 16745 5859 16779
rect 16405 16745 16439 16779
rect 4997 16609 5031 16643
rect 5733 16609 5767 16643
rect 9965 16609 9999 16643
rect 10241 16609 10275 16643
rect 10425 16609 10459 16643
rect 10609 16609 10643 16643
rect 10793 16609 10827 16643
rect 16589 16609 16623 16643
rect 16773 16609 16807 16643
rect 16957 16609 16991 16643
rect 17141 16609 17175 16643
rect 18245 16609 18279 16643
rect 4721 16541 4755 16575
rect 4905 16541 4939 16575
rect 6561 16541 6595 16575
rect 6837 16541 6871 16575
rect 9505 16541 9539 16575
rect 16865 16541 16899 16575
rect 4813 16405 4847 16439
rect 8309 16405 8343 16439
rect 18061 16405 18095 16439
rect 6929 16201 6963 16235
rect 10517 16201 10551 16235
rect 10701 16201 10735 16235
rect 10885 16133 10919 16167
rect 7573 16065 7607 16099
rect 9229 16065 9263 16099
rect 9781 16065 9815 16099
rect 9965 16065 9999 16099
rect 16957 16065 16991 16099
rect 2789 15997 2823 16031
rect 7113 15997 7147 16031
rect 7205 15997 7239 16031
rect 9689 15997 9723 16031
rect 10057 15997 10091 16031
rect 10333 15997 10367 16031
rect 10425 15997 10459 16031
rect 10977 15997 11011 16031
rect 11897 15997 11931 16031
rect 12265 15997 12299 16031
rect 14473 15997 14507 16031
rect 14841 15997 14875 16031
rect 14933 15997 14967 16031
rect 15033 15997 15067 16031
rect 7297 15929 7331 15963
rect 7435 15929 7469 15963
rect 9413 15929 9447 15963
rect 12081 15929 12115 15963
rect 12173 15929 12207 15963
rect 14565 15929 14599 15963
rect 14657 15929 14691 15963
rect 17233 15929 17267 15963
rect 2973 15861 3007 15895
rect 12449 15861 12483 15895
rect 14289 15861 14323 15895
rect 15209 15861 15243 15895
rect 18705 15861 18739 15895
rect 7481 15657 7515 15691
rect 9597 15657 9631 15691
rect 11713 15657 11747 15691
rect 11989 15657 12023 15691
rect 17141 15657 17175 15691
rect 17233 15657 17267 15691
rect 4629 15589 4663 15623
rect 4813 15589 4847 15623
rect 13461 15589 13495 15623
rect 14657 15589 14691 15623
rect 16865 15589 16899 15623
rect 1409 15521 1443 15555
rect 1869 15521 1903 15555
rect 4077 15521 4111 15555
rect 4169 15521 4203 15555
rect 4261 15521 4295 15555
rect 4399 15521 4433 15555
rect 4537 15521 4571 15555
rect 4997 15521 5031 15555
rect 5181 15521 5215 15555
rect 5457 15521 5491 15555
rect 7481 15521 7515 15555
rect 7665 15521 7699 15555
rect 9505 15521 9539 15555
rect 11772 15521 11806 15555
rect 16589 15521 16623 15555
rect 16773 15521 16807 15555
rect 16957 15521 16991 15555
rect 17417 15521 17451 15555
rect 17601 15521 17635 15555
rect 17693 15521 17727 15555
rect 17969 15521 18003 15555
rect 18705 15521 18739 15555
rect 2145 15453 2179 15487
rect 3893 15453 3927 15487
rect 11253 15453 11287 15487
rect 13737 15453 13771 15487
rect 14381 15453 14415 15487
rect 11345 15385 11379 15419
rect 1593 15317 1627 15351
rect 3617 15317 3651 15351
rect 5273 15317 5307 15351
rect 5549 15317 5583 15351
rect 11897 15317 11931 15351
rect 16129 15317 16163 15351
rect 17877 15317 17911 15351
rect 18521 15317 18555 15351
rect 4721 15113 4755 15147
rect 5365 15113 5399 15147
rect 7849 15113 7883 15147
rect 9689 15113 9723 15147
rect 10425 15113 10459 15147
rect 7941 15045 7975 15079
rect 14473 15045 14507 15079
rect 5181 14977 5215 15011
rect 9873 14977 9907 15011
rect 10333 14977 10367 15011
rect 12357 14977 12391 15011
rect 4905 14909 4939 14943
rect 4997 14909 5031 14943
rect 5273 14909 5307 14943
rect 5549 14909 5583 14943
rect 5733 14909 5767 14943
rect 7297 14909 7331 14943
rect 7665 14909 7699 14943
rect 8309 14909 8343 14943
rect 9965 14909 9999 14943
rect 10793 14909 10827 14943
rect 11897 14909 11931 14943
rect 12173 14909 12207 14943
rect 12265 14909 12299 14943
rect 12461 14909 12495 14943
rect 14749 14909 14783 14943
rect 15025 14909 15059 14943
rect 17049 14909 17083 14943
rect 17233 14909 17267 14943
rect 7481 14841 7515 14875
rect 7573 14841 7607 14875
rect 8125 14841 8159 14875
rect 10609 14841 10643 14875
rect 12081 14841 12115 14875
rect 17325 14841 17359 14875
rect 11713 14773 11747 14807
rect 14657 14773 14691 14807
rect 14841 14773 14875 14807
rect 5825 14569 5859 14603
rect 10977 14569 11011 14603
rect 11161 14569 11195 14603
rect 17049 14569 17083 14603
rect 7297 14501 7331 14535
rect 1501 14433 1535 14467
rect 2053 14433 2087 14467
rect 5089 14433 5123 14467
rect 5181 14433 5215 14467
rect 5457 14433 5491 14467
rect 5641 14433 5675 14467
rect 7021 14433 7055 14467
rect 7389 14433 7423 14467
rect 7665 14433 7699 14467
rect 8125 14433 8159 14467
rect 11158 14433 11192 14467
rect 16773 14433 16807 14467
rect 16957 14433 16991 14467
rect 17233 14433 17267 14467
rect 17325 14433 17359 14467
rect 4813 14365 4847 14399
rect 5365 14365 5399 14399
rect 7297 14365 7331 14399
rect 7849 14365 7883 14399
rect 7941 14365 7975 14399
rect 11529 14365 11563 14399
rect 11621 14365 11655 14399
rect 4997 14297 5031 14331
rect 5549 14297 5583 14331
rect 7113 14297 7147 14331
rect 8033 14297 8067 14331
rect 2053 14229 2087 14263
rect 4905 14229 4939 14263
rect 7481 14229 7515 14263
rect 8309 14229 8343 14263
rect 12633 14025 12667 14059
rect 14933 14025 14967 14059
rect 15485 14025 15519 14059
rect 16405 14025 16439 14059
rect 18521 14025 18555 14059
rect 10057 13957 10091 13991
rect 17233 13957 17267 13991
rect 12817 13889 12851 13923
rect 13185 13889 13219 13923
rect 1409 13821 1443 13855
rect 2053 13821 2087 13855
rect 2513 13821 2547 13855
rect 2605 13821 2639 13855
rect 2881 13821 2915 13855
rect 4900 13821 4934 13855
rect 5272 13821 5306 13855
rect 5358 13821 5392 13855
rect 5449 13821 5483 13855
rect 5733 13821 5767 13855
rect 7200 13821 7234 13855
rect 7517 13821 7551 13855
rect 7665 13821 7699 13855
rect 7941 13821 7975 13855
rect 8953 13821 8987 13855
rect 9046 13821 9080 13855
rect 9229 13821 9263 13855
rect 9459 13821 9493 13855
rect 9681 13821 9715 13855
rect 9965 13821 9999 13855
rect 12909 13821 12943 13855
rect 13553 13821 13587 13855
rect 15025 13821 15059 13855
rect 15301 13821 15335 13855
rect 15485 13821 15519 13855
rect 16129 13821 16163 13855
rect 16305 13821 16339 13855
rect 17417 13821 17451 13855
rect 17601 13821 17635 13855
rect 17785 13821 17819 13855
rect 18705 13821 18739 13855
rect 4997 13753 5031 13787
rect 5089 13753 5123 13787
rect 5825 13753 5859 13787
rect 7297 13753 7331 13787
rect 7389 13753 7423 13787
rect 9321 13753 9355 13787
rect 9781 13753 9815 13787
rect 13277 13753 13311 13787
rect 16037 13753 16071 13787
rect 17509 13753 17543 13787
rect 1593 13685 1627 13719
rect 3065 13685 3099 13719
rect 4721 13685 4755 13719
rect 5549 13685 5583 13719
rect 7021 13685 7055 13719
rect 7849 13685 7883 13719
rect 9597 13685 9631 13719
rect 13461 13685 13495 13719
rect 15117 13685 15151 13719
rect 1501 13481 1535 13515
rect 1961 13481 1995 13515
rect 3617 13481 3651 13515
rect 9689 13481 9723 13515
rect 12541 13481 12575 13515
rect 12725 13481 12759 13515
rect 13461 13481 13495 13515
rect 17693 13481 17727 13515
rect 2697 13413 2731 13447
rect 9781 13413 9815 13447
rect 10425 13413 10459 13447
rect 13277 13413 13311 13447
rect 13737 13413 13771 13447
rect 14657 13413 14691 13447
rect 16589 13413 16623 13447
rect 1869 13345 1903 13379
rect 2605 13345 2639 13379
rect 3157 13345 3191 13379
rect 4077 13345 4111 13379
rect 9137 13345 9171 13379
rect 9413 13345 9447 13379
rect 9505 13345 9539 13379
rect 10057 13345 10091 13379
rect 12722 13345 12756 13379
rect 13185 13345 13219 13379
rect 13553 13345 13587 13379
rect 13645 13345 13679 13379
rect 13829 13345 13863 13379
rect 14381 13345 14415 13379
rect 14841 13345 14875 13379
rect 15025 13345 15059 13379
rect 15129 13345 15163 13379
rect 15577 13345 15611 13379
rect 15761 13345 15795 13379
rect 15853 13345 15887 13379
rect 16129 13345 16163 13379
rect 16313 13345 16347 13379
rect 16405 13345 16439 13379
rect 17634 13345 17668 13379
rect 18153 13345 18187 13379
rect 2053 13277 2087 13311
rect 3249 13277 3283 13311
rect 9229 13277 9263 13311
rect 9781 13277 9815 13311
rect 10149 13277 10183 13311
rect 14657 13277 14691 13311
rect 14933 13277 14967 13311
rect 15301 13277 15335 13311
rect 15945 13277 15979 13311
rect 3617 13209 3651 13243
rect 3893 13209 3927 13243
rect 9965 13209 9999 13243
rect 13093 13209 13127 13243
rect 17509 13209 17543 13243
rect 11897 13141 11931 13175
rect 13277 13141 13311 13175
rect 14473 13141 14507 13175
rect 16773 13141 16807 13175
rect 18061 13141 18095 13175
rect 8953 12937 8987 12971
rect 11345 12937 11379 12971
rect 15209 12937 15243 12971
rect 4997 12869 5031 12903
rect 5181 12869 5215 12903
rect 5641 12869 5675 12903
rect 7205 12869 7239 12903
rect 7481 12869 7515 12903
rect 7941 12869 7975 12903
rect 4813 12801 4847 12835
rect 7021 12801 7055 12835
rect 9413 12801 9447 12835
rect 5089 12733 5123 12767
rect 5365 12733 5399 12767
rect 5457 12733 5491 12767
rect 5733 12733 5767 12767
rect 7297 12733 7331 12767
rect 7665 12733 7699 12767
rect 7757 12733 7791 12767
rect 8033 12733 8067 12767
rect 11161 12733 11195 12767
rect 12173 12733 12207 12767
rect 15117 12733 15151 12767
rect 16957 12733 16991 12767
rect 17141 12733 17175 12767
rect 17325 12733 17359 12767
rect 9505 12665 9539 12699
rect 12265 12665 12299 12699
rect 17233 12665 17267 12699
rect 4813 12597 4847 12631
rect 7021 12597 7055 12631
rect 9413 12597 9447 12631
rect 17509 12597 17543 12631
rect 5825 12393 5859 12427
rect 6285 12393 6319 12427
rect 18705 12393 18739 12427
rect 1593 12325 1627 12359
rect 2881 12325 2915 12359
rect 4353 12325 4387 12359
rect 12909 12325 12943 12359
rect 17233 12325 17267 12359
rect 3065 12257 3099 12291
rect 6193 12257 6227 12291
rect 7481 12257 7515 12291
rect 10517 12257 10551 12291
rect 12679 12257 12713 12291
rect 12817 12257 12851 12291
rect 13093 12257 13127 12291
rect 13369 12257 13403 12291
rect 15301 12257 15335 12291
rect 16957 12257 16991 12291
rect 4077 12189 4111 12223
rect 1501 12053 1535 12087
rect 7665 12053 7699 12087
rect 10609 12053 10643 12087
rect 12541 12053 12575 12087
rect 13553 12053 13587 12087
rect 15117 12053 15151 12087
rect 2881 11849 2915 11883
rect 2973 11849 3007 11883
rect 4537 11849 4571 11883
rect 5181 11849 5215 11883
rect 9873 11849 9907 11883
rect 14105 11849 14139 11883
rect 18153 11849 18187 11883
rect 2237 11781 2271 11815
rect 9413 11781 9447 11815
rect 1593 11713 1627 11747
rect 1777 11713 1811 11747
rect 3341 11713 3375 11747
rect 4813 11713 4847 11747
rect 6653 11713 6687 11747
rect 6929 11713 6963 11747
rect 9321 11713 9355 11747
rect 12633 11713 12667 11747
rect 14197 11713 14231 11747
rect 15945 11713 15979 11747
rect 2329 11645 2363 11679
rect 2881 11645 2915 11679
rect 2973 11645 3007 11679
rect 4721 11645 4755 11679
rect 4905 11645 4939 11679
rect 4997 11645 5031 11679
rect 5365 11645 5399 11679
rect 9137 11645 9171 11679
rect 9505 11645 9539 11679
rect 9597 11645 9631 11679
rect 12357 11645 12391 11679
rect 16221 11645 16255 11679
rect 17049 11645 17083 11679
rect 17969 11645 18003 11679
rect 18705 11645 18739 11679
rect 1869 11577 1903 11611
rect 8401 11509 8435 11543
rect 17233 11509 17267 11543
rect 18521 11509 18555 11543
rect 2881 11305 2915 11339
rect 4169 11305 4203 11339
rect 5181 11305 5215 11339
rect 8217 11305 8251 11339
rect 17877 11305 17911 11339
rect 6101 11237 6135 11271
rect 6285 11237 6319 11271
rect 11345 11237 11379 11271
rect 16405 11237 16439 11271
rect 2789 11169 2823 11203
rect 4537 11169 4571 11203
rect 5089 11169 5123 11203
rect 8125 11169 8159 11203
rect 10425 11169 10459 11203
rect 10609 11169 10643 11203
rect 11437 11169 11471 11203
rect 16129 11169 16163 11203
rect 4445 11101 4479 11135
rect 11253 11101 11287 11135
rect 6469 11033 6503 11067
rect 10793 11033 10827 11067
rect 11805 11033 11839 11067
rect 4537 10965 4571 10999
rect 4905 10761 4939 10795
rect 6193 10761 6227 10795
rect 6745 10761 6779 10795
rect 7297 10761 7331 10795
rect 8493 10761 8527 10795
rect 9597 10761 9631 10795
rect 9965 10761 9999 10795
rect 11713 10761 11747 10795
rect 8861 10693 8895 10727
rect 11529 10693 11563 10727
rect 9413 10625 9447 10659
rect 10885 10625 10919 10659
rect 11069 10625 11103 10659
rect 12081 10625 12115 10659
rect 13461 10625 13495 10659
rect 13645 10625 13679 10659
rect 4629 10557 4663 10591
rect 6101 10557 6135 10591
rect 6653 10557 6687 10591
rect 7205 10557 7239 10591
rect 8125 10557 8159 10591
rect 8309 10557 8343 10591
rect 8493 10557 8527 10591
rect 8677 10557 8711 10591
rect 9137 10557 9171 10591
rect 9229 10557 9263 10591
rect 9505 10557 9539 10591
rect 9689 10557 9723 10591
rect 10517 10557 10551 10591
rect 10701 10557 10735 10591
rect 11161 10557 11195 10591
rect 11897 10557 11931 10591
rect 12449 10557 12483 10591
rect 15025 10557 15059 10591
rect 15393 10557 15427 10591
rect 4813 10489 4847 10523
rect 6469 10489 6503 10523
rect 9045 10489 9079 10523
rect 12633 10489 12667 10523
rect 12817 10489 12851 10523
rect 13369 10489 13403 10523
rect 8125 10421 8159 10455
rect 10609 10421 10643 10455
rect 13001 10421 13035 10455
rect 15393 10421 15427 10455
rect 3249 10217 3283 10251
rect 4721 10217 4755 10251
rect 6837 10217 6871 10251
rect 10867 10217 10901 10251
rect 11345 10217 11379 10251
rect 12817 10217 12851 10251
rect 13461 10217 13495 10251
rect 15117 10217 15151 10251
rect 15485 10217 15519 10251
rect 15577 10217 15611 10251
rect 17049 10217 17083 10251
rect 11161 10149 11195 10183
rect 13277 10149 13311 10183
rect 2237 10081 2271 10115
rect 2789 10081 2823 10115
rect 3525 10081 3559 10115
rect 4813 10081 4847 10115
rect 5457 10081 5491 10115
rect 6561 10081 6595 10115
rect 9137 10081 9171 10115
rect 9229 10081 9263 10115
rect 9413 10081 9447 10115
rect 9873 10081 9907 10115
rect 10057 10081 10091 10115
rect 10241 10081 10275 10115
rect 12633 10081 12667 10115
rect 13553 10081 13587 10115
rect 14473 10081 14507 10115
rect 15025 10081 15059 10115
rect 17141 10081 17175 10115
rect 2881 10013 2915 10047
rect 4721 10013 4755 10047
rect 5181 10013 5215 10047
rect 5273 10013 5307 10047
rect 5365 10013 5399 10047
rect 6837 10013 6871 10047
rect 9965 10013 9999 10047
rect 11437 10013 11471 10047
rect 15669 10013 15703 10047
rect 16865 10013 16899 10047
rect 2789 9945 2823 9979
rect 3249 9945 3283 9979
rect 3341 9945 3375 9979
rect 4997 9945 5031 9979
rect 10425 9945 10459 9979
rect 4261 9877 4295 9911
rect 6653 9877 6687 9911
rect 13001 9877 13035 9911
rect 14473 9877 14507 9911
rect 17509 9877 17543 9911
rect 15485 9673 15519 9707
rect 6745 9605 6779 9639
rect 6929 9605 6963 9639
rect 7665 9605 7699 9639
rect 18521 9605 18555 9639
rect 1685 9537 1719 9571
rect 4721 9537 4755 9571
rect 4813 9537 4847 9571
rect 6193 9537 6227 9571
rect 6561 9537 6595 9571
rect 7205 9537 7239 9571
rect 7389 9537 7423 9571
rect 7481 9537 7515 9571
rect 4629 9469 4663 9503
rect 4905 9469 4939 9503
rect 6101 9469 6135 9503
rect 6837 9469 6871 9503
rect 6929 9469 6963 9503
rect 7297 9469 7331 9503
rect 15669 9469 15703 9503
rect 15761 9469 15795 9503
rect 18705 9469 18739 9503
rect 1777 9401 1811 9435
rect 5089 9401 5123 9435
rect 5273 9401 5307 9435
rect 5457 9401 5491 9435
rect 15853 9401 15887 9435
rect 1869 9333 1903 9367
rect 2237 9333 2271 9367
rect 4445 9333 4479 9367
rect 6561 9333 6595 9367
rect 3893 9129 3927 9163
rect 11253 9129 11287 9163
rect 13185 9129 13219 9163
rect 14565 9129 14599 9163
rect 2605 9061 2639 9095
rect 7205 9061 7239 9095
rect 9413 9061 9447 9095
rect 9629 9061 9663 9095
rect 12633 9061 12667 9095
rect 14473 9061 14507 9095
rect 1593 8993 1627 9027
rect 4077 8993 4111 9027
rect 4353 8993 4387 9027
rect 5273 8993 5307 9027
rect 5365 8993 5399 9027
rect 6653 8993 6687 9027
rect 7297 8993 7331 9027
rect 8493 8993 8527 9027
rect 9137 8993 9171 9027
rect 11345 8993 11379 9027
rect 12541 8993 12575 9027
rect 13093 8993 13127 9027
rect 13553 8993 13587 9027
rect 5089 8925 5123 8959
rect 5181 8925 5215 8959
rect 6929 8925 6963 8959
rect 8769 8925 8803 8959
rect 9229 8925 9263 8959
rect 11161 8925 11195 8959
rect 13185 8925 13219 8959
rect 1409 8857 1443 8891
rect 2789 8857 2823 8891
rect 4261 8857 4295 8891
rect 6745 8857 6779 8891
rect 6837 8857 6871 8891
rect 8677 8857 8711 8891
rect 4905 8789 4939 8823
rect 8309 8789 8343 8823
rect 9597 8789 9631 8823
rect 9781 8789 9815 8823
rect 11713 8789 11747 8823
rect 8861 8585 8895 8619
rect 9321 8585 9355 8619
rect 12909 8585 12943 8619
rect 15025 8585 15059 8619
rect 15485 8585 15519 8619
rect 2697 8517 2731 8551
rect 2789 8517 2823 8551
rect 4445 8517 4479 8551
rect 12081 8517 12115 8551
rect 12173 8517 12207 8551
rect 18061 8517 18095 8551
rect 18153 8517 18187 8551
rect 2329 8449 2363 8483
rect 4077 8449 4111 8483
rect 5917 8449 5951 8483
rect 8217 8449 8251 8483
rect 8401 8449 8435 8483
rect 9229 8449 9263 8483
rect 11713 8449 11747 8483
rect 15117 8449 15151 8483
rect 1685 8381 1719 8415
rect 2237 8381 2271 8415
rect 2973 8381 3007 8415
rect 5825 8381 5859 8415
rect 9505 8381 9539 8415
rect 10885 8381 10919 8415
rect 11437 8381 11471 8415
rect 12357 8381 12391 8415
rect 14473 8381 14507 8415
rect 15025 8381 15059 8415
rect 15485 8381 15519 8415
rect 16497 8381 16531 8415
rect 16681 8381 16715 8415
rect 17049 8381 17083 8415
rect 17601 8381 17635 8415
rect 17693 8381 17727 8415
rect 18337 8381 18371 8415
rect 2145 8313 2179 8347
rect 3893 8313 3927 8347
rect 3985 8313 4019 8347
rect 5733 8313 5767 8347
rect 9689 8313 9723 8347
rect 11345 8313 11379 8347
rect 12817 8313 12851 8347
rect 17141 8313 17175 8347
rect 2697 8245 2731 8279
rect 5365 8245 5399 8279
rect 8493 8245 8527 8279
rect 12081 8245 12115 8279
rect 18061 8245 18095 8279
rect 2513 8041 2547 8075
rect 4353 8041 4387 8075
rect 8493 8041 8527 8075
rect 17601 8041 17635 8075
rect 4537 7973 4571 8007
rect 7481 7973 7515 8007
rect 10885 7973 10919 8007
rect 11069 7973 11103 8007
rect 7389 7905 7423 7939
rect 7573 7905 7607 7939
rect 7849 7905 7883 7939
rect 8677 7905 8711 7939
rect 8861 7905 8895 7939
rect 8953 7905 8987 7939
rect 9137 7905 9171 7939
rect 4261 7837 4295 7871
rect 9229 7837 9263 7871
rect 4813 7769 4847 7803
rect 2605 7701 2639 7735
rect 9137 7701 9171 7735
rect 9505 7701 9539 7735
rect 17509 7701 17543 7735
rect 13369 7497 13403 7531
rect 13829 7497 13863 7531
rect 2513 7429 2547 7463
rect 16773 7429 16807 7463
rect 13461 7361 13495 7395
rect 2145 7293 2179 7327
rect 3985 7293 4019 7327
rect 4261 7293 4295 7327
rect 6653 7293 6687 7327
rect 7297 7293 7331 7327
rect 10977 7293 11011 7327
rect 12817 7293 12851 7327
rect 13369 7293 13403 7327
rect 13829 7293 13863 7327
rect 15761 7293 15795 7327
rect 16307 7293 16341 7327
rect 16405 7293 16439 7327
rect 11161 7225 11195 7259
rect 16221 7225 16255 7259
rect 2513 7157 2547 7191
rect 3801 7157 3835 7191
rect 4169 7157 4203 7191
rect 7757 7157 7791 7191
rect 11345 7157 11379 7191
rect 16773 7157 16807 7191
rect 2145 6953 2179 6987
rect 8769 6953 8803 6987
rect 12081 6953 12115 6987
rect 13369 6953 13403 6987
rect 13829 6953 13863 6987
rect 4813 6885 4847 6919
rect 7297 6885 7331 6919
rect 16497 6885 16531 6919
rect 1409 6817 1443 6851
rect 2605 6817 2639 6851
rect 3157 6817 3191 6851
rect 4721 6817 4755 6851
rect 4997 6817 5031 6851
rect 5733 6817 5767 6851
rect 5917 6817 5951 6851
rect 6285 6817 6319 6851
rect 6653 6817 6687 6851
rect 7573 6817 7607 6851
rect 7665 6817 7699 6851
rect 8401 6817 8435 6851
rect 9965 6817 9999 6851
rect 10701 6817 10735 6851
rect 10885 6817 10919 6851
rect 13645 6817 13679 6851
rect 14749 6817 14783 6851
rect 16313 6817 16347 6851
rect 18705 6817 18739 6851
rect 1961 6749 1995 6783
rect 2053 6749 2087 6783
rect 11897 6749 11931 6783
rect 11989 6749 12023 6783
rect 14841 6749 14875 6783
rect 15025 6749 15059 6783
rect 1593 6681 1627 6715
rect 2513 6681 2547 6715
rect 5273 6681 5307 6715
rect 8769 6681 8803 6715
rect 18521 6681 18555 6715
rect 3157 6613 3191 6647
rect 12449 6613 12483 6647
rect 13277 6613 13311 6647
rect 14381 6613 14415 6647
rect 9781 6409 9815 6443
rect 12725 6341 12759 6375
rect 6929 6273 6963 6307
rect 14657 6273 14691 6307
rect 6561 6205 6595 6239
rect 7021 6205 7055 6239
rect 7941 6205 7975 6239
rect 8125 6205 8159 6239
rect 9137 6205 9171 6239
rect 9689 6205 9723 6239
rect 9965 6205 9999 6239
rect 10241 6205 10275 6239
rect 10977 6205 11011 6239
rect 12357 6205 12391 6239
rect 14841 6205 14875 6239
rect 15025 6205 15059 6239
rect 15301 6205 15335 6239
rect 6745 6137 6779 6171
rect 7665 6137 7699 6171
rect 8769 6137 8803 6171
rect 9045 6137 9079 6171
rect 9597 6137 9631 6171
rect 10885 6137 10919 6171
rect 12725 6069 12759 6103
rect 3157 5865 3191 5899
rect 6653 5865 6687 5899
rect 7021 5865 7055 5899
rect 8309 5865 8343 5899
rect 8401 5865 8435 5899
rect 10793 5865 10827 5899
rect 14657 5865 14691 5899
rect 15117 5865 15151 5899
rect 15301 5865 15335 5899
rect 3249 5797 3283 5831
rect 4629 5797 4663 5831
rect 5365 5797 5399 5831
rect 12541 5797 12575 5831
rect 16313 5797 16347 5831
rect 3893 5729 3927 5763
rect 4813 5729 4847 5763
rect 5457 5729 5491 5763
rect 5549 5729 5583 5763
rect 5733 5729 5767 5763
rect 10701 5729 10735 5763
rect 12081 5729 12115 5763
rect 12633 5729 12667 5763
rect 14749 5729 14783 5763
rect 15301 5729 15335 5763
rect 15485 5729 15519 5763
rect 15669 5729 15703 5763
rect 16129 5729 16163 5763
rect 16221 5729 16255 5763
rect 4905 5661 4939 5695
rect 7113 5661 7147 5695
rect 7297 5661 7331 5695
rect 14565 5661 14599 5695
rect 16037 5661 16071 5695
rect 5917 5253 5951 5287
rect 6009 5253 6043 5287
rect 16313 5185 16347 5219
rect 2938 5117 2972 5151
rect 4905 5117 4939 5151
rect 5457 5117 5491 5151
rect 5549 5117 5583 5151
rect 6193 5117 6227 5151
rect 12633 5117 12667 5151
rect 15301 5117 15335 5151
rect 15485 5117 15519 5151
rect 15669 5117 15703 5151
rect 15853 5117 15887 5151
rect 16221 5117 16255 5151
rect 4997 5049 5031 5083
rect 12449 5049 12483 5083
rect 2835 4981 2869 5015
rect 5917 4981 5951 5015
rect 15669 4981 15703 5015
rect 16405 4981 16439 5015
rect 1501 4777 1535 4811
rect 6377 4777 6411 4811
rect 7665 4777 7699 4811
rect 11069 4777 11103 4811
rect 15025 4777 15059 4811
rect 15393 4777 15427 4811
rect 16037 4777 16071 4811
rect 18521 4777 18555 4811
rect 3341 4709 3375 4743
rect 6469 4709 6503 4743
rect 1593 4641 1627 4675
rect 2421 4641 2455 4675
rect 10057 4641 10091 4675
rect 10609 4641 10643 4675
rect 10701 4641 10735 4675
rect 11345 4641 11379 4675
rect 12265 4641 12299 4675
rect 16405 4641 16439 4675
rect 18705 4641 18739 4675
rect 7297 4573 7331 4607
rect 11621 4573 11655 4607
rect 15485 4573 15519 4607
rect 15669 4573 15703 4607
rect 16497 4573 16531 4607
rect 16589 4573 16623 4607
rect 3525 4505 3559 4539
rect 7665 4505 7699 4539
rect 11069 4505 11103 4539
rect 11161 4505 11195 4539
rect 2329 4437 2363 4471
rect 10609 4437 10643 4471
rect 7665 4233 7699 4267
rect 10609 4233 10643 4267
rect 7113 4097 7147 4131
rect 8125 4097 8159 4131
rect 9965 4097 9999 4131
rect 11897 4097 11931 4131
rect 13185 4097 13219 4131
rect 7297 4029 7331 4063
rect 7757 4029 7791 4063
rect 8309 4029 8343 4063
rect 10241 4029 10275 4063
rect 12541 4029 12575 4063
rect 13093 4029 13127 4063
rect 13553 4029 13587 4063
rect 13829 4029 13863 4063
rect 10149 3961 10183 3995
rect 12081 3961 12115 3995
rect 13001 3961 13035 3995
rect 7205 3893 7239 3927
rect 11989 3893 12023 3927
rect 12449 3893 12483 3927
rect 13553 3893 13587 3927
rect 13645 3893 13679 3927
rect 11161 3689 11195 3723
rect 13921 3689 13955 3723
rect 6009 3621 6043 3655
rect 8125 3621 8159 3655
rect 8309 3553 8343 3587
rect 11069 3553 11103 3587
rect 14749 3553 14783 3587
rect 17601 3553 17635 3587
rect 6285 3485 6319 3519
rect 14841 3485 14875 3519
rect 15025 3485 15059 3519
rect 15577 3485 15611 3519
rect 15853 3485 15887 3519
rect 4277 3349 4311 3383
rect 14013 3349 14047 3383
rect 14381 3349 14415 3383
rect 5917 3145 5951 3179
rect 8401 3145 8435 3179
rect 9597 3145 9631 3179
rect 10517 3145 10551 3179
rect 10977 3145 11011 3179
rect 12081 3145 12115 3179
rect 13093 3145 13127 3179
rect 18521 3145 18555 3179
rect 5043 3077 5077 3111
rect 8861 3077 8895 3111
rect 8953 3077 8987 3111
rect 3065 3009 3099 3043
rect 3341 3009 3375 3043
rect 10609 3009 10643 3043
rect 12725 3009 12759 3043
rect 16773 3009 16807 3043
rect 1409 2941 1443 2975
rect 5825 2941 5859 2975
rect 7849 2941 7883 2975
rect 8401 2941 8435 2975
rect 8493 2941 8527 2975
rect 9137 2941 9171 2975
rect 9505 2941 9539 2975
rect 9965 2941 9999 2975
rect 10517 2941 10551 2975
rect 10977 2941 11011 2975
rect 11805 2941 11839 2975
rect 11989 2941 12023 2975
rect 12081 2941 12115 2975
rect 12633 2941 12667 2975
rect 13093 2941 13127 2975
rect 13737 2941 13771 2975
rect 14289 2941 14323 2975
rect 18705 2941 18739 2975
rect 13829 2873 13863 2907
rect 14565 2873 14599 2907
rect 16497 2873 16531 2907
rect 1593 2805 1627 2839
rect 8861 2805 8895 2839
rect 14473 2805 14507 2839
rect 14749 2805 14783 2839
rect 1593 2601 1627 2635
rect 3433 2601 3467 2635
rect 4813 2601 4847 2635
rect 6009 2601 6043 2635
rect 7941 2601 7975 2635
rect 8401 2601 8435 2635
rect 8677 2601 8711 2635
rect 9505 2601 9539 2635
rect 9597 2601 9631 2635
rect 9965 2601 9999 2635
rect 10609 2601 10643 2635
rect 12173 2601 12207 2635
rect 13001 2601 13035 2635
rect 14013 2601 14047 2635
rect 15577 2601 15611 2635
rect 16589 2601 16623 2635
rect 18521 2601 18555 2635
rect 2053 2533 2087 2567
rect 10333 2533 10367 2567
rect 15025 2533 15059 2567
rect 15485 2533 15519 2567
rect 18153 2533 18187 2567
rect 1409 2465 1443 2499
rect 3249 2465 3283 2499
rect 4629 2465 4663 2499
rect 6193 2465 6227 2499
rect 8033 2465 8067 2499
rect 8493 2465 8527 2499
rect 10149 2465 10183 2499
rect 10793 2465 10827 2499
rect 11989 2465 12023 2499
rect 12817 2465 12851 2499
rect 14013 2465 14047 2499
rect 14381 2465 14415 2499
rect 14657 2465 14691 2499
rect 16773 2465 16807 2499
rect 18705 2465 18739 2499
rect 19165 2465 19199 2499
rect 7757 2397 7791 2431
rect 9321 2397 9355 2431
rect 1869 2329 1903 2363
rect 17969 2329 18003 2363
rect 19165 1377 19199 1411
<< metal1 >>
rect 1104 20154 19044 20176
rect 1104 20102 6962 20154
rect 7014 20102 7026 20154
rect 7078 20102 7090 20154
rect 7142 20102 7154 20154
rect 7206 20102 12942 20154
rect 12994 20102 13006 20154
rect 13058 20102 13070 20154
rect 13122 20102 13134 20154
rect 13186 20102 19044 20154
rect 1104 20080 19044 20102
rect 1486 20040 1492 20052
rect 1447 20012 1492 20040
rect 1486 20000 1492 20012
rect 1544 20000 1550 20052
rect 934 19932 940 19984
rect 992 19972 998 19984
rect 18601 19975 18659 19981
rect 992 19944 1808 19972
rect 992 19932 998 19944
rect 1578 19904 1584 19916
rect 1539 19876 1584 19904
rect 1578 19864 1584 19876
rect 1636 19864 1642 19916
rect 1780 19913 1808 19944
rect 18601 19941 18613 19975
rect 18647 19972 18659 19975
rect 18874 19972 18880 19984
rect 18647 19944 18880 19972
rect 18647 19941 18659 19944
rect 18601 19935 18659 19941
rect 18874 19932 18880 19944
rect 18932 19932 18938 19984
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19873 1823 19907
rect 2314 19904 2320 19916
rect 2275 19876 2320 19904
rect 1765 19867 1823 19873
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 3694 19864 3700 19916
rect 3752 19904 3758 19916
rect 3881 19907 3939 19913
rect 3881 19904 3893 19907
rect 3752 19876 3893 19904
rect 3752 19864 3758 19876
rect 3881 19873 3893 19876
rect 3927 19873 3939 19907
rect 5534 19904 5540 19916
rect 5495 19876 5540 19904
rect 3881 19867 3939 19873
rect 5534 19864 5540 19876
rect 5592 19864 5598 19916
rect 6914 19904 6920 19916
rect 6875 19876 6920 19904
rect 6914 19864 6920 19876
rect 6972 19864 6978 19916
rect 8294 19904 8300 19916
rect 8255 19876 8300 19904
rect 8294 19864 8300 19876
rect 8352 19864 8358 19916
rect 9674 19864 9680 19916
rect 9732 19904 9738 19916
rect 9861 19907 9919 19913
rect 9861 19904 9873 19907
rect 9732 19876 9873 19904
rect 9732 19864 9738 19876
rect 9861 19873 9873 19876
rect 9907 19873 9919 19907
rect 9861 19867 9919 19873
rect 11514 19864 11520 19916
rect 11572 19904 11578 19916
rect 11701 19907 11759 19913
rect 11701 19904 11713 19907
rect 11572 19876 11713 19904
rect 11572 19864 11578 19876
rect 11701 19873 11713 19876
rect 11747 19873 11759 19907
rect 11701 19867 11759 19873
rect 12802 19864 12808 19916
rect 12860 19904 12866 19916
rect 13081 19907 13139 19913
rect 13081 19904 13093 19907
rect 12860 19876 13093 19904
rect 12860 19864 12866 19876
rect 13081 19873 13093 19876
rect 13127 19873 13139 19907
rect 13081 19867 13139 19873
rect 14274 19864 14280 19916
rect 14332 19904 14338 19916
rect 14737 19907 14795 19913
rect 14737 19904 14749 19907
rect 14332 19876 14749 19904
rect 14332 19864 14338 19876
rect 14737 19873 14749 19876
rect 14783 19873 14795 19907
rect 14737 19867 14795 19873
rect 15654 19864 15660 19916
rect 15712 19904 15718 19916
rect 15841 19907 15899 19913
rect 15841 19904 15853 19907
rect 15712 19876 15853 19904
rect 15712 19864 15718 19876
rect 15841 19873 15853 19876
rect 15887 19873 15899 19907
rect 15841 19867 15899 19873
rect 17494 19864 17500 19916
rect 17552 19904 17558 19916
rect 17681 19907 17739 19913
rect 17681 19904 17693 19907
rect 17552 19876 17693 19904
rect 17552 19864 17558 19876
rect 17681 19873 17693 19876
rect 17727 19873 17739 19907
rect 18322 19904 18328 19916
rect 18283 19876 18328 19904
rect 17681 19867 17739 19873
rect 18322 19864 18328 19876
rect 18380 19864 18386 19916
rect 7101 19771 7159 19777
rect 7101 19737 7113 19771
rect 7147 19768 7159 19771
rect 9582 19768 9588 19780
rect 7147 19740 9588 19768
rect 7147 19737 7159 19740
rect 7101 19731 7159 19737
rect 9582 19728 9588 19740
rect 9640 19728 9646 19780
rect 13630 19728 13636 19780
rect 13688 19768 13694 19780
rect 18141 19771 18199 19777
rect 18141 19768 18153 19771
rect 13688 19740 18153 19768
rect 13688 19728 13694 19740
rect 18141 19737 18153 19740
rect 18187 19737 18199 19771
rect 18414 19768 18420 19780
rect 18375 19740 18420 19768
rect 18141 19731 18199 19737
rect 18414 19728 18420 19740
rect 18472 19728 18478 19780
rect 1946 19700 1952 19712
rect 1907 19672 1952 19700
rect 1946 19660 1952 19672
rect 2004 19660 2010 19712
rect 2498 19700 2504 19712
rect 2459 19672 2504 19700
rect 2498 19660 2504 19672
rect 2556 19660 2562 19712
rect 3694 19660 3700 19712
rect 3752 19700 3758 19712
rect 4065 19703 4123 19709
rect 4065 19700 4077 19703
rect 3752 19672 4077 19700
rect 3752 19660 3758 19672
rect 4065 19669 4077 19672
rect 4111 19669 4123 19703
rect 4065 19663 4123 19669
rect 5721 19703 5779 19709
rect 5721 19669 5733 19703
rect 5767 19700 5779 19703
rect 5994 19700 6000 19712
rect 5767 19672 6000 19700
rect 5767 19669 5779 19672
rect 5721 19663 5779 19669
rect 5994 19660 6000 19672
rect 6052 19660 6058 19712
rect 8386 19660 8392 19712
rect 8444 19700 8450 19712
rect 8481 19703 8539 19709
rect 8481 19700 8493 19703
rect 8444 19672 8493 19700
rect 8444 19660 8450 19672
rect 8481 19669 8493 19672
rect 8527 19669 8539 19703
rect 8481 19663 8539 19669
rect 9677 19703 9735 19709
rect 9677 19669 9689 19703
rect 9723 19700 9735 19703
rect 10502 19700 10508 19712
rect 9723 19672 10508 19700
rect 9723 19669 9735 19672
rect 9677 19663 9735 19669
rect 10502 19660 10508 19672
rect 10560 19660 10566 19712
rect 11517 19703 11575 19709
rect 11517 19669 11529 19703
rect 11563 19700 11575 19703
rect 11606 19700 11612 19712
rect 11563 19672 11612 19700
rect 11563 19669 11575 19672
rect 11517 19663 11575 19669
rect 11606 19660 11612 19672
rect 11664 19660 11670 19712
rect 11882 19660 11888 19712
rect 11940 19700 11946 19712
rect 12897 19703 12955 19709
rect 12897 19700 12909 19703
rect 11940 19672 12909 19700
rect 11940 19660 11946 19672
rect 12897 19669 12909 19672
rect 12943 19669 12955 19703
rect 12897 19663 12955 19669
rect 14366 19660 14372 19712
rect 14424 19700 14430 19712
rect 14553 19703 14611 19709
rect 14553 19700 14565 19703
rect 14424 19672 14565 19700
rect 14424 19660 14430 19672
rect 14553 19669 14565 19672
rect 14599 19669 14611 19703
rect 15654 19700 15660 19712
rect 15615 19672 15660 19700
rect 14553 19663 14611 19669
rect 15654 19660 15660 19672
rect 15712 19660 15718 19712
rect 17494 19700 17500 19712
rect 17455 19672 17500 19700
rect 17494 19660 17500 19672
rect 17552 19660 17558 19712
rect 1104 19610 19044 19632
rect 1104 19558 3972 19610
rect 4024 19558 4036 19610
rect 4088 19558 4100 19610
rect 4152 19558 4164 19610
rect 4216 19558 9952 19610
rect 10004 19558 10016 19610
rect 10068 19558 10080 19610
rect 10132 19558 10144 19610
rect 10196 19558 15932 19610
rect 15984 19558 15996 19610
rect 16048 19558 16060 19610
rect 16112 19558 16124 19610
rect 16176 19558 19044 19610
rect 1104 19536 19044 19558
rect 1578 19456 1584 19508
rect 1636 19496 1642 19508
rect 1673 19499 1731 19505
rect 1673 19496 1685 19499
rect 1636 19468 1685 19496
rect 1636 19456 1642 19468
rect 1673 19465 1685 19468
rect 1719 19465 1731 19499
rect 1673 19459 1731 19465
rect 2685 19363 2743 19369
rect 2685 19329 2697 19363
rect 2731 19360 2743 19363
rect 3878 19360 3884 19372
rect 2731 19332 3884 19360
rect 2731 19329 2743 19332
rect 2685 19323 2743 19329
rect 3878 19320 3884 19332
rect 3936 19320 3942 19372
rect 4801 19363 4859 19369
rect 4801 19329 4813 19363
rect 4847 19360 4859 19363
rect 4847 19332 6040 19360
rect 4847 19329 4859 19332
rect 4801 19323 4859 19329
rect 1854 19292 1860 19304
rect 1767 19264 1860 19292
rect 1854 19252 1860 19264
rect 1912 19292 1918 19304
rect 2409 19295 2467 19301
rect 2409 19292 2421 19295
rect 1912 19264 2421 19292
rect 1912 19252 1918 19264
rect 2409 19261 2421 19264
rect 2455 19261 2467 19295
rect 2409 19255 2467 19261
rect 4525 19295 4583 19301
rect 4525 19261 4537 19295
rect 4571 19261 4583 19295
rect 6012 19292 6040 19332
rect 8036 19332 8248 19360
rect 6917 19295 6975 19301
rect 6917 19292 6929 19295
rect 6012 19264 6929 19292
rect 4525 19255 4583 19261
rect 6917 19261 6929 19264
rect 6963 19261 6975 19295
rect 8036 19292 8064 19332
rect 8220 19304 8248 19332
rect 8846 19320 8852 19372
rect 8904 19360 8910 19372
rect 9217 19363 9275 19369
rect 9217 19360 9229 19363
rect 8904 19332 9229 19360
rect 8904 19320 8910 19332
rect 9217 19329 9229 19332
rect 9263 19329 9275 19363
rect 9217 19323 9275 19329
rect 9953 19363 10011 19369
rect 9953 19329 9965 19363
rect 9999 19360 10011 19363
rect 11238 19360 11244 19372
rect 9999 19332 11244 19360
rect 9999 19329 10011 19332
rect 9953 19323 10011 19329
rect 11238 19320 11244 19332
rect 11296 19320 11302 19372
rect 17310 19320 17316 19372
rect 17368 19360 17374 19372
rect 17405 19363 17463 19369
rect 17405 19360 17417 19363
rect 17368 19332 17417 19360
rect 17368 19320 17374 19332
rect 17405 19329 17417 19332
rect 17451 19329 17463 19363
rect 17405 19323 17463 19329
rect 18340 19332 18552 19360
rect 6917 19255 6975 19261
rect 7024 19264 8064 19292
rect 2424 19156 2452 19255
rect 3418 19184 3424 19236
rect 3476 19184 3482 19236
rect 4540 19224 4568 19255
rect 4798 19224 4804 19236
rect 3988 19196 4804 19224
rect 3988 19156 4016 19196
rect 4798 19184 4804 19196
rect 4856 19184 4862 19236
rect 5810 19184 5816 19236
rect 5868 19184 5874 19236
rect 6454 19184 6460 19236
rect 6512 19224 6518 19236
rect 7024 19224 7052 19264
rect 8202 19252 8208 19304
rect 8260 19252 8266 19304
rect 9493 19295 9551 19301
rect 9493 19261 9505 19295
rect 9539 19292 9551 19295
rect 9677 19295 9735 19301
rect 9677 19292 9689 19295
rect 9539 19264 9689 19292
rect 9539 19261 9551 19264
rect 9493 19255 9551 19261
rect 6512 19196 7052 19224
rect 7101 19227 7159 19233
rect 6512 19184 6518 19196
rect 7101 19193 7113 19227
rect 7147 19193 7159 19227
rect 7282 19224 7288 19236
rect 7243 19196 7288 19224
rect 7101 19187 7159 19193
rect 2424 19128 4016 19156
rect 4157 19159 4215 19165
rect 4157 19125 4169 19159
rect 4203 19156 4215 19159
rect 4430 19156 4436 19168
rect 4203 19128 4436 19156
rect 4203 19125 4215 19128
rect 4157 19119 4215 19125
rect 4430 19116 4436 19128
rect 4488 19116 4494 19168
rect 6273 19159 6331 19165
rect 6273 19125 6285 19159
rect 6319 19156 6331 19159
rect 7116 19156 7144 19187
rect 7282 19184 7288 19196
rect 7340 19184 7346 19236
rect 9122 19224 9128 19236
rect 8786 19196 9128 19224
rect 9122 19184 9128 19196
rect 9180 19184 9186 19236
rect 7558 19156 7564 19168
rect 6319 19128 7564 19156
rect 6319 19125 6331 19128
rect 6273 19119 6331 19125
rect 7558 19116 7564 19128
rect 7616 19116 7622 19168
rect 7745 19159 7803 19165
rect 7745 19125 7757 19159
rect 7791 19156 7803 19159
rect 7926 19156 7932 19168
rect 7791 19128 7932 19156
rect 7791 19125 7803 19128
rect 7745 19119 7803 19125
rect 7926 19116 7932 19128
rect 7984 19116 7990 19168
rect 8202 19116 8208 19168
rect 8260 19156 8266 19168
rect 9600 19156 9628 19264
rect 9677 19261 9689 19264
rect 9723 19261 9735 19295
rect 12618 19292 12624 19304
rect 9677 19255 9735 19261
rect 11256 19264 12624 19292
rect 10594 19184 10600 19236
rect 10652 19184 10658 19236
rect 11256 19156 11284 19264
rect 12618 19252 12624 19264
rect 12676 19292 12682 19304
rect 12805 19295 12863 19301
rect 12805 19292 12817 19295
rect 12676 19264 12817 19292
rect 12676 19252 12682 19264
rect 12805 19261 12817 19264
rect 12851 19261 12863 19295
rect 12805 19255 12863 19261
rect 15010 19252 15016 19304
rect 15068 19292 15074 19304
rect 15289 19295 15347 19301
rect 15289 19292 15301 19295
rect 15068 19264 15301 19292
rect 15068 19252 15074 19264
rect 15289 19261 15301 19264
rect 15335 19292 15347 19295
rect 16577 19295 16635 19301
rect 16577 19292 16589 19295
rect 15335 19264 16589 19292
rect 15335 19261 15347 19264
rect 15289 19255 15347 19261
rect 16577 19261 16589 19264
rect 16623 19261 16635 19295
rect 16577 19255 16635 19261
rect 13081 19227 13139 19233
rect 13081 19193 13093 19227
rect 13127 19193 13139 19227
rect 13081 19187 13139 19193
rect 8260 19128 11284 19156
rect 11425 19159 11483 19165
rect 8260 19116 8266 19128
rect 11425 19125 11437 19159
rect 11471 19156 11483 19159
rect 11514 19156 11520 19168
rect 11471 19128 11520 19156
rect 11471 19125 11483 19128
rect 11425 19119 11483 19125
rect 11514 19116 11520 19128
rect 11572 19116 11578 19168
rect 12802 19116 12808 19168
rect 12860 19156 12866 19168
rect 13096 19156 13124 19187
rect 13814 19184 13820 19236
rect 13872 19184 13878 19236
rect 16592 19224 16620 19255
rect 17218 19252 17224 19304
rect 17276 19292 17282 19304
rect 17773 19295 17831 19301
rect 17773 19292 17785 19295
rect 17276 19264 17785 19292
rect 17276 19252 17282 19264
rect 17773 19261 17785 19264
rect 17819 19261 17831 19295
rect 17773 19255 17831 19261
rect 17957 19295 18015 19301
rect 17957 19261 17969 19295
rect 18003 19292 18015 19295
rect 18340 19292 18368 19332
rect 18524 19301 18552 19332
rect 18003 19264 18368 19292
rect 18417 19295 18475 19301
rect 18003 19261 18015 19264
rect 17957 19255 18015 19261
rect 18417 19261 18429 19295
rect 18463 19261 18475 19295
rect 18417 19255 18475 19261
rect 18509 19295 18567 19301
rect 18509 19261 18521 19295
rect 18555 19292 18567 19295
rect 19153 19295 19211 19301
rect 19153 19292 19165 19295
rect 18555 19264 19165 19292
rect 18555 19261 18567 19264
rect 18509 19255 18567 19261
rect 19153 19261 19165 19264
rect 19199 19261 19211 19295
rect 19153 19255 19211 19261
rect 17788 19224 17816 19255
rect 18432 19224 18460 19255
rect 16592 19196 17724 19224
rect 17788 19196 18460 19224
rect 12860 19128 13124 19156
rect 12860 19116 12866 19128
rect 13722 19116 13728 19168
rect 13780 19156 13786 19168
rect 14553 19159 14611 19165
rect 14553 19156 14565 19159
rect 13780 19128 14565 19156
rect 13780 19116 13786 19128
rect 14553 19125 14565 19128
rect 14599 19125 14611 19159
rect 15470 19156 15476 19168
rect 15431 19128 15476 19156
rect 14553 19119 14611 19125
rect 15470 19116 15476 19128
rect 15528 19116 15534 19168
rect 16761 19159 16819 19165
rect 16761 19125 16773 19159
rect 16807 19156 16819 19159
rect 17034 19156 17040 19168
rect 16807 19128 17040 19156
rect 16807 19125 16819 19128
rect 16761 19119 16819 19125
rect 17034 19116 17040 19128
rect 17092 19116 17098 19168
rect 17696 19156 17724 19196
rect 18046 19156 18052 19168
rect 17696 19128 18052 19156
rect 18046 19116 18052 19128
rect 18104 19116 18110 19168
rect 1104 19066 19044 19088
rect 1104 19014 6962 19066
rect 7014 19014 7026 19066
rect 7078 19014 7090 19066
rect 7142 19014 7154 19066
rect 7206 19014 12942 19066
rect 12994 19014 13006 19066
rect 13058 19014 13070 19066
rect 13122 19014 13134 19066
rect 13186 19014 19044 19066
rect 1104 18992 19044 19014
rect 3418 18952 3424 18964
rect 3379 18924 3424 18952
rect 3418 18912 3424 18924
rect 3476 18912 3482 18964
rect 3878 18952 3884 18964
rect 3839 18924 3884 18952
rect 3878 18912 3884 18924
rect 3936 18912 3942 18964
rect 5721 18955 5779 18961
rect 5721 18921 5733 18955
rect 5767 18952 5779 18955
rect 5810 18952 5816 18964
rect 5767 18924 5816 18952
rect 5767 18921 5779 18924
rect 5721 18915 5779 18921
rect 5810 18912 5816 18924
rect 5868 18912 5874 18964
rect 9122 18952 9128 18964
rect 8312 18924 8800 18952
rect 9083 18924 9128 18952
rect 4617 18887 4675 18893
rect 4617 18884 4629 18887
rect 4080 18856 4629 18884
rect 3237 18819 3295 18825
rect 3237 18785 3249 18819
rect 3283 18816 3295 18819
rect 3602 18816 3608 18828
rect 3283 18788 3608 18816
rect 3283 18785 3295 18788
rect 3237 18779 3295 18785
rect 3602 18776 3608 18788
rect 3660 18776 3666 18828
rect 4080 18825 4108 18856
rect 4617 18853 4629 18856
rect 4663 18853 4675 18887
rect 4617 18847 4675 18853
rect 7742 18844 7748 18896
rect 7800 18884 7806 18896
rect 8021 18887 8079 18893
rect 8021 18884 8033 18887
rect 7800 18856 8033 18884
rect 7800 18844 7806 18856
rect 8021 18853 8033 18856
rect 8067 18853 8079 18887
rect 8312 18884 8340 18924
rect 8021 18847 8079 18853
rect 8220 18856 8340 18884
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18785 4123 18819
rect 4065 18779 4123 18785
rect 4157 18819 4215 18825
rect 4157 18785 4169 18819
rect 4203 18785 4215 18819
rect 4430 18816 4436 18828
rect 4391 18788 4436 18816
rect 4157 18779 4215 18785
rect 4172 18748 4200 18779
rect 4430 18776 4436 18788
rect 4488 18816 4494 18828
rect 4709 18819 4767 18825
rect 4709 18816 4721 18819
rect 4488 18788 4721 18816
rect 4488 18776 4494 18788
rect 4709 18785 4721 18788
rect 4755 18785 4767 18819
rect 4709 18779 4767 18785
rect 5905 18819 5963 18825
rect 5905 18785 5917 18819
rect 5951 18785 5963 18819
rect 5905 18779 5963 18785
rect 4614 18748 4620 18760
rect 4172 18720 4620 18748
rect 4614 18708 4620 18720
rect 4672 18708 4678 18760
rect 5920 18748 5948 18779
rect 7282 18776 7288 18828
rect 7340 18816 7346 18828
rect 7837 18819 7895 18825
rect 7837 18816 7849 18819
rect 7340 18788 7849 18816
rect 7340 18776 7346 18788
rect 7837 18785 7849 18788
rect 7883 18785 7895 18819
rect 7837 18779 7895 18785
rect 7374 18748 7380 18760
rect 5920 18720 7380 18748
rect 7374 18708 7380 18720
rect 7432 18708 7438 18760
rect 7852 18748 7880 18779
rect 7926 18776 7932 18828
rect 7984 18816 7990 18828
rect 8220 18825 8248 18856
rect 8570 18844 8576 18896
rect 8628 18884 8634 18896
rect 8772 18884 8800 18924
rect 9122 18912 9128 18924
rect 9180 18912 9186 18964
rect 10594 18952 10600 18964
rect 10555 18924 10600 18952
rect 10594 18912 10600 18924
rect 10652 18912 10658 18964
rect 11238 18952 11244 18964
rect 11199 18924 11244 18952
rect 11238 18912 11244 18924
rect 11296 18912 11302 18964
rect 12342 18952 12348 18964
rect 11348 18924 12348 18952
rect 11348 18884 11376 18924
rect 12342 18912 12348 18924
rect 12400 18912 12406 18964
rect 13814 18952 13820 18964
rect 13775 18924 13820 18952
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 15654 18952 15660 18964
rect 14752 18924 15660 18952
rect 11514 18884 11520 18896
rect 8628 18856 8673 18884
rect 8772 18856 11376 18884
rect 11475 18856 11520 18884
rect 8628 18844 8634 18856
rect 8205 18819 8263 18825
rect 7984 18788 8029 18816
rect 7984 18776 7990 18788
rect 8205 18785 8217 18819
rect 8251 18785 8263 18819
rect 8205 18779 8263 18785
rect 8343 18819 8401 18825
rect 8343 18785 8355 18819
rect 8389 18785 8401 18819
rect 8343 18779 8401 18785
rect 8481 18819 8539 18825
rect 8481 18785 8493 18819
rect 8527 18785 8539 18819
rect 8481 18779 8539 18785
rect 8711 18819 8769 18825
rect 8711 18785 8723 18819
rect 8757 18816 8769 18819
rect 8864 18816 8892 18856
rect 9306 18816 9312 18828
rect 8757 18788 8892 18816
rect 9267 18788 9312 18816
rect 8757 18785 8769 18788
rect 8711 18779 8769 18785
rect 8358 18748 8386 18779
rect 7852 18720 8386 18748
rect 8220 18692 8248 18720
rect 7558 18640 7564 18692
rect 7616 18680 7622 18692
rect 7616 18652 7880 18680
rect 7616 18640 7622 18652
rect 4338 18612 4344 18624
rect 4299 18584 4344 18612
rect 4338 18572 4344 18584
rect 4396 18572 4402 18624
rect 6730 18572 6736 18624
rect 6788 18612 6794 18624
rect 7653 18615 7711 18621
rect 7653 18612 7665 18615
rect 6788 18584 7665 18612
rect 6788 18572 6794 18584
rect 7653 18581 7665 18584
rect 7699 18581 7711 18615
rect 7852 18612 7880 18652
rect 8202 18640 8208 18692
rect 8260 18640 8266 18692
rect 8294 18612 8300 18624
rect 7852 18584 8300 18612
rect 7653 18575 7711 18581
rect 8294 18572 8300 18584
rect 8352 18612 8358 18624
rect 8496 18612 8524 18779
rect 9306 18776 9312 18788
rect 9364 18816 9370 18828
rect 10413 18819 10471 18825
rect 10413 18816 10425 18819
rect 9364 18788 10425 18816
rect 9364 18776 9370 18788
rect 10413 18785 10425 18788
rect 10459 18785 10471 18819
rect 11348 18816 11376 18856
rect 11514 18844 11520 18856
rect 11572 18884 11578 18896
rect 14752 18893 14780 18924
rect 15654 18912 15660 18924
rect 15712 18912 15718 18964
rect 16209 18955 16267 18961
rect 16209 18921 16221 18955
rect 16255 18952 16267 18955
rect 16255 18924 16620 18952
rect 16255 18921 16267 18924
rect 16209 18915 16267 18921
rect 14737 18887 14795 18893
rect 11572 18856 12112 18884
rect 11572 18844 11578 18856
rect 12084 18828 12112 18856
rect 14737 18853 14749 18887
rect 14783 18853 14795 18887
rect 14737 18847 14795 18853
rect 15470 18844 15476 18896
rect 15528 18844 15534 18896
rect 16592 18893 16620 18924
rect 16577 18887 16635 18893
rect 16577 18853 16589 18887
rect 16623 18853 16635 18887
rect 16577 18847 16635 18853
rect 17034 18844 17040 18896
rect 17092 18844 17098 18896
rect 18138 18844 18144 18896
rect 18196 18884 18202 18896
rect 18509 18887 18567 18893
rect 18509 18884 18521 18887
rect 18196 18856 18521 18884
rect 18196 18844 18202 18856
rect 18509 18853 18521 18856
rect 18555 18853 18567 18887
rect 18509 18847 18567 18853
rect 11790 18825 11796 18828
rect 11425 18819 11483 18825
rect 11425 18816 11437 18819
rect 11348 18788 11437 18816
rect 10413 18779 10471 18785
rect 11425 18785 11437 18788
rect 11471 18785 11483 18819
rect 11425 18779 11483 18785
rect 11609 18819 11667 18825
rect 11609 18785 11621 18819
rect 11655 18785 11667 18819
rect 11609 18779 11667 18785
rect 11773 18819 11796 18825
rect 11773 18785 11785 18819
rect 11773 18779 11796 18785
rect 8570 18640 8576 18692
rect 8628 18680 8634 18692
rect 9122 18680 9128 18692
rect 8628 18652 9128 18680
rect 8628 18640 8634 18652
rect 9122 18640 9128 18652
rect 9180 18640 9186 18692
rect 11624 18680 11652 18779
rect 11790 18776 11796 18779
rect 11848 18776 11854 18828
rect 12066 18816 12072 18828
rect 11979 18788 12072 18816
rect 12066 18776 12072 18788
rect 12124 18776 12130 18828
rect 13633 18819 13691 18825
rect 13633 18785 13645 18819
rect 13679 18816 13691 18819
rect 14274 18816 14280 18828
rect 13679 18788 14280 18816
rect 13679 18785 13691 18788
rect 13633 18779 13691 18785
rect 14274 18776 14280 18788
rect 14332 18776 14338 18828
rect 18046 18776 18052 18828
rect 18104 18816 18110 18828
rect 18325 18819 18383 18825
rect 18325 18816 18337 18819
rect 18104 18788 18337 18816
rect 18104 18776 18110 18788
rect 18325 18785 18337 18788
rect 18371 18785 18383 18819
rect 18325 18779 18383 18785
rect 12710 18748 12716 18760
rect 12268 18720 12716 18748
rect 12268 18680 12296 18720
rect 12710 18708 12716 18720
rect 12768 18748 12774 18760
rect 13722 18748 13728 18760
rect 12768 18720 13728 18748
rect 12768 18708 12774 18720
rect 13722 18708 13728 18720
rect 13780 18708 13786 18760
rect 14461 18751 14519 18757
rect 14461 18717 14473 18751
rect 14507 18748 14519 18751
rect 16301 18751 16359 18757
rect 16301 18748 16313 18751
rect 14507 18720 16313 18748
rect 14507 18717 14519 18720
rect 14461 18711 14519 18717
rect 16301 18717 16313 18720
rect 16347 18748 16359 18751
rect 16942 18748 16948 18760
rect 16347 18720 16948 18748
rect 16347 18717 16359 18720
rect 16301 18711 16359 18717
rect 11624 18652 12296 18680
rect 12342 18640 12348 18692
rect 12400 18680 12406 18692
rect 12526 18680 12532 18692
rect 12400 18652 12532 18680
rect 12400 18640 12406 18652
rect 12526 18640 12532 18652
rect 12584 18640 12590 18692
rect 12618 18640 12624 18692
rect 12676 18680 12682 18692
rect 14476 18680 14504 18711
rect 16942 18708 16948 18720
rect 17000 18708 17006 18760
rect 18690 18680 18696 18692
rect 12676 18652 14504 18680
rect 18651 18652 18696 18680
rect 12676 18640 12682 18652
rect 13740 18624 13768 18652
rect 18690 18640 18696 18652
rect 18748 18640 18754 18692
rect 8846 18612 8852 18624
rect 8352 18584 8524 18612
rect 8807 18584 8852 18612
rect 8352 18572 8358 18584
rect 8846 18572 8852 18584
rect 8904 18572 8910 18624
rect 11698 18572 11704 18624
rect 11756 18612 11762 18624
rect 11977 18615 12035 18621
rect 11977 18612 11989 18615
rect 11756 18584 11989 18612
rect 11756 18572 11762 18584
rect 11977 18581 11989 18584
rect 12023 18581 12035 18615
rect 11977 18575 12035 18581
rect 13722 18572 13728 18624
rect 13780 18572 13786 18624
rect 17218 18572 17224 18624
rect 17276 18612 17282 18624
rect 18049 18615 18107 18621
rect 18049 18612 18061 18615
rect 17276 18584 18061 18612
rect 17276 18572 17282 18584
rect 18049 18581 18061 18584
rect 18095 18581 18107 18615
rect 18049 18575 18107 18581
rect 18141 18615 18199 18621
rect 18141 18581 18153 18615
rect 18187 18612 18199 18615
rect 18230 18612 18236 18624
rect 18187 18584 18236 18612
rect 18187 18581 18199 18584
rect 18141 18575 18199 18581
rect 18230 18572 18236 18584
rect 18288 18572 18294 18624
rect 1104 18522 19044 18544
rect 1104 18470 3972 18522
rect 4024 18470 4036 18522
rect 4088 18470 4100 18522
rect 4152 18470 4164 18522
rect 4216 18470 9952 18522
rect 10004 18470 10016 18522
rect 10068 18470 10080 18522
rect 10132 18470 10144 18522
rect 10196 18470 15932 18522
rect 15984 18470 15996 18522
rect 16048 18470 16060 18522
rect 16112 18470 16124 18522
rect 16176 18470 19044 18522
rect 1104 18448 19044 18470
rect 7742 18368 7748 18420
rect 7800 18408 7806 18420
rect 8205 18411 8263 18417
rect 8205 18408 8217 18411
rect 7800 18380 8217 18408
rect 7800 18368 7806 18380
rect 8205 18377 8217 18380
rect 8251 18377 8263 18411
rect 12802 18408 12808 18420
rect 12763 18380 12808 18408
rect 8205 18371 8263 18377
rect 6730 18272 6736 18284
rect 6691 18244 6736 18272
rect 6730 18232 6736 18244
rect 6788 18232 6794 18284
rect 8220 18272 8248 18371
rect 12802 18368 12808 18380
rect 12860 18368 12866 18420
rect 18693 18411 18751 18417
rect 18693 18377 18705 18411
rect 18739 18408 18751 18411
rect 19153 18411 19211 18417
rect 19153 18408 19165 18411
rect 18739 18380 19165 18408
rect 18739 18377 18751 18380
rect 18693 18371 18751 18377
rect 19153 18377 19165 18380
rect 19199 18377 19211 18411
rect 19153 18371 19211 18377
rect 11790 18340 11796 18352
rect 9646 18312 11796 18340
rect 9646 18272 9674 18312
rect 11790 18300 11796 18312
rect 11848 18300 11854 18352
rect 8220 18244 8524 18272
rect 4614 18164 4620 18216
rect 4672 18204 4678 18216
rect 4709 18207 4767 18213
rect 4709 18204 4721 18207
rect 4672 18176 4721 18204
rect 4672 18164 4678 18176
rect 4709 18173 4721 18176
rect 4755 18173 4767 18207
rect 4709 18167 4767 18173
rect 4798 18164 4804 18216
rect 4856 18204 4862 18216
rect 6454 18204 6460 18216
rect 4856 18176 6460 18204
rect 4856 18164 4862 18176
rect 6454 18164 6460 18176
rect 6512 18164 6518 18216
rect 8294 18204 8300 18216
rect 8255 18176 8300 18204
rect 8294 18164 8300 18176
rect 8352 18164 8358 18216
rect 8496 18213 8524 18244
rect 8864 18244 9674 18272
rect 8864 18213 8892 18244
rect 11514 18232 11520 18284
rect 11572 18272 11578 18284
rect 12621 18275 12679 18281
rect 12621 18272 12633 18275
rect 11572 18244 12633 18272
rect 11572 18232 11578 18244
rect 8481 18207 8539 18213
rect 8481 18173 8493 18207
rect 8527 18173 8539 18207
rect 8481 18167 8539 18173
rect 8849 18207 8907 18213
rect 8849 18173 8861 18207
rect 8895 18173 8907 18207
rect 9030 18204 9036 18216
rect 8991 18176 9036 18204
rect 8849 18167 8907 18173
rect 7282 18096 7288 18148
rect 7340 18096 7346 18148
rect 8202 18096 8208 18148
rect 8260 18136 8266 18148
rect 8864 18136 8892 18167
rect 9030 18164 9036 18176
rect 9088 18164 9094 18216
rect 9122 18164 9128 18216
rect 9180 18204 9186 18216
rect 11698 18204 11704 18216
rect 9180 18176 9225 18204
rect 11659 18176 11704 18204
rect 9180 18164 9186 18176
rect 11698 18164 11704 18176
rect 11756 18164 11762 18216
rect 11900 18213 11928 18244
rect 12621 18241 12633 18244
rect 12667 18272 12679 18275
rect 16942 18272 16948 18284
rect 12667 18244 13032 18272
rect 16903 18244 16948 18272
rect 12667 18241 12679 18244
rect 12621 18235 12679 18241
rect 11885 18207 11943 18213
rect 11885 18173 11897 18207
rect 11931 18173 11943 18207
rect 12066 18204 12072 18216
rect 12027 18176 12072 18204
rect 11885 18167 11943 18173
rect 12066 18164 12072 18176
rect 12124 18164 12130 18216
rect 12710 18204 12716 18216
rect 12406 18176 12716 18204
rect 8260 18108 8892 18136
rect 11977 18139 12035 18145
rect 8260 18096 8266 18108
rect 11977 18105 11989 18139
rect 12023 18136 12035 18139
rect 12406 18136 12434 18176
rect 12710 18164 12716 18176
rect 12768 18164 12774 18216
rect 13004 18213 13032 18244
rect 16942 18232 16948 18244
rect 17000 18232 17006 18284
rect 17218 18272 17224 18284
rect 17179 18244 17224 18272
rect 17218 18232 17224 18244
rect 17276 18232 17282 18284
rect 12989 18207 13047 18213
rect 12989 18173 13001 18207
rect 13035 18173 13047 18207
rect 12989 18167 13047 18173
rect 13081 18207 13139 18213
rect 13081 18173 13093 18207
rect 13127 18204 13139 18207
rect 13446 18204 13452 18216
rect 13127 18176 13452 18204
rect 13127 18173 13139 18176
rect 13081 18167 13139 18173
rect 13446 18164 13452 18176
rect 13504 18164 13510 18216
rect 12802 18136 12808 18148
rect 12023 18108 12434 18136
rect 12763 18108 12808 18136
rect 12023 18105 12035 18108
rect 11977 18099 12035 18105
rect 12802 18096 12808 18108
rect 12860 18096 12866 18148
rect 18230 18096 18236 18148
rect 18288 18096 18294 18148
rect 4338 18028 4344 18080
rect 4396 18068 4402 18080
rect 4801 18071 4859 18077
rect 4801 18068 4813 18071
rect 4396 18040 4813 18068
rect 4396 18028 4402 18040
rect 4801 18037 4813 18040
rect 4847 18037 4859 18071
rect 4801 18031 4859 18037
rect 7742 18028 7748 18080
rect 7800 18068 7806 18080
rect 9306 18068 9312 18080
rect 7800 18040 9312 18068
rect 7800 18028 7806 18040
rect 9306 18028 9312 18040
rect 9364 18028 9370 18080
rect 12250 18068 12256 18080
rect 12211 18040 12256 18068
rect 12250 18028 12256 18040
rect 12308 18028 12314 18080
rect 1104 17978 19044 18000
rect 1104 17926 6962 17978
rect 7014 17926 7026 17978
rect 7078 17926 7090 17978
rect 7142 17926 7154 17978
rect 7206 17926 12942 17978
rect 12994 17926 13006 17978
rect 13058 17926 13070 17978
rect 13122 17926 13134 17978
rect 13186 17926 19044 17978
rect 1104 17904 19044 17926
rect 6641 17867 6699 17873
rect 6641 17833 6653 17867
rect 6687 17864 6699 17867
rect 7282 17864 7288 17876
rect 6687 17836 7288 17864
rect 6687 17833 6699 17836
rect 6641 17827 6699 17833
rect 7282 17824 7288 17836
rect 7340 17824 7346 17876
rect 11790 17824 11796 17876
rect 11848 17864 11854 17876
rect 12802 17864 12808 17876
rect 11848 17836 12808 17864
rect 11848 17824 11854 17836
rect 12802 17824 12808 17836
rect 12860 17824 12866 17876
rect 4430 17796 4436 17808
rect 4391 17768 4436 17796
rect 4430 17756 4436 17768
rect 4488 17796 4494 17808
rect 4488 17768 4752 17796
rect 4488 17756 4494 17768
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 4614 17728 4620 17740
rect 4575 17700 4620 17728
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 4724 17737 4752 17768
rect 11072 17768 11928 17796
rect 4709 17731 4767 17737
rect 4709 17697 4721 17731
rect 4755 17697 4767 17731
rect 4709 17691 4767 17697
rect 4893 17731 4951 17737
rect 4893 17697 4905 17731
rect 4939 17697 4951 17731
rect 4893 17691 4951 17697
rect 6457 17731 6515 17737
rect 6457 17697 6469 17731
rect 6503 17728 6515 17731
rect 7374 17728 7380 17740
rect 6503 17700 7380 17728
rect 6503 17697 6515 17700
rect 6457 17691 6515 17697
rect 4632 17660 4660 17688
rect 4908 17660 4936 17691
rect 4632 17632 4936 17660
rect 3602 17552 3608 17604
rect 3660 17592 3666 17604
rect 6472 17592 6500 17691
rect 7374 17688 7380 17700
rect 7432 17728 7438 17740
rect 7742 17728 7748 17740
rect 7432 17700 7748 17728
rect 7432 17688 7438 17700
rect 7742 17688 7748 17700
rect 7800 17688 7806 17740
rect 11072 17737 11100 17768
rect 11900 17740 11928 17768
rect 12526 17756 12532 17808
rect 12584 17796 12590 17808
rect 12584 17768 13216 17796
rect 12584 17756 12590 17768
rect 13188 17740 13216 17768
rect 13262 17756 13268 17808
rect 13320 17796 13326 17808
rect 14918 17796 14924 17808
rect 13320 17768 14924 17796
rect 13320 17756 13326 17768
rect 11057 17731 11115 17737
rect 11057 17697 11069 17731
rect 11103 17697 11115 17731
rect 11057 17691 11115 17697
rect 11241 17731 11299 17737
rect 11241 17697 11253 17731
rect 11287 17697 11299 17731
rect 11514 17728 11520 17740
rect 11475 17700 11520 17728
rect 11241 17691 11299 17697
rect 11256 17660 11284 17691
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 11698 17728 11704 17740
rect 11659 17700 11704 17728
rect 11698 17688 11704 17700
rect 11756 17688 11762 17740
rect 11882 17728 11888 17740
rect 11843 17700 11888 17728
rect 11882 17688 11888 17700
rect 11940 17688 11946 17740
rect 12066 17728 12072 17740
rect 12027 17700 12072 17728
rect 12066 17688 12072 17700
rect 12124 17728 12130 17740
rect 12805 17731 12863 17737
rect 12805 17728 12817 17731
rect 12124 17700 12817 17728
rect 12124 17688 12130 17700
rect 12805 17697 12817 17700
rect 12851 17697 12863 17731
rect 13170 17728 13176 17740
rect 13131 17700 13176 17728
rect 12805 17691 12863 17697
rect 13170 17688 13176 17700
rect 13228 17688 13234 17740
rect 13357 17731 13415 17737
rect 13357 17728 13369 17731
rect 13280 17700 13369 17728
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 11256 17632 11805 17660
rect 11793 17629 11805 17632
rect 11839 17660 11851 17663
rect 12161 17663 12219 17669
rect 12161 17660 12173 17663
rect 11839 17632 12173 17660
rect 11839 17629 11851 17632
rect 11793 17623 11851 17629
rect 12161 17629 12173 17632
rect 12207 17629 12219 17663
rect 12342 17660 12348 17672
rect 12303 17632 12348 17660
rect 12161 17623 12219 17629
rect 12342 17620 12348 17632
rect 12400 17620 12406 17672
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17629 12495 17663
rect 12437 17623 12495 17629
rect 3660 17564 6500 17592
rect 3660 17552 3666 17564
rect 9674 17552 9680 17604
rect 9732 17592 9738 17604
rect 9732 17564 11284 17592
rect 9732 17552 9738 17564
rect 11256 17536 11284 17564
rect 12250 17552 12256 17604
rect 12308 17592 12314 17604
rect 12452 17592 12480 17623
rect 12710 17620 12716 17672
rect 12768 17660 12774 17672
rect 13280 17660 13308 17700
rect 13357 17697 13369 17700
rect 13403 17697 13415 17731
rect 13357 17691 13415 17697
rect 13446 17688 13452 17740
rect 13504 17728 13510 17740
rect 13740 17737 13768 17768
rect 14918 17756 14924 17768
rect 14976 17756 14982 17808
rect 13725 17731 13783 17737
rect 13504 17700 13549 17728
rect 13504 17688 13510 17700
rect 13725 17697 13737 17731
rect 13771 17697 13783 17731
rect 13725 17691 13783 17697
rect 14274 17688 14280 17740
rect 14332 17728 14338 17740
rect 14553 17731 14611 17737
rect 14553 17728 14565 17731
rect 14332 17700 14565 17728
rect 14332 17688 14338 17700
rect 14553 17697 14565 17700
rect 14599 17728 14611 17731
rect 15010 17728 15016 17740
rect 14599 17700 15016 17728
rect 14599 17697 14611 17700
rect 14553 17691 14611 17697
rect 15010 17688 15016 17700
rect 15068 17688 15074 17740
rect 12768 17632 13308 17660
rect 12768 17620 12774 17632
rect 12308 17564 12480 17592
rect 12308 17552 12314 17564
rect 1581 17527 1639 17533
rect 1581 17493 1593 17527
rect 1627 17524 1639 17527
rect 1670 17524 1676 17536
rect 1627 17496 1676 17524
rect 1627 17493 1639 17496
rect 1581 17487 1639 17493
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 3786 17484 3792 17536
rect 3844 17524 3850 17536
rect 4249 17527 4307 17533
rect 4249 17524 4261 17527
rect 3844 17496 4261 17524
rect 3844 17484 3850 17496
rect 4249 17493 4261 17496
rect 4295 17493 4307 17527
rect 4798 17524 4804 17536
rect 4759 17496 4804 17524
rect 4249 17487 4307 17493
rect 4798 17484 4804 17496
rect 4856 17484 4862 17536
rect 10318 17484 10324 17536
rect 10376 17524 10382 17536
rect 11149 17527 11207 17533
rect 11149 17524 11161 17527
rect 10376 17496 11161 17524
rect 10376 17484 10382 17496
rect 11149 17493 11161 17496
rect 11195 17493 11207 17527
rect 11149 17487 11207 17493
rect 11238 17484 11244 17536
rect 11296 17524 11302 17536
rect 11333 17527 11391 17533
rect 11333 17524 11345 17527
rect 11296 17496 11345 17524
rect 11296 17484 11302 17496
rect 11333 17493 11345 17496
rect 11379 17493 11391 17527
rect 11333 17487 11391 17493
rect 11698 17484 11704 17536
rect 11756 17524 11762 17536
rect 12342 17524 12348 17536
rect 11756 17496 12348 17524
rect 11756 17484 11762 17496
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 13280 17524 13308 17632
rect 13541 17663 13599 17669
rect 13541 17629 13553 17663
rect 13587 17660 13599 17663
rect 14642 17660 14648 17672
rect 13587 17632 14648 17660
rect 13587 17629 13599 17632
rect 13541 17623 13599 17629
rect 13354 17552 13360 17604
rect 13412 17592 13418 17604
rect 13556 17592 13584 17623
rect 14642 17620 14648 17632
rect 14700 17620 14706 17672
rect 13412 17564 13584 17592
rect 13412 17552 13418 17564
rect 13538 17524 13544 17536
rect 13280 17496 13544 17524
rect 13538 17484 13544 17496
rect 13596 17484 13602 17536
rect 13814 17484 13820 17536
rect 13872 17524 13878 17536
rect 13909 17527 13967 17533
rect 13909 17524 13921 17527
rect 13872 17496 13921 17524
rect 13872 17484 13878 17496
rect 13909 17493 13921 17496
rect 13955 17493 13967 17527
rect 13909 17487 13967 17493
rect 14737 17527 14795 17533
rect 14737 17493 14749 17527
rect 14783 17524 14795 17527
rect 14826 17524 14832 17536
rect 14783 17496 14832 17524
rect 14783 17493 14795 17496
rect 14737 17487 14795 17493
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 1104 17434 19044 17456
rect 1104 17382 3972 17434
rect 4024 17382 4036 17434
rect 4088 17382 4100 17434
rect 4152 17382 4164 17434
rect 4216 17382 9952 17434
rect 10004 17382 10016 17434
rect 10068 17382 10080 17434
rect 10132 17382 10144 17434
rect 10196 17382 15932 17434
rect 15984 17382 15996 17434
rect 16048 17382 16060 17434
rect 16112 17382 16124 17434
rect 16176 17382 19044 17434
rect 1104 17360 19044 17382
rect 4433 17323 4491 17329
rect 4433 17289 4445 17323
rect 4479 17320 4491 17323
rect 4614 17320 4620 17332
rect 4479 17292 4620 17320
rect 4479 17289 4491 17292
rect 4433 17283 4491 17289
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 12066 17320 12072 17332
rect 10060 17292 11468 17320
rect 12027 17292 12072 17320
rect 3329 17255 3387 17261
rect 3329 17221 3341 17255
rect 3375 17252 3387 17255
rect 10060 17252 10088 17292
rect 3375 17224 4200 17252
rect 3375 17221 3387 17224
rect 3329 17215 3387 17221
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17184 1915 17187
rect 3697 17187 3755 17193
rect 3697 17184 3709 17187
rect 1903 17156 3709 17184
rect 1903 17153 1915 17156
rect 1857 17147 1915 17153
rect 3697 17153 3709 17156
rect 3743 17153 3755 17187
rect 3697 17147 3755 17153
rect 4172 17184 4200 17224
rect 9968 17224 10088 17252
rect 10321 17255 10379 17261
rect 4890 17184 4896 17196
rect 4172 17156 4660 17184
rect 4851 17156 4896 17184
rect 1581 17119 1639 17125
rect 1581 17085 1593 17119
rect 1627 17085 1639 17119
rect 3602 17116 3608 17128
rect 3563 17088 3608 17116
rect 1581 17079 1639 17085
rect 1596 17048 1624 17079
rect 3602 17076 3608 17088
rect 3660 17076 3666 17128
rect 3786 17076 3792 17128
rect 3844 17116 3850 17128
rect 4172 17125 4200 17156
rect 3881 17119 3939 17125
rect 3881 17116 3893 17119
rect 3844 17088 3893 17116
rect 3844 17076 3850 17088
rect 3881 17085 3893 17088
rect 3927 17085 3939 17119
rect 4172 17119 4241 17125
rect 4172 17088 4195 17119
rect 3881 17079 3939 17085
rect 4183 17085 4195 17088
rect 4229 17085 4241 17119
rect 4183 17079 4241 17085
rect 4341 17119 4399 17125
rect 4341 17085 4353 17119
rect 4387 17116 4399 17119
rect 4522 17116 4528 17128
rect 4387 17088 4528 17116
rect 4387 17085 4399 17088
rect 4341 17079 4399 17085
rect 4522 17076 4528 17088
rect 4580 17076 4586 17128
rect 4632 17125 4660 17156
rect 4890 17144 4896 17156
rect 4948 17144 4954 17196
rect 5169 17187 5227 17193
rect 5169 17184 5181 17187
rect 5000 17156 5181 17184
rect 5000 17128 5028 17156
rect 5169 17153 5181 17156
rect 5215 17153 5227 17187
rect 9674 17184 9680 17196
rect 9635 17156 9680 17184
rect 5169 17147 5227 17153
rect 9674 17144 9680 17156
rect 9732 17144 9738 17196
rect 9766 17144 9772 17196
rect 9824 17184 9830 17196
rect 9968 17193 9996 17224
rect 10321 17221 10333 17255
rect 10367 17252 10379 17255
rect 11330 17252 11336 17264
rect 10367 17224 11336 17252
rect 10367 17221 10379 17224
rect 10321 17215 10379 17221
rect 11330 17212 11336 17224
rect 11388 17212 11394 17264
rect 11440 17252 11468 17292
rect 12066 17280 12072 17292
rect 12124 17280 12130 17332
rect 13078 17280 13084 17332
rect 13136 17320 13142 17332
rect 13262 17320 13268 17332
rect 13136 17292 13268 17320
rect 13136 17280 13142 17292
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 13357 17323 13415 17329
rect 13357 17289 13369 17323
rect 13403 17320 13415 17323
rect 13446 17320 13452 17332
rect 13403 17292 13452 17320
rect 13403 17289 13415 17292
rect 13357 17283 13415 17289
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 16025 17323 16083 17329
rect 16025 17320 16037 17323
rect 13648 17292 16037 17320
rect 13648 17252 13676 17292
rect 16025 17289 16037 17292
rect 16071 17289 16083 17323
rect 16025 17283 16083 17289
rect 11440 17224 13676 17252
rect 14918 17212 14924 17264
rect 14976 17252 14982 17264
rect 15289 17255 15347 17261
rect 15289 17252 15301 17255
rect 14976 17224 15301 17252
rect 14976 17212 14982 17224
rect 15289 17221 15301 17224
rect 15335 17221 15347 17255
rect 15289 17215 15347 17221
rect 9861 17187 9919 17193
rect 9861 17184 9873 17187
rect 9824 17156 9873 17184
rect 9824 17144 9830 17156
rect 9861 17153 9873 17156
rect 9907 17153 9919 17187
rect 9861 17147 9919 17153
rect 9953 17187 10011 17193
rect 9953 17153 9965 17187
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 10137 17187 10195 17193
rect 10137 17153 10149 17187
rect 10183 17153 10195 17187
rect 15841 17187 15899 17193
rect 15841 17184 15853 17187
rect 10137 17147 10195 17153
rect 13004 17156 15853 17184
rect 4617 17119 4675 17125
rect 4617 17085 4629 17119
rect 4663 17085 4675 17119
rect 4617 17079 4675 17085
rect 1854 17048 1860 17060
rect 1596 17020 1860 17048
rect 1854 17008 1860 17020
rect 1912 17008 1918 17060
rect 3973 17051 4031 17057
rect 3082 17020 3464 17048
rect 3436 16989 3464 17020
rect 3973 17017 3985 17051
rect 4019 17017 4031 17051
rect 3973 17011 4031 17017
rect 4065 17051 4123 17057
rect 4065 17017 4077 17051
rect 4111 17048 4123 17051
rect 4430 17048 4436 17060
rect 4111 17020 4436 17048
rect 4111 17017 4123 17020
rect 4065 17011 4123 17017
rect 3421 16983 3479 16989
rect 3421 16949 3433 16983
rect 3467 16949 3479 16983
rect 3988 16980 4016 17011
rect 4430 17008 4436 17020
rect 4488 17008 4494 17060
rect 4632 17048 4660 17079
rect 4706 17076 4712 17128
rect 4764 17116 4770 17128
rect 4982 17116 4988 17128
rect 4764 17088 4809 17116
rect 4895 17088 4988 17116
rect 4764 17076 4770 17088
rect 4982 17076 4988 17088
rect 5040 17076 5046 17128
rect 5077 17119 5135 17125
rect 5077 17085 5089 17119
rect 5123 17085 5135 17119
rect 5077 17079 5135 17085
rect 7377 17119 7435 17125
rect 7377 17085 7389 17119
rect 7423 17116 7435 17119
rect 7742 17116 7748 17128
rect 7423 17088 7748 17116
rect 7423 17085 7435 17088
rect 7377 17079 7435 17085
rect 5092 17048 5120 17079
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 9030 17076 9036 17128
rect 9088 17116 9094 17128
rect 9585 17119 9643 17125
rect 9585 17116 9597 17119
rect 9088 17088 9597 17116
rect 9088 17076 9094 17088
rect 9585 17085 9597 17088
rect 9631 17085 9643 17119
rect 9876 17116 9904 17147
rect 10152 17116 10180 17147
rect 9876 17088 10180 17116
rect 10413 17119 10471 17125
rect 9585 17079 9643 17085
rect 10413 17085 10425 17119
rect 10459 17116 10471 17119
rect 10594 17116 10600 17128
rect 10459 17088 10600 17116
rect 10459 17085 10471 17088
rect 10413 17079 10471 17085
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 10689 17119 10747 17125
rect 10689 17085 10701 17119
rect 10735 17116 10747 17119
rect 11238 17116 11244 17128
rect 10735 17088 11244 17116
rect 10735 17085 10747 17088
rect 10689 17079 10747 17085
rect 11238 17076 11244 17088
rect 11296 17076 11302 17128
rect 11330 17076 11336 17128
rect 11388 17116 11394 17128
rect 13004 17116 13032 17156
rect 15841 17153 15853 17156
rect 15887 17184 15899 17187
rect 16390 17184 16396 17196
rect 15887 17156 16396 17184
rect 15887 17153 15899 17156
rect 15841 17147 15899 17153
rect 16390 17144 16396 17156
rect 16448 17144 16454 17196
rect 17218 17184 17224 17196
rect 16500 17156 17224 17184
rect 11388 17088 13032 17116
rect 11388 17076 11394 17088
rect 13078 17076 13084 17128
rect 13136 17116 13142 17128
rect 13265 17119 13323 17125
rect 13265 17116 13277 17119
rect 13136 17088 13277 17116
rect 13136 17076 13142 17088
rect 13265 17085 13277 17088
rect 13311 17085 13323 17119
rect 13265 17079 13323 17085
rect 13354 17076 13360 17128
rect 13412 17116 13418 17128
rect 13449 17119 13507 17125
rect 13449 17116 13461 17119
rect 13412 17088 13461 17116
rect 13412 17076 13418 17088
rect 13449 17085 13461 17088
rect 13495 17085 13507 17119
rect 13449 17079 13507 17085
rect 13541 17119 13599 17125
rect 13541 17085 13553 17119
rect 13587 17085 13599 17119
rect 13541 17079 13599 17085
rect 16301 17119 16359 17125
rect 16301 17085 16313 17119
rect 16347 17116 16359 17119
rect 16500 17116 16528 17156
rect 17218 17144 17224 17156
rect 17276 17144 17282 17196
rect 16347 17088 16528 17116
rect 16577 17119 16635 17125
rect 16347 17085 16359 17088
rect 16301 17079 16359 17085
rect 16577 17085 16589 17119
rect 16623 17085 16635 17119
rect 16577 17079 16635 17085
rect 4632 17020 5120 17048
rect 8110 17008 8116 17060
rect 8168 17048 8174 17060
rect 9401 17051 9459 17057
rect 9401 17048 9413 17051
rect 8168 17020 9413 17048
rect 8168 17008 8174 17020
rect 9401 17017 9413 17020
rect 9447 17017 9459 17051
rect 10042 17048 10048 17060
rect 10003 17020 10048 17048
rect 9401 17011 9459 17017
rect 10042 17008 10048 17020
rect 10100 17008 10106 17060
rect 10137 17051 10195 17057
rect 10137 17017 10149 17051
rect 10183 17048 10195 17051
rect 10778 17048 10784 17060
rect 10183 17020 10784 17048
rect 10183 17017 10195 17020
rect 10137 17011 10195 17017
rect 10778 17008 10784 17020
rect 10836 17008 10842 17060
rect 11698 17048 11704 17060
rect 11659 17020 11704 17048
rect 11698 17008 11704 17020
rect 11756 17008 11762 17060
rect 11885 17051 11943 17057
rect 11885 17017 11897 17051
rect 11931 17048 11943 17051
rect 12250 17048 12256 17060
rect 11931 17020 12256 17048
rect 11931 17017 11943 17020
rect 11885 17011 11943 17017
rect 12250 17008 12256 17020
rect 12308 17008 12314 17060
rect 13556 17048 13584 17079
rect 13722 17048 13728 17060
rect 13556 17020 13728 17048
rect 13722 17008 13728 17020
rect 13780 17008 13786 17060
rect 13814 17008 13820 17060
rect 13872 17048 13878 17060
rect 13872 17020 13917 17048
rect 13872 17008 13878 17020
rect 14826 17008 14832 17060
rect 14884 17008 14890 17060
rect 16485 17051 16543 17057
rect 16485 17048 16497 17051
rect 15120 17020 16497 17048
rect 4798 16980 4804 16992
rect 3988 16952 4804 16980
rect 3421 16943 3479 16949
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 7558 16980 7564 16992
rect 7519 16952 7564 16980
rect 7558 16940 7564 16952
rect 7616 16940 7622 16992
rect 9950 16940 9956 16992
rect 10008 16980 10014 16992
rect 10597 16983 10655 16989
rect 10597 16980 10609 16983
rect 10008 16952 10609 16980
rect 10008 16940 10014 16952
rect 10597 16949 10609 16952
rect 10643 16949 10655 16983
rect 10597 16943 10655 16949
rect 10686 16940 10692 16992
rect 10744 16980 10750 16992
rect 15120 16980 15148 17020
rect 16485 17017 16497 17020
rect 16531 17017 16543 17051
rect 16592 17048 16620 17079
rect 16758 17076 16764 17128
rect 16816 17116 16822 17128
rect 16945 17119 17003 17125
rect 16945 17116 16957 17119
rect 16816 17088 16957 17116
rect 16816 17076 16822 17088
rect 16945 17085 16957 17088
rect 16991 17085 17003 17119
rect 16945 17079 17003 17085
rect 17129 17119 17187 17125
rect 17129 17085 17141 17119
rect 17175 17116 17187 17119
rect 17494 17116 17500 17128
rect 17175 17088 17500 17116
rect 17175 17085 17187 17088
rect 17129 17079 17187 17085
rect 17034 17048 17040 17060
rect 16592 17020 17040 17048
rect 16485 17011 16543 17017
rect 17034 17008 17040 17020
rect 17092 17008 17098 17060
rect 10744 16952 15148 16980
rect 16209 16983 16267 16989
rect 10744 16940 10750 16952
rect 16209 16949 16221 16983
rect 16255 16980 16267 16983
rect 16574 16980 16580 16992
rect 16255 16952 16580 16980
rect 16255 16949 16267 16952
rect 16209 16943 16267 16949
rect 16574 16940 16580 16952
rect 16632 16940 16638 16992
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 17144 16980 17172 17079
rect 17494 17076 17500 17088
rect 17552 17076 17558 17128
rect 16724 16952 17172 16980
rect 16724 16940 16730 16952
rect 1104 16890 19044 16912
rect 1104 16838 6962 16890
rect 7014 16838 7026 16890
rect 7078 16838 7090 16890
rect 7142 16838 7154 16890
rect 7206 16838 12942 16890
rect 12994 16838 13006 16890
rect 13058 16838 13070 16890
rect 13122 16838 13134 16890
rect 13186 16838 19044 16890
rect 1104 16816 19044 16838
rect 4706 16736 4712 16788
rect 4764 16776 4770 16788
rect 5813 16779 5871 16785
rect 5813 16776 5825 16779
rect 4764 16748 5825 16776
rect 4764 16736 4770 16748
rect 5813 16745 5825 16748
rect 5859 16745 5871 16779
rect 16390 16776 16396 16788
rect 16351 16748 16396 16776
rect 5813 16739 5871 16745
rect 16390 16736 16396 16748
rect 16448 16736 16454 16788
rect 16574 16736 16580 16788
rect 16632 16776 16638 16788
rect 18506 16776 18512 16788
rect 16632 16748 18512 16776
rect 16632 16736 16638 16748
rect 7558 16668 7564 16720
rect 7616 16668 7622 16720
rect 16666 16708 16672 16720
rect 16592 16680 16672 16708
rect 4798 16640 4804 16652
rect 4724 16612 4804 16640
rect 4724 16581 4752 16612
rect 4798 16600 4804 16612
rect 4856 16600 4862 16652
rect 4982 16640 4988 16652
rect 4943 16612 4988 16640
rect 4982 16600 4988 16612
rect 5040 16600 5046 16652
rect 5721 16643 5779 16649
rect 5721 16609 5733 16643
rect 5767 16640 5779 16643
rect 5902 16640 5908 16652
rect 5767 16612 5908 16640
rect 5767 16609 5779 16612
rect 5721 16603 5779 16609
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16541 4767 16575
rect 4890 16572 4896 16584
rect 4803 16544 4896 16572
rect 4709 16535 4767 16541
rect 4890 16532 4896 16544
rect 4948 16572 4954 16584
rect 5736 16572 5764 16603
rect 5902 16600 5908 16612
rect 5960 16600 5966 16652
rect 9950 16640 9956 16652
rect 9911 16612 9956 16640
rect 9950 16600 9956 16612
rect 10008 16600 10014 16652
rect 10226 16640 10232 16652
rect 10187 16612 10232 16640
rect 10226 16600 10232 16612
rect 10284 16600 10290 16652
rect 10410 16640 10416 16652
rect 10371 16612 10416 16640
rect 10410 16600 10416 16612
rect 10468 16600 10474 16652
rect 10594 16640 10600 16652
rect 10555 16612 10600 16640
rect 10594 16600 10600 16612
rect 10652 16600 10658 16652
rect 10778 16640 10784 16652
rect 10739 16612 10784 16640
rect 10778 16600 10784 16612
rect 10836 16600 10842 16652
rect 16592 16649 16620 16680
rect 16666 16668 16672 16680
rect 16724 16668 16730 16720
rect 16577 16643 16635 16649
rect 16577 16609 16589 16643
rect 16623 16609 16635 16643
rect 16758 16640 16764 16652
rect 16719 16612 16764 16640
rect 16577 16603 16635 16609
rect 16758 16600 16764 16612
rect 16816 16600 16822 16652
rect 16960 16649 16988 16748
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 16945 16643 17003 16649
rect 16945 16609 16957 16643
rect 16991 16609 17003 16643
rect 16945 16603 17003 16609
rect 17034 16600 17040 16652
rect 17092 16640 17098 16652
rect 17129 16643 17187 16649
rect 17129 16640 17141 16643
rect 17092 16612 17141 16640
rect 17092 16600 17098 16612
rect 17129 16609 17141 16612
rect 17175 16609 17187 16643
rect 17129 16603 17187 16609
rect 18046 16600 18052 16652
rect 18104 16640 18110 16652
rect 18233 16643 18291 16649
rect 18233 16640 18245 16643
rect 18104 16612 18245 16640
rect 18104 16600 18110 16612
rect 18233 16609 18245 16612
rect 18279 16609 18291 16643
rect 18233 16603 18291 16609
rect 6546 16572 6552 16584
rect 4948 16544 5764 16572
rect 6507 16544 6552 16572
rect 4948 16532 4954 16544
rect 6546 16532 6552 16544
rect 6604 16532 6610 16584
rect 6825 16575 6883 16581
rect 6825 16541 6837 16575
rect 6871 16572 6883 16575
rect 6914 16572 6920 16584
rect 6871 16544 6920 16572
rect 6871 16541 6883 16544
rect 6825 16535 6883 16541
rect 6914 16532 6920 16544
rect 6972 16532 6978 16584
rect 9398 16532 9404 16584
rect 9456 16572 9462 16584
rect 9493 16575 9551 16581
rect 9493 16572 9505 16575
rect 9456 16544 9505 16572
rect 9456 16532 9462 16544
rect 9493 16541 9505 16544
rect 9539 16541 9551 16575
rect 9493 16535 9551 16541
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16572 16911 16575
rect 17218 16572 17224 16584
rect 16899 16544 17224 16572
rect 16899 16541 16911 16544
rect 16853 16535 16911 16541
rect 17218 16532 17224 16544
rect 17276 16532 17282 16584
rect 4798 16436 4804 16448
rect 4759 16408 4804 16436
rect 4798 16396 4804 16408
rect 4856 16396 4862 16448
rect 8294 16436 8300 16448
rect 8255 16408 8300 16436
rect 8294 16396 8300 16408
rect 8352 16396 8358 16448
rect 17954 16396 17960 16448
rect 18012 16436 18018 16448
rect 18049 16439 18107 16445
rect 18049 16436 18061 16439
rect 18012 16408 18061 16436
rect 18012 16396 18018 16408
rect 18049 16405 18061 16408
rect 18095 16405 18107 16439
rect 18049 16399 18107 16405
rect 1104 16346 19044 16368
rect 1104 16294 3972 16346
rect 4024 16294 4036 16346
rect 4088 16294 4100 16346
rect 4152 16294 4164 16346
rect 4216 16294 9952 16346
rect 10004 16294 10016 16346
rect 10068 16294 10080 16346
rect 10132 16294 10144 16346
rect 10196 16294 15932 16346
rect 15984 16294 15996 16346
rect 16048 16294 16060 16346
rect 16112 16294 16124 16346
rect 16176 16294 19044 16346
rect 1104 16272 19044 16294
rect 6914 16232 6920 16244
rect 6875 16204 6920 16232
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 10505 16235 10563 16241
rect 10505 16201 10517 16235
rect 10551 16201 10563 16235
rect 10505 16195 10563 16201
rect 4522 16124 4528 16176
rect 4580 16164 4586 16176
rect 8110 16164 8116 16176
rect 4580 16136 8116 16164
rect 4580 16124 4586 16136
rect 7466 16096 7472 16108
rect 7116 16068 7472 16096
rect 2777 16031 2835 16037
rect 2777 15997 2789 16031
rect 2823 16028 2835 16031
rect 3602 16028 3608 16040
rect 2823 16000 3608 16028
rect 2823 15997 2835 16000
rect 2777 15991 2835 15997
rect 3602 15988 3608 16000
rect 3660 15988 3666 16040
rect 7116 16037 7144 16068
rect 7466 16056 7472 16068
rect 7524 16056 7530 16108
rect 7576 16105 7604 16136
rect 8110 16124 8116 16136
rect 8168 16124 8174 16176
rect 9674 16164 9680 16176
rect 9232 16136 9680 16164
rect 9232 16105 9260 16136
rect 9674 16124 9680 16136
rect 9732 16164 9738 16176
rect 10318 16164 10324 16176
rect 9732 16136 10324 16164
rect 9732 16124 9738 16136
rect 10318 16124 10324 16136
rect 10376 16124 10382 16176
rect 10520 16164 10548 16195
rect 10594 16192 10600 16244
rect 10652 16232 10658 16244
rect 10689 16235 10747 16241
rect 10689 16232 10701 16235
rect 10652 16204 10701 16232
rect 10652 16192 10658 16204
rect 10689 16201 10701 16204
rect 10735 16201 10747 16235
rect 10689 16195 10747 16201
rect 10873 16167 10931 16173
rect 10873 16164 10885 16167
rect 10520 16136 10885 16164
rect 7561 16099 7619 16105
rect 7561 16065 7573 16099
rect 7607 16065 7619 16099
rect 7561 16059 7619 16065
rect 9217 16099 9275 16105
rect 9217 16065 9229 16099
rect 9263 16065 9275 16099
rect 9217 16059 9275 16065
rect 9769 16099 9827 16105
rect 9769 16065 9781 16099
rect 9815 16096 9827 16099
rect 9953 16099 10011 16105
rect 9815 16068 9904 16096
rect 9815 16065 9827 16068
rect 9769 16059 9827 16065
rect 7101 16031 7159 16037
rect 7101 15997 7113 16031
rect 7147 15997 7159 16031
rect 7101 15991 7159 15997
rect 7190 15988 7196 16040
rect 7248 16028 7254 16040
rect 7248 16000 7293 16028
rect 7248 15988 7254 16000
rect 9582 15988 9588 16040
rect 9640 16028 9646 16040
rect 9677 16031 9735 16037
rect 9677 16028 9689 16031
rect 9640 16000 9689 16028
rect 9640 15988 9646 16000
rect 9677 15997 9689 16000
rect 9723 15997 9735 16031
rect 9677 15991 9735 15997
rect 4246 15920 4252 15972
rect 4304 15960 4310 15972
rect 4430 15960 4436 15972
rect 4304 15932 4436 15960
rect 4304 15920 4310 15932
rect 4430 15920 4436 15932
rect 4488 15960 4494 15972
rect 5166 15960 5172 15972
rect 4488 15932 5172 15960
rect 4488 15920 4494 15932
rect 5166 15920 5172 15932
rect 5224 15960 5230 15972
rect 7285 15963 7343 15969
rect 7285 15960 7297 15963
rect 5224 15932 7297 15960
rect 5224 15920 5230 15932
rect 7285 15929 7297 15932
rect 7331 15929 7343 15963
rect 7285 15923 7343 15929
rect 7423 15963 7481 15969
rect 7423 15929 7435 15963
rect 7469 15960 7481 15963
rect 8294 15960 8300 15972
rect 7469 15932 8300 15960
rect 7469 15929 7481 15932
rect 7423 15923 7481 15929
rect 8294 15920 8300 15932
rect 8352 15920 8358 15972
rect 9401 15963 9459 15969
rect 9401 15929 9413 15963
rect 9447 15960 9459 15963
rect 9766 15960 9772 15972
rect 9447 15932 9772 15960
rect 9447 15929 9459 15932
rect 9401 15923 9459 15929
rect 9766 15920 9772 15932
rect 9824 15920 9830 15972
rect 2866 15852 2872 15904
rect 2924 15892 2930 15904
rect 2961 15895 3019 15901
rect 2961 15892 2973 15895
rect 2924 15864 2973 15892
rect 2924 15852 2930 15864
rect 2961 15861 2973 15864
rect 3007 15861 3019 15895
rect 9876 15892 9904 16068
rect 9953 16065 9965 16099
rect 9999 16096 10011 16099
rect 10520 16096 10548 16136
rect 10873 16133 10885 16136
rect 10919 16133 10931 16167
rect 10873 16127 10931 16133
rect 13722 16124 13728 16176
rect 13780 16164 13786 16176
rect 13780 16136 16988 16164
rect 13780 16124 13786 16136
rect 12802 16096 12808 16108
rect 9999 16068 10548 16096
rect 11992 16068 12808 16096
rect 9999 16065 10011 16068
rect 9953 16059 10011 16065
rect 11992 16040 12020 16068
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 16390 16096 16396 16108
rect 14844 16068 16396 16096
rect 10042 16028 10048 16040
rect 10003 16000 10048 16028
rect 10042 15988 10048 16000
rect 10100 15988 10106 16040
rect 10318 16028 10324 16040
rect 10279 16000 10324 16028
rect 10318 15988 10324 16000
rect 10376 15988 10382 16040
rect 10413 16031 10471 16037
rect 10413 15997 10425 16031
rect 10459 15997 10471 16031
rect 10413 15991 10471 15997
rect 10965 16031 11023 16037
rect 10965 15997 10977 16031
rect 11011 16028 11023 16031
rect 11054 16028 11060 16040
rect 11011 16000 11060 16028
rect 11011 15997 11023 16000
rect 10965 15991 11023 15997
rect 10060 15960 10088 15988
rect 10428 15960 10456 15991
rect 10060 15932 10456 15960
rect 10980 15892 11008 15991
rect 11054 15988 11060 16000
rect 11112 15988 11118 16040
rect 11885 16031 11943 16037
rect 11885 15997 11897 16031
rect 11931 16028 11943 16031
rect 11974 16028 11980 16040
rect 11931 16000 11980 16028
rect 11931 15997 11943 16000
rect 11885 15991 11943 15997
rect 11974 15988 11980 16000
rect 12032 15988 12038 16040
rect 12253 16031 12311 16037
rect 12253 15997 12265 16031
rect 12299 16028 12311 16031
rect 13262 16028 13268 16040
rect 12299 16000 13268 16028
rect 12299 15997 12311 16000
rect 12253 15991 12311 15997
rect 13262 15988 13268 16000
rect 13320 15988 13326 16040
rect 13538 15988 13544 16040
rect 13596 16028 13602 16040
rect 14458 16028 14464 16040
rect 13596 16000 14464 16028
rect 13596 15988 13602 16000
rect 14458 15988 14464 16000
rect 14516 15988 14522 16040
rect 14844 16037 14872 16068
rect 16390 16056 16396 16068
rect 16448 16056 16454 16108
rect 16960 16105 16988 16136
rect 16945 16099 17003 16105
rect 16945 16065 16957 16099
rect 16991 16065 17003 16099
rect 16945 16059 17003 16065
rect 14829 16031 14887 16037
rect 14829 15997 14841 16031
rect 14875 15997 14887 16031
rect 14829 15991 14887 15997
rect 14921 16031 14979 16037
rect 14921 15997 14933 16031
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 12066 15960 12072 15972
rect 12027 15932 12072 15960
rect 12066 15920 12072 15932
rect 12124 15920 12130 15972
rect 12158 15920 12164 15972
rect 12216 15960 12222 15972
rect 14550 15960 14556 15972
rect 12216 15932 12261 15960
rect 14511 15932 14556 15960
rect 12216 15920 12222 15932
rect 14550 15920 14556 15932
rect 14608 15920 14614 15972
rect 14645 15963 14703 15969
rect 14645 15929 14657 15963
rect 14691 15960 14703 15963
rect 14936 15960 14964 15991
rect 15010 15988 15016 16040
rect 15068 16037 15074 16040
rect 15068 16028 15079 16037
rect 15068 16000 15113 16028
rect 15068 15991 15079 16000
rect 15068 15988 15074 15991
rect 16574 15960 16580 15972
rect 14691 15932 14872 15960
rect 14936 15932 16580 15960
rect 14691 15929 14703 15932
rect 14645 15923 14703 15929
rect 14844 15904 14872 15932
rect 16574 15920 16580 15932
rect 16632 15920 16638 15972
rect 17126 15920 17132 15972
rect 17184 15960 17190 15972
rect 17221 15963 17279 15969
rect 17221 15960 17233 15963
rect 17184 15932 17233 15960
rect 17184 15920 17190 15932
rect 17221 15929 17233 15932
rect 17267 15929 17279 15963
rect 17221 15923 17279 15929
rect 17954 15920 17960 15972
rect 18012 15920 18018 15972
rect 9876 15864 11008 15892
rect 12437 15895 12495 15901
rect 2961 15855 3019 15861
rect 12437 15861 12449 15895
rect 12483 15892 12495 15895
rect 13446 15892 13452 15904
rect 12483 15864 13452 15892
rect 12483 15861 12495 15864
rect 12437 15855 12495 15861
rect 13446 15852 13452 15864
rect 13504 15852 13510 15904
rect 14274 15892 14280 15904
rect 14235 15864 14280 15892
rect 14274 15852 14280 15864
rect 14332 15852 14338 15904
rect 14826 15852 14832 15904
rect 14884 15852 14890 15904
rect 15194 15892 15200 15904
rect 15155 15864 15200 15892
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 18693 15895 18751 15901
rect 18693 15861 18705 15895
rect 18739 15892 18751 15895
rect 18739 15864 19104 15892
rect 18739 15861 18751 15864
rect 18693 15855 18751 15861
rect 1104 15802 19044 15824
rect 1104 15750 6962 15802
rect 7014 15750 7026 15802
rect 7078 15750 7090 15802
rect 7142 15750 7154 15802
rect 7206 15750 12942 15802
rect 12994 15750 13006 15802
rect 13058 15750 13070 15802
rect 13122 15750 13134 15802
rect 13186 15750 19044 15802
rect 1104 15728 19044 15750
rect 7466 15688 7472 15700
rect 7427 15660 7472 15688
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 9585 15691 9643 15697
rect 9585 15657 9597 15691
rect 9631 15688 9643 15691
rect 10042 15688 10048 15700
rect 9631 15660 10048 15688
rect 9631 15657 9643 15660
rect 9585 15651 9643 15657
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 11701 15691 11759 15697
rect 11701 15657 11713 15691
rect 11747 15688 11759 15691
rect 11977 15691 12035 15697
rect 11977 15688 11989 15691
rect 11747 15660 11989 15688
rect 11747 15657 11759 15660
rect 11701 15651 11759 15657
rect 11977 15657 11989 15660
rect 12023 15688 12035 15691
rect 12158 15688 12164 15700
rect 12023 15660 12164 15688
rect 12023 15657 12035 15660
rect 11977 15651 12035 15657
rect 12158 15648 12164 15660
rect 12216 15648 12222 15700
rect 13262 15648 13268 15700
rect 13320 15688 13326 15700
rect 14918 15688 14924 15700
rect 13320 15660 14924 15688
rect 13320 15648 13326 15660
rect 14918 15648 14924 15660
rect 14976 15688 14982 15700
rect 16942 15688 16948 15700
rect 14976 15660 16948 15688
rect 14976 15648 14982 15660
rect 16942 15648 16948 15660
rect 17000 15648 17006 15700
rect 17126 15688 17132 15700
rect 17087 15660 17132 15688
rect 17126 15648 17132 15660
rect 17184 15648 17190 15700
rect 17218 15648 17224 15700
rect 17276 15688 17282 15700
rect 17276 15660 17321 15688
rect 17276 15648 17282 15660
rect 2866 15580 2872 15632
rect 2924 15580 2930 15632
rect 4617 15623 4675 15629
rect 4617 15620 4629 15623
rect 4080 15592 4629 15620
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 1854 15552 1860 15564
rect 1815 15524 1860 15552
rect 1854 15512 1860 15524
rect 1912 15512 1918 15564
rect 4080 15561 4108 15592
rect 4617 15589 4629 15592
rect 4663 15589 4675 15623
rect 4798 15620 4804 15632
rect 4759 15592 4804 15620
rect 4617 15583 4675 15589
rect 4798 15580 4804 15592
rect 4856 15620 4862 15632
rect 4856 15592 5212 15620
rect 4856 15580 4862 15592
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15521 4123 15555
rect 4065 15515 4123 15521
rect 4157 15555 4215 15561
rect 4157 15521 4169 15555
rect 4203 15521 4215 15555
rect 4157 15515 4215 15521
rect 2133 15487 2191 15493
rect 2133 15453 2145 15487
rect 2179 15484 2191 15487
rect 3881 15487 3939 15493
rect 3881 15484 3893 15487
rect 2179 15456 3893 15484
rect 2179 15453 2191 15456
rect 2133 15447 2191 15453
rect 3881 15453 3893 15456
rect 3927 15453 3939 15487
rect 3881 15447 3939 15453
rect 4172 15416 4200 15515
rect 4246 15512 4252 15564
rect 4304 15552 4310 15564
rect 4430 15561 4436 15564
rect 4387 15555 4436 15561
rect 4304 15524 4349 15552
rect 4304 15512 4310 15524
rect 4387 15521 4399 15555
rect 4433 15521 4436 15555
rect 4387 15515 4436 15521
rect 4430 15512 4436 15515
rect 4488 15512 4494 15564
rect 4522 15512 4528 15564
rect 4580 15552 4586 15564
rect 4982 15552 4988 15564
rect 4580 15524 4625 15552
rect 4943 15524 4988 15552
rect 4580 15512 4586 15524
rect 4982 15512 4988 15524
rect 5040 15512 5046 15564
rect 5184 15561 5212 15592
rect 12710 15580 12716 15632
rect 12768 15580 12774 15632
rect 13446 15620 13452 15632
rect 13407 15592 13452 15620
rect 13446 15580 13452 15592
rect 13504 15580 13510 15632
rect 14274 15580 14280 15632
rect 14332 15620 14338 15632
rect 14645 15623 14703 15629
rect 14645 15620 14657 15623
rect 14332 15592 14657 15620
rect 14332 15580 14338 15592
rect 14645 15589 14657 15592
rect 14691 15589 14703 15623
rect 14645 15583 14703 15589
rect 15194 15580 15200 15632
rect 15252 15580 15258 15632
rect 16853 15623 16911 15629
rect 16853 15589 16865 15623
rect 16899 15620 16911 15623
rect 19076 15620 19104 15864
rect 16899 15592 19104 15620
rect 16899 15589 16911 15592
rect 16853 15583 16911 15589
rect 5169 15555 5227 15561
rect 5169 15521 5181 15555
rect 5215 15521 5227 15555
rect 5169 15515 5227 15521
rect 5445 15555 5503 15561
rect 5445 15521 5457 15555
rect 5491 15521 5503 15555
rect 7466 15552 7472 15564
rect 7427 15524 7472 15552
rect 5445 15515 5503 15521
rect 5000 15484 5028 15512
rect 5460 15484 5488 15515
rect 7466 15512 7472 15524
rect 7524 15512 7530 15564
rect 7650 15552 7656 15564
rect 7611 15524 7656 15552
rect 7650 15512 7656 15524
rect 7708 15512 7714 15564
rect 9493 15555 9551 15561
rect 9493 15521 9505 15555
rect 9539 15552 9551 15555
rect 9582 15552 9588 15564
rect 9539 15524 9588 15552
rect 9539 15521 9551 15524
rect 9493 15515 9551 15521
rect 9582 15512 9588 15524
rect 9640 15512 9646 15564
rect 11760 15555 11818 15561
rect 11760 15521 11772 15555
rect 11806 15552 11818 15555
rect 12066 15552 12072 15564
rect 11806 15524 12072 15552
rect 11806 15521 11818 15524
rect 11760 15515 11818 15521
rect 12066 15512 12072 15524
rect 12124 15512 12130 15564
rect 16574 15552 16580 15564
rect 16535 15524 16580 15552
rect 16574 15512 16580 15524
rect 16632 15512 16638 15564
rect 16761 15555 16819 15561
rect 16761 15521 16773 15555
rect 16807 15521 16819 15555
rect 16942 15552 16948 15564
rect 16855 15524 16948 15552
rect 16761 15515 16819 15521
rect 5000 15456 5488 15484
rect 11241 15487 11299 15493
rect 11241 15453 11253 15487
rect 11287 15484 11299 15487
rect 11882 15484 11888 15496
rect 11287 15456 11888 15484
rect 11287 15453 11299 15456
rect 11241 15447 11299 15453
rect 11882 15444 11888 15456
rect 11940 15444 11946 15496
rect 13722 15484 13728 15496
rect 13683 15456 13728 15484
rect 13722 15444 13728 15456
rect 13780 15484 13786 15496
rect 14369 15487 14427 15493
rect 14369 15484 14381 15487
rect 13780 15456 14381 15484
rect 13780 15444 13786 15456
rect 14369 15453 14381 15456
rect 14415 15453 14427 15487
rect 16776 15484 16804 15515
rect 16942 15512 16948 15524
rect 17000 15552 17006 15564
rect 17218 15552 17224 15564
rect 17000 15524 17224 15552
rect 17000 15512 17006 15524
rect 17218 15512 17224 15524
rect 17276 15512 17282 15564
rect 17402 15552 17408 15564
rect 17363 15524 17408 15552
rect 17402 15512 17408 15524
rect 17460 15512 17466 15564
rect 17586 15552 17592 15564
rect 17547 15524 17592 15552
rect 17586 15512 17592 15524
rect 17644 15512 17650 15564
rect 17681 15555 17739 15561
rect 17681 15521 17693 15555
rect 17727 15552 17739 15555
rect 17862 15552 17868 15564
rect 17727 15524 17868 15552
rect 17727 15521 17739 15524
rect 17681 15515 17739 15521
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 17972 15561 18000 15592
rect 17957 15555 18015 15561
rect 17957 15521 17969 15555
rect 18003 15521 18015 15555
rect 18690 15552 18696 15564
rect 18651 15524 18696 15552
rect 17957 15515 18015 15521
rect 18690 15512 18696 15524
rect 18748 15512 18754 15564
rect 14369 15447 14427 15453
rect 16132 15456 16804 15484
rect 4798 15416 4804 15428
rect 4172 15388 4804 15416
rect 4798 15376 4804 15388
rect 4856 15416 4862 15428
rect 5350 15416 5356 15428
rect 4856 15388 5356 15416
rect 4856 15376 4862 15388
rect 5350 15376 5356 15388
rect 5408 15376 5414 15428
rect 11333 15419 11391 15425
rect 11333 15385 11345 15419
rect 11379 15416 11391 15419
rect 11379 15388 12112 15416
rect 11379 15385 11391 15388
rect 11333 15379 11391 15385
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15348 1639 15351
rect 1762 15348 1768 15360
rect 1627 15320 1768 15348
rect 1627 15317 1639 15320
rect 1581 15311 1639 15317
rect 1762 15308 1768 15320
rect 1820 15308 1826 15360
rect 3605 15351 3663 15357
rect 3605 15317 3617 15351
rect 3651 15348 3663 15351
rect 4430 15348 4436 15360
rect 3651 15320 4436 15348
rect 3651 15317 3663 15320
rect 3605 15311 3663 15317
rect 4430 15308 4436 15320
rect 4488 15308 4494 15360
rect 5261 15351 5319 15357
rect 5261 15317 5273 15351
rect 5307 15348 5319 15351
rect 5442 15348 5448 15360
rect 5307 15320 5448 15348
rect 5307 15317 5319 15320
rect 5261 15311 5319 15317
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 5537 15351 5595 15357
rect 5537 15317 5549 15351
rect 5583 15348 5595 15351
rect 5718 15348 5724 15360
rect 5583 15320 5724 15348
rect 5583 15317 5595 15320
rect 5537 15311 5595 15317
rect 5718 15308 5724 15320
rect 5776 15308 5782 15360
rect 11698 15308 11704 15360
rect 11756 15348 11762 15360
rect 11885 15351 11943 15357
rect 11885 15348 11897 15351
rect 11756 15320 11897 15348
rect 11756 15308 11762 15320
rect 11885 15317 11897 15320
rect 11931 15317 11943 15351
rect 12084 15348 12112 15388
rect 12434 15348 12440 15360
rect 12084 15320 12440 15348
rect 11885 15311 11943 15317
rect 12434 15308 12440 15320
rect 12492 15308 12498 15360
rect 12710 15308 12716 15360
rect 12768 15348 12774 15360
rect 15010 15348 15016 15360
rect 12768 15320 15016 15348
rect 12768 15308 12774 15320
rect 15010 15308 15016 15320
rect 15068 15308 15074 15360
rect 15746 15308 15752 15360
rect 15804 15348 15810 15360
rect 16132 15357 16160 15456
rect 16117 15351 16175 15357
rect 16117 15348 16129 15351
rect 15804 15320 16129 15348
rect 15804 15308 15810 15320
rect 16117 15317 16129 15320
rect 16163 15317 16175 15351
rect 17862 15348 17868 15360
rect 17823 15320 17868 15348
rect 16117 15311 16175 15317
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 17954 15308 17960 15360
rect 18012 15348 18018 15360
rect 18509 15351 18567 15357
rect 18509 15348 18521 15351
rect 18012 15320 18521 15348
rect 18012 15308 18018 15320
rect 18509 15317 18521 15320
rect 18555 15317 18567 15351
rect 18509 15311 18567 15317
rect 1104 15258 19044 15280
rect 1104 15206 3972 15258
rect 4024 15206 4036 15258
rect 4088 15206 4100 15258
rect 4152 15206 4164 15258
rect 4216 15206 9952 15258
rect 10004 15206 10016 15258
rect 10068 15206 10080 15258
rect 10132 15206 10144 15258
rect 10196 15206 15932 15258
rect 15984 15206 15996 15258
rect 16048 15206 16060 15258
rect 16112 15206 16124 15258
rect 16176 15206 19044 15258
rect 1104 15184 19044 15206
rect 4709 15147 4767 15153
rect 4709 15113 4721 15147
rect 4755 15144 4767 15147
rect 4982 15144 4988 15156
rect 4755 15116 4988 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 4982 15104 4988 15116
rect 5040 15104 5046 15156
rect 5350 15144 5356 15156
rect 5311 15116 5356 15144
rect 5350 15104 5356 15116
rect 5408 15104 5414 15156
rect 7650 15104 7656 15156
rect 7708 15144 7714 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7708 15116 7849 15144
rect 7708 15104 7714 15116
rect 7837 15113 7849 15116
rect 7883 15144 7895 15147
rect 9674 15144 9680 15156
rect 7883 15116 8340 15144
rect 9635 15116 9680 15144
rect 7883 15113 7895 15116
rect 7837 15107 7895 15113
rect 5626 15076 5632 15088
rect 5000 15048 5632 15076
rect 4706 14968 4712 15020
rect 4764 15008 4770 15020
rect 5000 15008 5028 15048
rect 5626 15036 5632 15048
rect 5684 15076 5690 15088
rect 5684 15048 7236 15076
rect 5684 15036 5690 15048
rect 4764 14980 5028 15008
rect 4764 14968 4770 14980
rect 4430 14900 4436 14952
rect 4488 14940 4494 14952
rect 5000 14949 5028 14980
rect 5169 15011 5227 15017
rect 5169 14977 5181 15011
rect 5215 15008 5227 15011
rect 7208 15008 7236 15048
rect 7282 15036 7288 15088
rect 7340 15076 7346 15088
rect 7558 15076 7564 15088
rect 7340 15048 7564 15076
rect 7340 15036 7346 15048
rect 7558 15036 7564 15048
rect 7616 15076 7622 15088
rect 7929 15079 7987 15085
rect 7929 15076 7941 15079
rect 7616 15048 7941 15076
rect 7616 15036 7622 15048
rect 7929 15045 7941 15048
rect 7975 15045 7987 15079
rect 7929 15039 7987 15045
rect 5215 14980 5396 15008
rect 7208 14980 7696 15008
rect 5215 14977 5227 14980
rect 5169 14971 5227 14977
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4488 14912 4905 14940
rect 4488 14900 4494 14912
rect 4893 14909 4905 14912
rect 4939 14909 4951 14943
rect 4893 14903 4951 14909
rect 4985 14943 5043 14949
rect 4985 14909 4997 14943
rect 5031 14909 5043 14943
rect 4985 14903 5043 14909
rect 4908 14872 4936 14903
rect 5074 14900 5080 14952
rect 5132 14940 5138 14952
rect 5261 14943 5319 14949
rect 5261 14940 5273 14943
rect 5132 14912 5273 14940
rect 5132 14900 5138 14912
rect 5261 14909 5273 14912
rect 5307 14909 5319 14943
rect 5261 14903 5319 14909
rect 5368 14872 5396 14980
rect 5442 14900 5448 14952
rect 5500 14940 5506 14952
rect 5537 14943 5595 14949
rect 5537 14940 5549 14943
rect 5500 14912 5549 14940
rect 5500 14900 5506 14912
rect 5537 14909 5549 14912
rect 5583 14909 5595 14943
rect 5718 14940 5724 14952
rect 5679 14912 5724 14940
rect 5537 14903 5595 14909
rect 5718 14900 5724 14912
rect 5776 14900 5782 14952
rect 5902 14900 5908 14952
rect 5960 14940 5966 14952
rect 7285 14943 7343 14949
rect 7285 14940 7297 14943
rect 5960 14912 7297 14940
rect 5960 14900 5966 14912
rect 7285 14909 7297 14912
rect 7331 14940 7343 14943
rect 7374 14940 7380 14952
rect 7331 14912 7380 14940
rect 7331 14909 7343 14912
rect 7285 14903 7343 14909
rect 7374 14900 7380 14912
rect 7432 14900 7438 14952
rect 7668 14949 7696 14980
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14940 7711 14943
rect 7926 14940 7932 14952
rect 7699 14912 7932 14940
rect 7699 14909 7711 14912
rect 7653 14903 7711 14909
rect 7926 14900 7932 14912
rect 7984 14900 7990 14952
rect 8202 14900 8208 14952
rect 8260 14940 8266 14952
rect 8312 14949 8340 15116
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 10410 15144 10416 15156
rect 10371 15116 10416 15144
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 9861 15011 9919 15017
rect 9861 14977 9873 15011
rect 9907 15008 9919 15011
rect 10321 15011 10379 15017
rect 9907 14980 10272 15008
rect 9907 14977 9919 14980
rect 9861 14971 9919 14977
rect 8297 14943 8355 14949
rect 8297 14940 8309 14943
rect 8260 14912 8309 14940
rect 8260 14900 8266 14912
rect 8297 14909 8309 14912
rect 8343 14909 8355 14943
rect 8297 14903 8355 14909
rect 9953 14943 10011 14949
rect 9953 14909 9965 14943
rect 9999 14909 10011 14943
rect 10244 14940 10272 14980
rect 10321 14977 10333 15011
rect 10367 15008 10379 15011
rect 10428 15008 10456 15104
rect 14461 15079 14519 15085
rect 14461 15045 14473 15079
rect 14507 15076 14519 15079
rect 14826 15076 14832 15088
rect 14507 15048 14832 15076
rect 14507 15045 14519 15048
rect 14461 15039 14519 15045
rect 12345 15011 12403 15017
rect 12345 15008 12357 15011
rect 10367 14980 10456 15008
rect 11900 14980 12357 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 11900 14952 11928 14980
rect 12345 14977 12357 14980
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 10781 14943 10839 14949
rect 10781 14940 10793 14943
rect 10244 14912 10793 14940
rect 9953 14903 10011 14909
rect 10781 14909 10793 14912
rect 10827 14940 10839 14943
rect 10962 14940 10968 14952
rect 10827 14912 10968 14940
rect 10827 14909 10839 14912
rect 10781 14903 10839 14909
rect 5920 14872 5948 14900
rect 7469 14875 7527 14881
rect 7469 14872 7481 14875
rect 4908 14844 5304 14872
rect 5368 14844 5948 14872
rect 7300 14844 7481 14872
rect 5276 14816 5304 14844
rect 7300 14816 7328 14844
rect 7469 14841 7481 14844
rect 7515 14841 7527 14875
rect 7469 14835 7527 14841
rect 7561 14875 7619 14881
rect 7561 14841 7573 14875
rect 7607 14841 7619 14875
rect 8110 14872 8116 14884
rect 8071 14844 8116 14872
rect 7561 14835 7619 14841
rect 5258 14764 5264 14816
rect 5316 14764 5322 14816
rect 7282 14764 7288 14816
rect 7340 14764 7346 14816
rect 7576 14804 7604 14835
rect 8110 14832 8116 14844
rect 8168 14832 8174 14884
rect 9968 14872 9996 14903
rect 10962 14900 10968 14912
rect 11020 14900 11026 14952
rect 11882 14940 11888 14952
rect 11843 14912 11888 14940
rect 11882 14900 11888 14912
rect 11940 14900 11946 14952
rect 12158 14940 12164 14952
rect 12119 14912 12164 14940
rect 12158 14900 12164 14912
rect 12216 14940 12222 14952
rect 12253 14943 12311 14949
rect 12253 14940 12265 14943
rect 12216 14912 12265 14940
rect 12216 14900 12222 14912
rect 12253 14909 12265 14912
rect 12299 14909 12311 14943
rect 12253 14903 12311 14909
rect 12449 14943 12507 14949
rect 12449 14909 12461 14943
rect 12495 14909 12507 14943
rect 12449 14903 12507 14909
rect 10318 14872 10324 14884
rect 9968 14844 10324 14872
rect 10318 14832 10324 14844
rect 10376 14872 10382 14884
rect 10597 14875 10655 14881
rect 10597 14872 10609 14875
rect 10376 14844 10609 14872
rect 10376 14832 10382 14844
rect 10597 14841 10609 14844
rect 10643 14841 10655 14875
rect 12066 14872 12072 14884
rect 11979 14844 12072 14872
rect 10597 14835 10655 14841
rect 12066 14832 12072 14844
rect 12124 14872 12130 14884
rect 12452 14872 12480 14903
rect 14476 14872 14504 15039
rect 14826 15036 14832 15048
rect 14884 15036 14890 15088
rect 17586 15008 17592 15020
rect 17052 14980 17592 15008
rect 14550 14900 14556 14952
rect 14608 14940 14614 14952
rect 14737 14943 14795 14949
rect 14737 14940 14749 14943
rect 14608 14912 14749 14940
rect 14608 14900 14614 14912
rect 14737 14909 14749 14912
rect 14783 14909 14795 14943
rect 14737 14903 14795 14909
rect 14826 14900 14832 14952
rect 14884 14940 14890 14952
rect 15013 14943 15071 14949
rect 15013 14940 15025 14943
rect 14884 14912 15025 14940
rect 14884 14900 14890 14912
rect 15013 14909 15025 14912
rect 15059 14909 15071 14943
rect 15013 14903 15071 14909
rect 16390 14900 16396 14952
rect 16448 14940 16454 14952
rect 17052 14949 17080 14980
rect 17586 14968 17592 14980
rect 17644 14968 17650 15020
rect 17037 14943 17095 14949
rect 17037 14940 17049 14943
rect 16448 14912 17049 14940
rect 16448 14900 16454 14912
rect 17037 14909 17049 14912
rect 17083 14909 17095 14943
rect 17037 14903 17095 14909
rect 17221 14943 17279 14949
rect 17221 14909 17233 14943
rect 17267 14940 17279 14943
rect 17862 14940 17868 14952
rect 17267 14912 17868 14940
rect 17267 14909 17279 14912
rect 17221 14903 17279 14909
rect 17862 14900 17868 14912
rect 17920 14900 17926 14952
rect 12124 14844 14504 14872
rect 17313 14875 17371 14881
rect 12124 14832 12130 14844
rect 17313 14841 17325 14875
rect 17359 14872 17371 14875
rect 17402 14872 17408 14884
rect 17359 14844 17408 14872
rect 17359 14841 17371 14844
rect 17313 14835 17371 14841
rect 17402 14832 17408 14844
rect 17460 14872 17466 14884
rect 17586 14872 17592 14884
rect 17460 14844 17592 14872
rect 17460 14832 17466 14844
rect 17586 14832 17592 14844
rect 17644 14832 17650 14884
rect 8294 14804 8300 14816
rect 7576 14776 8300 14804
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 11514 14764 11520 14816
rect 11572 14804 11578 14816
rect 11701 14807 11759 14813
rect 11701 14804 11713 14807
rect 11572 14776 11713 14804
rect 11572 14764 11578 14776
rect 11701 14773 11713 14776
rect 11747 14773 11759 14807
rect 14642 14804 14648 14816
rect 14603 14776 14648 14804
rect 11701 14767 11759 14773
rect 14642 14764 14648 14776
rect 14700 14764 14706 14816
rect 14734 14764 14740 14816
rect 14792 14804 14798 14816
rect 14829 14807 14887 14813
rect 14829 14804 14841 14807
rect 14792 14776 14841 14804
rect 14792 14764 14798 14776
rect 14829 14773 14841 14776
rect 14875 14804 14887 14807
rect 14918 14804 14924 14816
rect 14875 14776 14924 14804
rect 14875 14773 14887 14776
rect 14829 14767 14887 14773
rect 14918 14764 14924 14776
rect 14976 14764 14982 14816
rect 1104 14714 19044 14736
rect 1104 14662 6962 14714
rect 7014 14662 7026 14714
rect 7078 14662 7090 14714
rect 7142 14662 7154 14714
rect 7206 14662 12942 14714
rect 12994 14662 13006 14714
rect 13058 14662 13070 14714
rect 13122 14662 13134 14714
rect 13186 14662 19044 14714
rect 1104 14640 19044 14662
rect 5813 14603 5871 14609
rect 5813 14569 5825 14603
rect 5859 14600 5871 14603
rect 7466 14600 7472 14612
rect 5859 14572 7472 14600
rect 5859 14569 5871 14572
rect 5813 14563 5871 14569
rect 7466 14560 7472 14572
rect 7524 14600 7530 14612
rect 8110 14600 8116 14612
rect 7524 14572 8116 14600
rect 7524 14560 7530 14572
rect 5902 14532 5908 14544
rect 5184 14504 5908 14532
rect 1486 14464 1492 14476
rect 1447 14436 1492 14464
rect 1486 14424 1492 14436
rect 1544 14424 1550 14476
rect 2041 14467 2099 14473
rect 2041 14433 2053 14467
rect 2087 14464 2099 14467
rect 2590 14464 2596 14476
rect 2087 14436 2596 14464
rect 2087 14433 2099 14436
rect 2041 14427 2099 14433
rect 2590 14424 2596 14436
rect 2648 14424 2654 14476
rect 4982 14424 4988 14476
rect 5040 14464 5046 14476
rect 5184 14473 5212 14504
rect 5902 14492 5908 14504
rect 5960 14492 5966 14544
rect 7285 14535 7343 14541
rect 7285 14501 7297 14535
rect 7331 14532 7343 14535
rect 7331 14504 7420 14532
rect 7331 14501 7343 14504
rect 7285 14495 7343 14501
rect 5077 14467 5135 14473
rect 5077 14464 5089 14467
rect 5040 14436 5089 14464
rect 5040 14424 5046 14436
rect 5077 14433 5089 14436
rect 5123 14433 5135 14467
rect 5077 14427 5135 14433
rect 5169 14467 5227 14473
rect 5169 14433 5181 14467
rect 5215 14433 5227 14467
rect 5442 14464 5448 14476
rect 5403 14436 5448 14464
rect 5169 14427 5227 14433
rect 4798 14396 4804 14408
rect 4759 14368 4804 14396
rect 4798 14356 4804 14368
rect 4856 14356 4862 14408
rect 4985 14331 5043 14337
rect 4985 14297 4997 14331
rect 5031 14328 5043 14331
rect 5184 14328 5212 14427
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14464 5687 14467
rect 5718 14464 5724 14476
rect 5675 14436 5724 14464
rect 5675 14433 5687 14436
rect 5629 14427 5687 14433
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 7006 14464 7012 14476
rect 6967 14436 7012 14464
rect 7006 14424 7012 14436
rect 7064 14424 7070 14476
rect 7190 14424 7196 14476
rect 7248 14464 7254 14476
rect 7392 14473 7420 14504
rect 7377 14467 7435 14473
rect 7377 14464 7389 14467
rect 7248 14436 7389 14464
rect 7248 14424 7254 14436
rect 7377 14433 7389 14436
rect 7423 14433 7435 14467
rect 7377 14427 7435 14433
rect 7653 14467 7711 14473
rect 7653 14433 7665 14467
rect 7699 14433 7711 14467
rect 7653 14427 7711 14433
rect 5353 14399 5411 14405
rect 5353 14365 5365 14399
rect 5399 14396 5411 14399
rect 6178 14396 6184 14408
rect 5399 14368 6184 14396
rect 5399 14365 5411 14368
rect 5353 14359 5411 14365
rect 6178 14356 6184 14368
rect 6236 14356 6242 14408
rect 7285 14399 7343 14405
rect 7285 14365 7297 14399
rect 7331 14396 7343 14399
rect 7558 14396 7564 14408
rect 7331 14368 7564 14396
rect 7331 14365 7343 14368
rect 7285 14359 7343 14365
rect 7558 14356 7564 14368
rect 7616 14356 7622 14408
rect 5031 14300 5212 14328
rect 5031 14297 5043 14300
rect 4985 14291 5043 14297
rect 5442 14288 5448 14340
rect 5500 14328 5506 14340
rect 5537 14331 5595 14337
rect 5537 14328 5549 14331
rect 5500 14300 5549 14328
rect 5500 14288 5506 14300
rect 5537 14297 5549 14300
rect 5583 14297 5595 14331
rect 5537 14291 5595 14297
rect 7101 14331 7159 14337
rect 7101 14297 7113 14331
rect 7147 14328 7159 14331
rect 7374 14328 7380 14340
rect 7147 14300 7380 14328
rect 7147 14297 7159 14300
rect 7101 14291 7159 14297
rect 7374 14288 7380 14300
rect 7432 14328 7438 14340
rect 7668 14328 7696 14427
rect 7834 14396 7840 14408
rect 7795 14368 7840 14396
rect 7834 14356 7840 14368
rect 7892 14356 7898 14408
rect 7929 14399 7987 14405
rect 7929 14365 7941 14399
rect 7975 14396 7987 14399
rect 8036 14396 8064 14572
rect 8110 14560 8116 14572
rect 8168 14560 8174 14612
rect 10962 14600 10968 14612
rect 10923 14572 10968 14600
rect 10962 14560 10968 14572
rect 11020 14560 11026 14612
rect 11149 14603 11207 14609
rect 11149 14569 11161 14603
rect 11195 14600 11207 14603
rect 11514 14600 11520 14612
rect 11195 14572 11520 14600
rect 11195 14569 11207 14572
rect 11149 14563 11207 14569
rect 11514 14560 11520 14572
rect 11572 14560 11578 14612
rect 16758 14560 16764 14612
rect 16816 14600 16822 14612
rect 17037 14603 17095 14609
rect 17037 14600 17049 14603
rect 16816 14572 17049 14600
rect 16816 14560 16822 14572
rect 17037 14569 17049 14572
rect 17083 14569 17095 14603
rect 17037 14563 17095 14569
rect 16776 14504 17356 14532
rect 8113 14467 8171 14473
rect 8113 14433 8125 14467
rect 8159 14464 8171 14467
rect 8202 14464 8208 14476
rect 8159 14436 8208 14464
rect 8159 14433 8171 14436
rect 8113 14427 8171 14433
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 16776 14473 16804 14504
rect 17328 14473 17356 14504
rect 11146 14467 11204 14473
rect 11146 14433 11158 14467
rect 11192 14464 11204 14467
rect 16761 14467 16819 14473
rect 11192 14436 11652 14464
rect 11192 14433 11204 14436
rect 11146 14427 11204 14433
rect 11514 14396 11520 14408
rect 7975 14368 8064 14396
rect 11475 14368 11520 14396
rect 7975 14365 7987 14368
rect 7929 14359 7987 14365
rect 11514 14356 11520 14368
rect 11572 14356 11578 14408
rect 11624 14405 11652 14436
rect 16761 14433 16773 14467
rect 16807 14433 16819 14467
rect 16761 14427 16819 14433
rect 16945 14467 17003 14473
rect 16945 14433 16957 14467
rect 16991 14464 17003 14467
rect 17221 14467 17279 14473
rect 17221 14464 17233 14467
rect 16991 14436 17233 14464
rect 16991 14433 17003 14436
rect 16945 14427 17003 14433
rect 17221 14433 17233 14436
rect 17267 14433 17279 14467
rect 17221 14427 17279 14433
rect 17313 14467 17371 14473
rect 17313 14433 17325 14467
rect 17359 14464 17371 14467
rect 17586 14464 17592 14476
rect 17359 14436 17592 14464
rect 17359 14433 17371 14436
rect 17313 14427 17371 14433
rect 11609 14399 11667 14405
rect 11609 14365 11621 14399
rect 11655 14396 11667 14399
rect 12526 14396 12532 14408
rect 11655 14368 12532 14396
rect 11655 14365 11667 14368
rect 11609 14359 11667 14365
rect 12526 14356 12532 14368
rect 12584 14356 12590 14408
rect 17236 14396 17264 14427
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 17770 14396 17776 14408
rect 17236 14368 17776 14396
rect 17770 14356 17776 14368
rect 17828 14356 17834 14408
rect 8018 14328 8024 14340
rect 7432 14300 7696 14328
rect 7979 14300 8024 14328
rect 7432 14288 7438 14300
rect 7668 14272 7696 14300
rect 8018 14288 8024 14300
rect 8076 14288 8082 14340
rect 9398 14328 9404 14340
rect 8128 14300 9404 14328
rect 2041 14263 2099 14269
rect 2041 14229 2053 14263
rect 2087 14260 2099 14263
rect 2498 14260 2504 14272
rect 2087 14232 2504 14260
rect 2087 14229 2099 14232
rect 2041 14223 2099 14229
rect 2498 14220 2504 14232
rect 2556 14220 2562 14272
rect 4890 14260 4896 14272
rect 4851 14232 4896 14260
rect 4890 14220 4896 14232
rect 4948 14260 4954 14272
rect 5718 14260 5724 14272
rect 4948 14232 5724 14260
rect 4948 14220 4954 14232
rect 5718 14220 5724 14232
rect 5776 14220 5782 14272
rect 7466 14260 7472 14272
rect 7427 14232 7472 14260
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 7650 14260 7656 14272
rect 7563 14232 7656 14260
rect 7650 14220 7656 14232
rect 7708 14260 7714 14272
rect 8128 14260 8156 14300
rect 9398 14288 9404 14300
rect 9456 14288 9462 14340
rect 7708 14232 8156 14260
rect 8297 14263 8355 14269
rect 7708 14220 7714 14232
rect 8297 14229 8309 14263
rect 8343 14260 8355 14263
rect 9214 14260 9220 14272
rect 8343 14232 9220 14260
rect 8343 14229 8355 14232
rect 8297 14223 8355 14229
rect 9214 14220 9220 14232
rect 9272 14220 9278 14272
rect 1104 14170 19044 14192
rect 1104 14118 3972 14170
rect 4024 14118 4036 14170
rect 4088 14118 4100 14170
rect 4152 14118 4164 14170
rect 4216 14118 9952 14170
rect 10004 14118 10016 14170
rect 10068 14118 10080 14170
rect 10132 14118 10144 14170
rect 10196 14118 15932 14170
rect 15984 14118 15996 14170
rect 16048 14118 16060 14170
rect 16112 14118 16124 14170
rect 16176 14118 19044 14170
rect 1104 14096 19044 14118
rect 7006 14016 7012 14068
rect 7064 14056 7070 14068
rect 7282 14056 7288 14068
rect 7064 14028 7288 14056
rect 7064 14016 7070 14028
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 12621 14059 12679 14065
rect 12621 14056 12633 14059
rect 11112 14028 12633 14056
rect 11112 14016 11118 14028
rect 12621 14025 12633 14028
rect 12667 14025 12679 14059
rect 12621 14019 12679 14025
rect 14642 14016 14648 14068
rect 14700 14056 14706 14068
rect 14921 14059 14979 14065
rect 14921 14056 14933 14059
rect 14700 14028 14933 14056
rect 14700 14016 14706 14028
rect 14921 14025 14933 14028
rect 14967 14025 14979 14059
rect 14921 14019 14979 14025
rect 15473 14059 15531 14065
rect 15473 14025 15485 14059
rect 15519 14056 15531 14059
rect 15654 14056 15660 14068
rect 15519 14028 15660 14056
rect 15519 14025 15531 14028
rect 15473 14019 15531 14025
rect 15654 14016 15660 14028
rect 15712 14056 15718 14068
rect 16390 14056 16396 14068
rect 15712 14028 16396 14056
rect 15712 14016 15718 14028
rect 16390 14016 16396 14028
rect 16448 14016 16454 14068
rect 18506 14056 18512 14068
rect 18467 14028 18512 14056
rect 18506 14016 18512 14028
rect 18564 14016 18570 14068
rect 10045 13991 10103 13997
rect 10045 13988 10057 13991
rect 5361 13960 7696 13988
rect 4522 13880 4528 13932
rect 4580 13920 4586 13932
rect 5361 13920 5389 13960
rect 4580 13892 5389 13920
rect 4580 13880 4586 13892
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 1486 13812 1492 13864
rect 1544 13852 1550 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1544 13824 2053 13852
rect 1544 13812 1550 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2498 13852 2504 13864
rect 2459 13824 2504 13852
rect 2041 13815 2099 13821
rect 2498 13812 2504 13824
rect 2556 13812 2562 13864
rect 4890 13861 4896 13864
rect 2593 13855 2651 13861
rect 2593 13821 2605 13855
rect 2639 13852 2651 13855
rect 2869 13855 2927 13861
rect 2869 13852 2881 13855
rect 2639 13824 2881 13852
rect 2639 13821 2651 13824
rect 2593 13815 2651 13821
rect 2869 13821 2881 13824
rect 2915 13821 2927 13855
rect 4888 13852 4896 13861
rect 4851 13824 4896 13852
rect 2869 13815 2927 13821
rect 4888 13815 4896 13824
rect 4890 13812 4896 13815
rect 4948 13812 4954 13864
rect 5361 13861 5389 13892
rect 7668 13920 7696 13960
rect 9048 13960 10057 13988
rect 7668 13892 8984 13920
rect 5442 13861 5448 13864
rect 5260 13855 5318 13861
rect 5260 13821 5272 13855
rect 5306 13821 5318 13855
rect 5260 13815 5318 13821
rect 5346 13855 5404 13861
rect 5346 13821 5358 13855
rect 5392 13821 5404 13855
rect 5346 13815 5404 13821
rect 5437 13815 5448 13861
rect 5500 13852 5506 13864
rect 5718 13852 5724 13864
rect 5500 13824 5537 13852
rect 5679 13824 5724 13852
rect 4985 13787 5043 13793
rect 4985 13753 4997 13787
rect 5031 13753 5043 13787
rect 4985 13747 5043 13753
rect 1578 13716 1584 13728
rect 1539 13688 1584 13716
rect 1578 13676 1584 13688
rect 1636 13676 1642 13728
rect 3050 13716 3056 13728
rect 3011 13688 3056 13716
rect 3050 13676 3056 13688
rect 3108 13676 3114 13728
rect 4709 13719 4767 13725
rect 4709 13685 4721 13719
rect 4755 13716 4767 13719
rect 4798 13716 4804 13728
rect 4755 13688 4804 13716
rect 4755 13685 4767 13688
rect 4709 13679 4767 13685
rect 4798 13676 4804 13688
rect 4856 13676 4862 13728
rect 5000 13716 5028 13747
rect 5074 13744 5080 13796
rect 5132 13784 5138 13796
rect 5275 13784 5303 13815
rect 5442 13812 5448 13815
rect 5500 13812 5506 13824
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 7190 13861 7196 13864
rect 7188 13852 7196 13861
rect 7151 13824 7196 13852
rect 7188 13815 7196 13824
rect 7190 13812 7196 13815
rect 7248 13812 7254 13864
rect 7466 13812 7472 13864
rect 7524 13861 7530 13864
rect 7668 13861 7696 13892
rect 7524 13855 7563 13861
rect 7551 13821 7563 13855
rect 7524 13815 7563 13821
rect 7653 13855 7711 13861
rect 7653 13821 7665 13855
rect 7699 13821 7711 13855
rect 7653 13815 7711 13821
rect 7929 13855 7987 13861
rect 7929 13821 7941 13855
rect 7975 13852 7987 13855
rect 8018 13852 8024 13864
rect 7975 13824 8024 13852
rect 7975 13821 7987 13824
rect 7929 13815 7987 13821
rect 7524 13812 7530 13815
rect 5813 13787 5871 13793
rect 5813 13784 5825 13787
rect 5132 13756 5177 13784
rect 5275 13756 5825 13784
rect 5132 13744 5138 13756
rect 5813 13753 5825 13756
rect 5859 13753 5871 13787
rect 5813 13747 5871 13753
rect 7285 13787 7343 13793
rect 7285 13753 7297 13787
rect 7331 13753 7343 13787
rect 7285 13747 7343 13753
rect 5537 13719 5595 13725
rect 5537 13716 5549 13719
rect 5000 13688 5549 13716
rect 5537 13685 5549 13688
rect 5583 13685 5595 13719
rect 5537 13679 5595 13685
rect 6822 13676 6828 13728
rect 6880 13716 6886 13728
rect 7009 13719 7067 13725
rect 7009 13716 7021 13719
rect 6880 13688 7021 13716
rect 6880 13676 6886 13688
rect 7009 13685 7021 13688
rect 7055 13685 7067 13719
rect 7300 13716 7328 13747
rect 7374 13744 7380 13796
rect 7432 13784 7438 13796
rect 7944 13784 7972 13815
rect 8018 13812 8024 13824
rect 8076 13812 8082 13864
rect 8956 13861 8984 13892
rect 9048 13861 9076 13960
rect 10045 13957 10057 13960
rect 10091 13957 10103 13991
rect 17221 13991 17279 13997
rect 17221 13988 17233 13991
rect 10045 13951 10103 13957
rect 12820 13960 17233 13988
rect 12820 13929 12848 13960
rect 12805 13923 12863 13929
rect 9232 13892 9720 13920
rect 9232 13864 9260 13892
rect 8941 13855 8999 13861
rect 8941 13821 8953 13855
rect 8987 13821 8999 13855
rect 8941 13815 8999 13821
rect 9034 13855 9092 13861
rect 9034 13821 9046 13855
rect 9080 13821 9092 13855
rect 9214 13852 9220 13864
rect 9175 13824 9220 13852
rect 9034 13815 9092 13821
rect 9214 13812 9220 13824
rect 9272 13812 9278 13864
rect 9490 13861 9496 13864
rect 9447 13855 9496 13861
rect 9447 13821 9459 13855
rect 9493 13821 9496 13855
rect 9447 13815 9496 13821
rect 9490 13812 9496 13815
rect 9548 13812 9554 13864
rect 9692 13861 9720 13892
rect 12805 13889 12817 13923
rect 12851 13889 12863 13923
rect 13173 13923 13231 13929
rect 13173 13920 13185 13923
rect 12805 13883 12863 13889
rect 12912 13892 13185 13920
rect 9669 13855 9727 13861
rect 9669 13821 9681 13855
rect 9715 13821 9727 13855
rect 9669 13815 9727 13821
rect 9858 13812 9864 13864
rect 9916 13852 9922 13864
rect 12912 13861 12940 13892
rect 13173 13889 13185 13892
rect 13219 13920 13231 13923
rect 13262 13920 13268 13932
rect 13219 13892 13268 13920
rect 13219 13889 13231 13892
rect 13173 13883 13231 13889
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 13556 13861 13584 13960
rect 17221 13957 17233 13960
rect 17267 13957 17279 13991
rect 17221 13951 17279 13957
rect 15838 13880 15844 13932
rect 15896 13920 15902 13932
rect 15896 13892 16252 13920
rect 15896 13880 15902 13892
rect 9953 13855 10011 13861
rect 9953 13852 9965 13855
rect 9916 13824 9965 13852
rect 9916 13812 9922 13824
rect 9953 13821 9965 13824
rect 9999 13821 10011 13855
rect 9953 13815 10011 13821
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13821 12955 13855
rect 13541 13855 13599 13861
rect 13541 13852 13553 13855
rect 12897 13815 12955 13821
rect 13280 13824 13553 13852
rect 13280 13793 13308 13824
rect 13541 13821 13553 13824
rect 13587 13821 13599 13855
rect 13541 13815 13599 13821
rect 15013 13855 15071 13861
rect 15013 13821 15025 13855
rect 15059 13852 15071 13855
rect 15286 13852 15292 13864
rect 15059 13824 15148 13852
rect 15247 13824 15292 13852
rect 15059 13821 15071 13824
rect 15013 13815 15071 13821
rect 7432 13756 7972 13784
rect 9309 13787 9367 13793
rect 7432 13744 7438 13756
rect 9309 13753 9321 13787
rect 9355 13784 9367 13787
rect 9769 13787 9827 13793
rect 9769 13784 9781 13787
rect 9355 13756 9781 13784
rect 9355 13753 9367 13756
rect 9309 13747 9367 13753
rect 9769 13753 9781 13756
rect 9815 13753 9827 13787
rect 9769 13747 9827 13753
rect 13265 13787 13323 13793
rect 13265 13753 13277 13787
rect 13311 13753 13323 13787
rect 13265 13747 13323 13753
rect 7837 13719 7895 13725
rect 7837 13716 7849 13719
rect 7300 13688 7849 13716
rect 7009 13679 7067 13685
rect 7837 13685 7849 13688
rect 7883 13685 7895 13719
rect 9582 13716 9588 13728
rect 9543 13688 9588 13716
rect 7837 13679 7895 13685
rect 9582 13676 9588 13688
rect 9640 13676 9646 13728
rect 13446 13716 13452 13728
rect 13407 13688 13452 13716
rect 13446 13676 13452 13688
rect 13504 13676 13510 13728
rect 15010 13676 15016 13728
rect 15068 13716 15074 13728
rect 15120 13725 15148 13824
rect 15286 13812 15292 13824
rect 15344 13812 15350 13864
rect 15470 13852 15476 13864
rect 15431 13824 15476 13852
rect 15470 13812 15476 13824
rect 15528 13812 15534 13864
rect 15746 13812 15752 13864
rect 15804 13852 15810 13864
rect 16117 13855 16175 13861
rect 16117 13852 16129 13855
rect 15804 13824 16129 13852
rect 15804 13812 15810 13824
rect 16117 13821 16129 13824
rect 16163 13821 16175 13855
rect 16224 13852 16252 13892
rect 16293 13855 16351 13861
rect 16293 13852 16305 13855
rect 16224 13824 16305 13852
rect 16117 13815 16175 13821
rect 16293 13821 16305 13824
rect 16339 13821 16351 13855
rect 17402 13852 17408 13864
rect 17363 13824 17408 13852
rect 16293 13815 16351 13821
rect 15304 13784 15332 13812
rect 16025 13787 16083 13793
rect 16025 13784 16037 13787
rect 15304 13756 16037 13784
rect 16025 13753 16037 13756
rect 16071 13753 16083 13787
rect 16132 13784 16160 13815
rect 17402 13812 17408 13824
rect 17460 13812 17466 13864
rect 17586 13852 17592 13864
rect 17547 13824 17592 13852
rect 17586 13812 17592 13824
rect 17644 13812 17650 13864
rect 17770 13852 17776 13864
rect 17731 13824 17776 13852
rect 17770 13812 17776 13824
rect 17828 13812 17834 13864
rect 18690 13852 18696 13864
rect 18651 13824 18696 13852
rect 18690 13812 18696 13824
rect 18748 13812 18754 13864
rect 17494 13784 17500 13796
rect 16132 13756 17500 13784
rect 16025 13747 16083 13753
rect 17494 13744 17500 13756
rect 17552 13744 17558 13796
rect 15105 13719 15163 13725
rect 15105 13716 15117 13719
rect 15068 13688 15117 13716
rect 15068 13676 15074 13688
rect 15105 13685 15117 13688
rect 15151 13685 15163 13719
rect 15105 13679 15163 13685
rect 1104 13626 19044 13648
rect 1104 13574 6962 13626
rect 7014 13574 7026 13626
rect 7078 13574 7090 13626
rect 7142 13574 7154 13626
rect 7206 13574 12942 13626
rect 12994 13574 13006 13626
rect 13058 13574 13070 13626
rect 13122 13574 13134 13626
rect 13186 13574 19044 13626
rect 1104 13552 19044 13574
rect 1486 13512 1492 13524
rect 1447 13484 1492 13512
rect 1486 13472 1492 13484
rect 1544 13472 1550 13524
rect 1946 13512 1952 13524
rect 1907 13484 1952 13512
rect 1946 13472 1952 13484
rect 2004 13472 2010 13524
rect 3050 13512 3056 13524
rect 2700 13484 3056 13512
rect 2700 13453 2728 13484
rect 3050 13472 3056 13484
rect 3108 13512 3114 13524
rect 3605 13515 3663 13521
rect 3605 13512 3617 13515
rect 3108 13484 3617 13512
rect 3108 13472 3114 13484
rect 3605 13481 3617 13484
rect 3651 13481 3663 13515
rect 3605 13475 3663 13481
rect 5074 13472 5080 13524
rect 5132 13512 5138 13524
rect 5442 13512 5448 13524
rect 5132 13484 5448 13512
rect 5132 13472 5138 13484
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 9674 13512 9680 13524
rect 9635 13484 9680 13512
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 12526 13512 12532 13524
rect 12487 13484 12532 13512
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 12713 13515 12771 13521
rect 12713 13481 12725 13515
rect 12759 13512 12771 13515
rect 12802 13512 12808 13524
rect 12759 13484 12808 13512
rect 12759 13481 12771 13484
rect 12713 13475 12771 13481
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 13449 13515 13507 13521
rect 13449 13512 13461 13515
rect 13096 13484 13461 13512
rect 2685 13447 2743 13453
rect 2685 13413 2697 13447
rect 2731 13413 2743 13447
rect 9769 13447 9827 13453
rect 2685 13407 2743 13413
rect 3068 13416 4108 13444
rect 1857 13379 1915 13385
rect 1857 13345 1869 13379
rect 1903 13345 1915 13379
rect 2590 13376 2596 13388
rect 2551 13348 2596 13376
rect 1857 13339 1915 13345
rect 1872 13172 1900 13339
rect 2590 13336 2596 13348
rect 2648 13376 2654 13388
rect 2866 13376 2872 13388
rect 2648 13348 2872 13376
rect 2648 13336 2654 13348
rect 2866 13336 2872 13348
rect 2924 13376 2930 13388
rect 3068 13376 3096 13416
rect 4080 13385 4108 13416
rect 9769 13413 9781 13447
rect 9815 13444 9827 13447
rect 10413 13447 10471 13453
rect 10413 13444 10425 13447
rect 9815 13416 10425 13444
rect 9815 13413 9827 13416
rect 9769 13407 9827 13413
rect 10413 13413 10425 13416
rect 10459 13413 10471 13447
rect 10413 13407 10471 13413
rect 11422 13404 11428 13456
rect 11480 13404 11486 13456
rect 2924 13348 3096 13376
rect 3145 13379 3203 13385
rect 2924 13336 2930 13348
rect 3145 13345 3157 13379
rect 3191 13345 3203 13379
rect 3145 13339 3203 13345
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13345 4123 13379
rect 9122 13376 9128 13388
rect 9083 13348 9128 13376
rect 4065 13339 4123 13345
rect 2038 13308 2044 13320
rect 1999 13280 2044 13308
rect 2038 13268 2044 13280
rect 2096 13268 2102 13320
rect 3160 13308 3188 13339
rect 9122 13336 9128 13348
rect 9180 13336 9186 13388
rect 9398 13376 9404 13388
rect 9359 13348 9404 13376
rect 9398 13336 9404 13348
rect 9456 13336 9462 13388
rect 9490 13336 9496 13388
rect 9548 13376 9554 13388
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 9548 13348 10057 13376
rect 9548 13336 9554 13348
rect 10045 13345 10057 13348
rect 10091 13345 10103 13379
rect 10045 13339 10103 13345
rect 12710 13379 12768 13385
rect 12710 13345 12722 13379
rect 12756 13376 12768 13379
rect 13096 13376 13124 13484
rect 13449 13481 13461 13484
rect 13495 13512 13507 13515
rect 15286 13512 15292 13524
rect 13495 13484 13860 13512
rect 13495 13481 13507 13484
rect 13449 13475 13507 13481
rect 13265 13447 13323 13453
rect 13265 13444 13277 13447
rect 13188 13416 13277 13444
rect 13188 13385 13216 13416
rect 13265 13413 13277 13416
rect 13311 13444 13323 13447
rect 13725 13447 13783 13453
rect 13725 13444 13737 13447
rect 13311 13416 13737 13444
rect 13311 13413 13323 13416
rect 13265 13407 13323 13413
rect 13725 13413 13737 13416
rect 13771 13413 13783 13447
rect 13725 13407 13783 13413
rect 13832 13388 13860 13484
rect 14384 13484 15292 13512
rect 12756 13348 13124 13376
rect 13173 13379 13231 13385
rect 12756 13345 12768 13348
rect 12710 13339 12768 13345
rect 13173 13345 13185 13379
rect 13219 13345 13231 13379
rect 13173 13339 13231 13345
rect 13541 13379 13599 13385
rect 13541 13345 13553 13379
rect 13587 13376 13599 13379
rect 13633 13379 13691 13385
rect 13633 13376 13645 13379
rect 13587 13348 13645 13376
rect 13587 13345 13599 13348
rect 13541 13339 13599 13345
rect 13633 13345 13645 13348
rect 13679 13345 13691 13379
rect 13814 13376 13820 13388
rect 13775 13348 13820 13376
rect 13633 13339 13691 13345
rect 3234 13308 3240 13320
rect 3160 13280 3240 13308
rect 3234 13268 3240 13280
rect 3292 13268 3298 13320
rect 7926 13268 7932 13320
rect 7984 13308 7990 13320
rect 9217 13311 9275 13317
rect 9217 13308 9229 13311
rect 7984 13280 9229 13308
rect 7984 13268 7990 13280
rect 9217 13277 9229 13280
rect 9263 13277 9275 13311
rect 9217 13271 9275 13277
rect 9582 13268 9588 13320
rect 9640 13308 9646 13320
rect 9769 13311 9827 13317
rect 9769 13308 9781 13311
rect 9640 13280 9781 13308
rect 9640 13268 9646 13280
rect 9769 13277 9781 13280
rect 9815 13277 9827 13311
rect 9769 13271 9827 13277
rect 10137 13311 10195 13317
rect 10137 13277 10149 13311
rect 10183 13308 10195 13311
rect 10410 13308 10416 13320
rect 10183 13280 10416 13308
rect 10183 13277 10195 13280
rect 10137 13271 10195 13277
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 12802 13268 12808 13320
rect 12860 13308 12866 13320
rect 13556 13308 13584 13339
rect 13814 13336 13820 13348
rect 13872 13336 13878 13388
rect 14384 13385 14412 13484
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 15378 13472 15384 13524
rect 15436 13512 15442 13524
rect 15436 13484 16620 13512
rect 15436 13472 15442 13484
rect 14645 13447 14703 13453
rect 14645 13413 14657 13447
rect 14691 13444 14703 13447
rect 15304 13444 15332 13472
rect 16592 13453 16620 13484
rect 17402 13472 17408 13524
rect 17460 13512 17466 13524
rect 17681 13515 17739 13521
rect 17681 13512 17693 13515
rect 17460 13484 17693 13512
rect 17460 13472 17466 13484
rect 17681 13481 17693 13484
rect 17727 13512 17739 13515
rect 18046 13512 18052 13524
rect 17727 13484 18052 13512
rect 17727 13481 17739 13484
rect 17681 13475 17739 13481
rect 18046 13472 18052 13484
rect 18104 13472 18110 13524
rect 16577 13447 16635 13453
rect 14691 13416 15148 13444
rect 15304 13416 16160 13444
rect 14691 13413 14703 13416
rect 14645 13407 14703 13413
rect 14369 13379 14427 13385
rect 14369 13345 14381 13379
rect 14415 13345 14427 13379
rect 14826 13376 14832 13388
rect 14787 13348 14832 13376
rect 14369 13339 14427 13345
rect 14826 13336 14832 13348
rect 14884 13336 14890 13388
rect 15010 13376 15016 13388
rect 14971 13348 15016 13376
rect 15010 13336 15016 13348
rect 15068 13336 15074 13388
rect 15120 13385 15148 13416
rect 15117 13379 15175 13385
rect 15117 13345 15129 13379
rect 15163 13345 15175 13379
rect 15565 13379 15623 13385
rect 15565 13376 15577 13379
rect 15117 13339 15175 13345
rect 15212 13348 15577 13376
rect 12860 13280 13584 13308
rect 14645 13311 14703 13317
rect 12860 13268 12866 13280
rect 14645 13277 14657 13311
rect 14691 13277 14703 13311
rect 14645 13271 14703 13277
rect 3605 13243 3663 13249
rect 3605 13209 3617 13243
rect 3651 13240 3663 13243
rect 3881 13243 3939 13249
rect 3881 13240 3893 13243
rect 3651 13212 3893 13240
rect 3651 13209 3663 13212
rect 3605 13203 3663 13209
rect 3881 13209 3893 13212
rect 3927 13209 3939 13243
rect 3881 13203 3939 13209
rect 4890 13200 4896 13252
rect 4948 13240 4954 13252
rect 5166 13240 5172 13252
rect 4948 13212 5172 13240
rect 4948 13200 4954 13212
rect 5166 13200 5172 13212
rect 5224 13240 5230 13252
rect 7190 13240 7196 13252
rect 5224 13212 7196 13240
rect 5224 13200 5230 13212
rect 7190 13200 7196 13212
rect 7248 13240 7254 13252
rect 9953 13243 10011 13249
rect 9953 13240 9965 13243
rect 7248 13212 9965 13240
rect 7248 13200 7254 13212
rect 9953 13209 9965 13212
rect 9999 13209 10011 13243
rect 9953 13203 10011 13209
rect 13081 13243 13139 13249
rect 13081 13209 13093 13243
rect 13127 13240 13139 13243
rect 13446 13240 13452 13252
rect 13127 13212 13452 13240
rect 13127 13209 13139 13212
rect 13081 13203 13139 13209
rect 13446 13200 13452 13212
rect 13504 13200 13510 13252
rect 14660 13240 14688 13271
rect 14734 13268 14740 13320
rect 14792 13308 14798 13320
rect 14921 13311 14979 13317
rect 14921 13308 14933 13311
rect 14792 13280 14933 13308
rect 14792 13268 14798 13280
rect 14921 13277 14933 13280
rect 14967 13308 14979 13311
rect 15212 13308 15240 13348
rect 15565 13345 15577 13348
rect 15611 13345 15623 13379
rect 15746 13376 15752 13388
rect 15707 13348 15752 13376
rect 15565 13339 15623 13345
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 15838 13336 15844 13388
rect 15896 13376 15902 13388
rect 16132 13385 16160 13416
rect 16577 13413 16589 13447
rect 16623 13413 16635 13447
rect 16577 13407 16635 13413
rect 16117 13379 16175 13385
rect 15896 13348 15941 13376
rect 15896 13336 15902 13348
rect 16117 13345 16129 13379
rect 16163 13345 16175 13379
rect 16117 13339 16175 13345
rect 16301 13379 16359 13385
rect 16301 13345 16313 13379
rect 16347 13376 16359 13379
rect 16393 13379 16451 13385
rect 16393 13376 16405 13379
rect 16347 13348 16405 13376
rect 16347 13345 16359 13348
rect 16301 13339 16359 13345
rect 16393 13345 16405 13348
rect 16439 13345 16451 13379
rect 16393 13339 16451 13345
rect 17126 13336 17132 13388
rect 17184 13376 17190 13388
rect 17494 13376 17500 13388
rect 17184 13348 17500 13376
rect 17184 13336 17190 13348
rect 17494 13336 17500 13348
rect 17552 13376 17558 13388
rect 17622 13379 17680 13385
rect 17622 13376 17634 13379
rect 17552 13348 17634 13376
rect 17552 13336 17558 13348
rect 17622 13345 17634 13348
rect 17668 13376 17680 13379
rect 18141 13379 18199 13385
rect 18141 13376 18153 13379
rect 17668 13348 18153 13376
rect 17668 13345 17680 13348
rect 17622 13339 17680 13345
rect 18141 13345 18153 13348
rect 18187 13345 18199 13379
rect 18141 13339 18199 13345
rect 14967 13280 15240 13308
rect 15289 13311 15347 13317
rect 14967 13277 14979 13280
rect 14921 13271 14979 13277
rect 15289 13277 15301 13311
rect 15335 13308 15347 13311
rect 15378 13308 15384 13320
rect 15335 13280 15384 13308
rect 15335 13277 15347 13280
rect 15289 13271 15347 13277
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 15654 13268 15660 13320
rect 15712 13308 15718 13320
rect 15933 13311 15991 13317
rect 15933 13308 15945 13311
rect 15712 13280 15945 13308
rect 15712 13268 15718 13280
rect 15933 13277 15945 13280
rect 15979 13277 15991 13311
rect 15933 13271 15991 13277
rect 15470 13240 15476 13252
rect 14660 13212 15476 13240
rect 15470 13200 15476 13212
rect 15528 13200 15534 13252
rect 4522 13172 4528 13184
rect 1872 13144 4528 13172
rect 4522 13132 4528 13144
rect 4580 13132 4586 13184
rect 11882 13172 11888 13184
rect 11843 13144 11888 13172
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 13262 13172 13268 13184
rect 13223 13144 13268 13172
rect 13262 13132 13268 13144
rect 13320 13132 13326 13184
rect 14461 13175 14519 13181
rect 14461 13141 14473 13175
rect 14507 13172 14519 13175
rect 15672 13172 15700 13268
rect 17497 13243 17555 13249
rect 17497 13209 17509 13243
rect 17543 13240 17555 13243
rect 17770 13240 17776 13252
rect 17543 13212 17776 13240
rect 17543 13209 17555 13212
rect 17497 13203 17555 13209
rect 17770 13200 17776 13212
rect 17828 13200 17834 13252
rect 14507 13144 15700 13172
rect 14507 13141 14519 13144
rect 14461 13135 14519 13141
rect 16390 13132 16396 13184
rect 16448 13172 16454 13184
rect 16761 13175 16819 13181
rect 16761 13172 16773 13175
rect 16448 13144 16773 13172
rect 16448 13132 16454 13144
rect 16761 13141 16773 13144
rect 16807 13141 16819 13175
rect 18046 13172 18052 13184
rect 18007 13144 18052 13172
rect 16761 13135 16819 13141
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 1104 13082 19044 13104
rect 1104 13030 3972 13082
rect 4024 13030 4036 13082
rect 4088 13030 4100 13082
rect 4152 13030 4164 13082
rect 4216 13030 9952 13082
rect 10004 13030 10016 13082
rect 10068 13030 10080 13082
rect 10132 13030 10144 13082
rect 10196 13030 15932 13082
rect 15984 13030 15996 13082
rect 16048 13030 16060 13082
rect 16112 13030 16124 13082
rect 16176 13030 19044 13082
rect 1104 13008 19044 13030
rect 3234 12928 3240 12980
rect 3292 12968 3298 12980
rect 8941 12971 8999 12977
rect 8941 12968 8953 12971
rect 3292 12940 8953 12968
rect 3292 12928 3298 12940
rect 8941 12937 8953 12940
rect 8987 12937 8999 12971
rect 8941 12931 8999 12937
rect 11333 12971 11391 12977
rect 11333 12937 11345 12971
rect 11379 12968 11391 12971
rect 11422 12968 11428 12980
rect 11379 12940 11428 12968
rect 11379 12937 11391 12940
rect 11333 12931 11391 12937
rect 11422 12928 11428 12940
rect 11480 12928 11486 12980
rect 15197 12971 15255 12977
rect 15197 12937 15209 12971
rect 15243 12968 15255 12971
rect 15470 12968 15476 12980
rect 15243 12940 15476 12968
rect 15243 12937 15255 12940
rect 15197 12931 15255 12937
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 4890 12860 4896 12912
rect 4948 12900 4954 12912
rect 4985 12903 5043 12909
rect 4985 12900 4997 12903
rect 4948 12872 4997 12900
rect 4948 12860 4954 12872
rect 4985 12869 4997 12872
rect 5031 12869 5043 12903
rect 4985 12863 5043 12869
rect 5074 12860 5080 12912
rect 5132 12900 5138 12912
rect 5169 12903 5227 12909
rect 5169 12900 5181 12903
rect 5132 12872 5181 12900
rect 5132 12860 5138 12872
rect 5169 12869 5181 12872
rect 5215 12869 5227 12903
rect 5626 12900 5632 12912
rect 5587 12872 5632 12900
rect 5169 12863 5227 12869
rect 5626 12860 5632 12872
rect 5684 12860 5690 12912
rect 7190 12860 7196 12912
rect 7248 12900 7254 12912
rect 7248 12872 7293 12900
rect 7248 12860 7254 12872
rect 7374 12860 7380 12912
rect 7432 12900 7438 12912
rect 7469 12903 7527 12909
rect 7469 12900 7481 12903
rect 7432 12872 7481 12900
rect 7432 12860 7438 12872
rect 7469 12869 7481 12872
rect 7515 12869 7527 12903
rect 7469 12863 7527 12869
rect 7650 12860 7656 12912
rect 7708 12900 7714 12912
rect 7926 12900 7932 12912
rect 7708 12872 7788 12900
rect 7887 12872 7932 12900
rect 7708 12860 7714 12872
rect 4798 12832 4804 12844
rect 4759 12804 4804 12832
rect 4798 12792 4804 12804
rect 4856 12792 4862 12844
rect 5902 12832 5908 12844
rect 5460 12804 5908 12832
rect 5077 12767 5135 12773
rect 5077 12733 5089 12767
rect 5123 12733 5135 12767
rect 5350 12764 5356 12776
rect 5311 12736 5356 12764
rect 5077 12727 5135 12733
rect 5092 12696 5120 12727
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 5460 12773 5488 12804
rect 5902 12792 5908 12804
rect 5960 12792 5966 12844
rect 6914 12792 6920 12844
rect 6972 12832 6978 12844
rect 7009 12835 7067 12841
rect 7009 12832 7021 12835
rect 6972 12804 7021 12832
rect 6972 12792 6978 12804
rect 7009 12801 7021 12804
rect 7055 12801 7067 12835
rect 7009 12795 7067 12801
rect 5445 12767 5503 12773
rect 5445 12733 5457 12767
rect 5491 12733 5503 12767
rect 5445 12727 5503 12733
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12764 5779 12767
rect 6270 12764 6276 12776
rect 5767 12736 6276 12764
rect 5767 12733 5779 12736
rect 5721 12727 5779 12733
rect 5736 12696 5764 12727
rect 6270 12724 6276 12736
rect 6328 12724 6334 12776
rect 7285 12767 7343 12773
rect 7285 12733 7297 12767
rect 7331 12733 7343 12767
rect 7285 12727 7343 12733
rect 5092 12668 5764 12696
rect 7300 12696 7328 12727
rect 7558 12724 7564 12776
rect 7616 12764 7622 12776
rect 7760 12773 7788 12872
rect 7926 12860 7932 12872
rect 7984 12860 7990 12912
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12832 9459 12835
rect 9766 12832 9772 12844
rect 9447 12804 9772 12832
rect 9447 12801 9459 12804
rect 9401 12795 9459 12801
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 12618 12832 12624 12844
rect 12176 12804 12624 12832
rect 7653 12767 7711 12773
rect 7653 12764 7665 12767
rect 7616 12736 7665 12764
rect 7616 12724 7622 12736
rect 7653 12733 7665 12736
rect 7699 12733 7711 12767
rect 7653 12727 7711 12733
rect 7745 12767 7803 12773
rect 7745 12733 7757 12767
rect 7791 12733 7803 12767
rect 7745 12727 7803 12733
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12764 8079 12767
rect 8202 12764 8208 12776
rect 8067 12736 8208 12764
rect 8067 12733 8079 12736
rect 8021 12727 8079 12733
rect 8036 12696 8064 12727
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 11054 12724 11060 12776
rect 11112 12764 11118 12776
rect 12176 12773 12204 12804
rect 12618 12792 12624 12804
rect 12676 12832 12682 12844
rect 14734 12832 14740 12844
rect 12676 12804 14740 12832
rect 12676 12792 12682 12804
rect 14734 12792 14740 12804
rect 14792 12832 14798 12844
rect 14792 12804 17356 12832
rect 14792 12792 14798 12804
rect 11149 12767 11207 12773
rect 11149 12764 11161 12767
rect 11112 12736 11161 12764
rect 11112 12724 11118 12736
rect 11149 12733 11161 12736
rect 11195 12733 11207 12767
rect 11149 12727 11207 12733
rect 12161 12767 12219 12773
rect 12161 12733 12173 12767
rect 12207 12733 12219 12767
rect 12161 12727 12219 12733
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 15105 12767 15163 12773
rect 15105 12764 15117 12767
rect 13872 12736 15117 12764
rect 13872 12724 13878 12736
rect 15105 12733 15117 12736
rect 15151 12733 15163 12767
rect 15105 12727 15163 12733
rect 16574 12724 16580 12776
rect 16632 12764 16638 12776
rect 16945 12767 17003 12773
rect 16945 12764 16957 12767
rect 16632 12736 16957 12764
rect 16632 12724 16638 12736
rect 16945 12733 16957 12736
rect 16991 12733 17003 12767
rect 17126 12764 17132 12776
rect 17087 12736 17132 12764
rect 16945 12727 17003 12733
rect 17126 12724 17132 12736
rect 17184 12724 17190 12776
rect 17328 12773 17356 12804
rect 17313 12767 17371 12773
rect 17313 12733 17325 12767
rect 17359 12733 17371 12767
rect 17313 12727 17371 12733
rect 7300 12668 8064 12696
rect 9493 12699 9551 12705
rect 9493 12665 9505 12699
rect 9539 12696 9551 12699
rect 11238 12696 11244 12708
rect 9539 12668 11244 12696
rect 9539 12665 9551 12668
rect 9493 12659 9551 12665
rect 11238 12656 11244 12668
rect 11296 12656 11302 12708
rect 11974 12656 11980 12708
rect 12032 12696 12038 12708
rect 12253 12699 12311 12705
rect 12253 12696 12265 12699
rect 12032 12668 12265 12696
rect 12032 12656 12038 12668
rect 12253 12665 12265 12668
rect 12299 12696 12311 12699
rect 13262 12696 13268 12708
rect 12299 12668 13268 12696
rect 12299 12665 12311 12668
rect 12253 12659 12311 12665
rect 13262 12656 13268 12668
rect 13320 12696 13326 12708
rect 16592 12696 16620 12724
rect 13320 12668 16620 12696
rect 17221 12699 17279 12705
rect 13320 12656 13326 12668
rect 17221 12665 17233 12699
rect 17267 12696 17279 12699
rect 18046 12696 18052 12708
rect 17267 12668 18052 12696
rect 17267 12665 17279 12668
rect 17221 12659 17279 12665
rect 18046 12656 18052 12668
rect 18104 12656 18110 12708
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4801 12631 4859 12637
rect 4801 12628 4813 12631
rect 4212 12600 4813 12628
rect 4212 12588 4218 12600
rect 4801 12597 4813 12600
rect 4847 12597 4859 12631
rect 4801 12591 4859 12597
rect 6822 12588 6828 12640
rect 6880 12628 6886 12640
rect 7009 12631 7067 12637
rect 7009 12628 7021 12631
rect 6880 12600 7021 12628
rect 6880 12588 6886 12600
rect 7009 12597 7021 12600
rect 7055 12597 7067 12631
rect 7009 12591 7067 12597
rect 9401 12631 9459 12637
rect 9401 12597 9413 12631
rect 9447 12628 9459 12631
rect 10502 12628 10508 12640
rect 9447 12600 10508 12628
rect 9447 12597 9459 12600
rect 9401 12591 9459 12597
rect 10502 12588 10508 12600
rect 10560 12588 10566 12640
rect 17494 12628 17500 12640
rect 17455 12600 17500 12628
rect 17494 12588 17500 12600
rect 17552 12588 17558 12640
rect 1104 12538 19044 12560
rect 1104 12486 6962 12538
rect 7014 12486 7026 12538
rect 7078 12486 7090 12538
rect 7142 12486 7154 12538
rect 7206 12486 12942 12538
rect 12994 12486 13006 12538
rect 13058 12486 13070 12538
rect 13122 12486 13134 12538
rect 13186 12486 19044 12538
rect 1104 12464 19044 12486
rect 1596 12396 2774 12424
rect 1596 12365 1624 12396
rect 1581 12359 1639 12365
rect 1581 12325 1593 12359
rect 1627 12325 1639 12359
rect 1581 12319 1639 12325
rect 1486 12084 1492 12096
rect 1447 12056 1492 12084
rect 1486 12044 1492 12056
rect 1544 12044 1550 12096
rect 2746 12084 2774 12396
rect 4154 12384 4160 12436
rect 4212 12384 4218 12436
rect 5350 12384 5356 12436
rect 5408 12424 5414 12436
rect 5813 12427 5871 12433
rect 5813 12424 5825 12427
rect 5408 12396 5825 12424
rect 5408 12384 5414 12396
rect 5813 12393 5825 12396
rect 5859 12393 5871 12427
rect 6270 12424 6276 12436
rect 6231 12396 6276 12424
rect 5813 12387 5871 12393
rect 2866 12356 2872 12368
rect 2827 12328 2872 12356
rect 2866 12316 2872 12328
rect 2924 12316 2930 12368
rect 4172 12356 4200 12384
rect 4341 12359 4399 12365
rect 4341 12356 4353 12359
rect 4172 12328 4353 12356
rect 4341 12325 4353 12328
rect 4387 12325 4399 12359
rect 4341 12319 4399 12325
rect 5074 12316 5080 12368
rect 5132 12316 5138 12368
rect 5828 12356 5856 12387
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 16298 12384 16304 12436
rect 16356 12424 16362 12436
rect 16356 12396 16988 12424
rect 16356 12384 16362 12396
rect 11054 12356 11060 12368
rect 5828 12328 6224 12356
rect 2958 12248 2964 12300
rect 3016 12288 3022 12300
rect 6196 12297 6224 12328
rect 7760 12328 11060 12356
rect 7760 12300 7788 12328
rect 11054 12316 11060 12328
rect 11112 12356 11118 12368
rect 12897 12359 12955 12365
rect 11112 12328 12434 12356
rect 11112 12316 11118 12328
rect 3053 12291 3111 12297
rect 3053 12288 3065 12291
rect 3016 12260 3065 12288
rect 3016 12248 3022 12260
rect 3053 12257 3065 12260
rect 3099 12257 3111 12291
rect 3053 12251 3111 12257
rect 6181 12291 6239 12297
rect 6181 12257 6193 12291
rect 6227 12288 6239 12291
rect 6227 12260 6776 12288
rect 6227 12257 6239 12260
rect 6181 12251 6239 12257
rect 4065 12223 4123 12229
rect 4065 12189 4077 12223
rect 4111 12220 4123 12223
rect 5534 12220 5540 12232
rect 4111 12192 5540 12220
rect 4111 12189 4123 12192
rect 4065 12183 4123 12189
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 6748 12220 6776 12260
rect 7006 12248 7012 12300
rect 7064 12288 7070 12300
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 7064 12260 7481 12288
rect 7064 12248 7070 12260
rect 7469 12257 7481 12260
rect 7515 12288 7527 12291
rect 7742 12288 7748 12300
rect 7515 12260 7748 12288
rect 7515 12257 7527 12260
rect 7469 12251 7527 12257
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 9122 12248 9128 12300
rect 9180 12288 9186 12300
rect 10505 12291 10563 12297
rect 10505 12288 10517 12291
rect 9180 12260 10517 12288
rect 9180 12248 9186 12260
rect 10505 12257 10517 12260
rect 10551 12288 10563 12291
rect 11146 12288 11152 12300
rect 10551 12260 11152 12288
rect 10551 12257 10563 12260
rect 10505 12251 10563 12257
rect 11146 12248 11152 12260
rect 11204 12288 11210 12300
rect 11882 12288 11888 12300
rect 11204 12260 11888 12288
rect 11204 12248 11210 12260
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 9306 12220 9312 12232
rect 6748 12192 9312 12220
rect 9306 12180 9312 12192
rect 9364 12180 9370 12232
rect 12406 12220 12434 12328
rect 12897 12325 12909 12359
rect 12943 12356 12955 12359
rect 13814 12356 13820 12368
rect 12943 12328 13820 12356
rect 12943 12325 12955 12328
rect 12897 12319 12955 12325
rect 13814 12316 13820 12328
rect 13872 12356 13878 12368
rect 14182 12356 14188 12368
rect 13872 12328 14188 12356
rect 13872 12316 13878 12328
rect 14182 12316 14188 12328
rect 14240 12316 14246 12368
rect 12618 12248 12624 12300
rect 12676 12297 12682 12300
rect 12676 12291 12725 12297
rect 12676 12257 12679 12291
rect 12713 12257 12725 12291
rect 12802 12288 12808 12300
rect 12763 12260 12808 12288
rect 12676 12251 12725 12257
rect 12676 12248 12682 12251
rect 12802 12248 12808 12260
rect 12860 12248 12866 12300
rect 13081 12291 13139 12297
rect 13081 12257 13093 12291
rect 13127 12288 13139 12291
rect 13262 12288 13268 12300
rect 13127 12260 13268 12288
rect 13127 12257 13139 12260
rect 13081 12251 13139 12257
rect 13262 12248 13268 12260
rect 13320 12248 13326 12300
rect 13357 12291 13415 12297
rect 13357 12257 13369 12291
rect 13403 12288 13415 12291
rect 15289 12291 15347 12297
rect 15289 12288 15301 12291
rect 13403 12260 15301 12288
rect 13403 12257 13415 12260
rect 13357 12251 13415 12257
rect 15289 12257 15301 12260
rect 15335 12288 15347 12291
rect 16850 12288 16856 12300
rect 15335 12260 16856 12288
rect 15335 12257 15347 12260
rect 15289 12251 15347 12257
rect 13372 12220 13400 12251
rect 16850 12248 16856 12260
rect 16908 12248 16914 12300
rect 16960 12297 16988 12396
rect 18046 12384 18052 12436
rect 18104 12424 18110 12436
rect 18693 12427 18751 12433
rect 18693 12424 18705 12427
rect 18104 12396 18705 12424
rect 18104 12384 18110 12396
rect 18693 12393 18705 12396
rect 18739 12393 18751 12427
rect 18693 12387 18751 12393
rect 17221 12359 17279 12365
rect 17221 12325 17233 12359
rect 17267 12356 17279 12359
rect 17494 12356 17500 12368
rect 17267 12328 17500 12356
rect 17267 12325 17279 12328
rect 17221 12319 17279 12325
rect 17494 12316 17500 12328
rect 17552 12316 17558 12368
rect 18230 12316 18236 12368
rect 18288 12316 18294 12368
rect 16945 12291 17003 12297
rect 16945 12257 16957 12291
rect 16991 12257 17003 12291
rect 16945 12251 17003 12257
rect 12406 12192 13400 12220
rect 12728 12164 12756 12192
rect 12710 12112 12716 12164
rect 12768 12112 12774 12164
rect 4890 12084 4896 12096
rect 2746 12056 4896 12084
rect 4890 12044 4896 12056
rect 4948 12044 4954 12096
rect 7650 12084 7656 12096
rect 7611 12056 7656 12084
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 9490 12044 9496 12096
rect 9548 12084 9554 12096
rect 10597 12087 10655 12093
rect 10597 12084 10609 12087
rect 9548 12056 10609 12084
rect 9548 12044 9554 12056
rect 10597 12053 10609 12056
rect 10643 12053 10655 12087
rect 10597 12047 10655 12053
rect 12529 12087 12587 12093
rect 12529 12053 12541 12087
rect 12575 12084 12587 12087
rect 12618 12084 12624 12096
rect 12575 12056 12624 12084
rect 12575 12053 12587 12056
rect 12529 12047 12587 12053
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 13541 12087 13599 12093
rect 13541 12053 13553 12087
rect 13587 12084 13599 12087
rect 13630 12084 13636 12096
rect 13587 12056 13636 12084
rect 13587 12053 13599 12056
rect 13541 12047 13599 12053
rect 13630 12044 13636 12056
rect 13688 12044 13694 12096
rect 14918 12044 14924 12096
rect 14976 12084 14982 12096
rect 15105 12087 15163 12093
rect 15105 12084 15117 12087
rect 14976 12056 15117 12084
rect 14976 12044 14982 12056
rect 15105 12053 15117 12056
rect 15151 12053 15163 12087
rect 15105 12047 15163 12053
rect 1104 11994 19044 12016
rect 1104 11942 3972 11994
rect 4024 11942 4036 11994
rect 4088 11942 4100 11994
rect 4152 11942 4164 11994
rect 4216 11942 9952 11994
rect 10004 11942 10016 11994
rect 10068 11942 10080 11994
rect 10132 11942 10144 11994
rect 10196 11942 15932 11994
rect 15984 11942 15996 11994
rect 16048 11942 16060 11994
rect 16112 11942 16124 11994
rect 16176 11942 19044 11994
rect 1104 11920 19044 11942
rect 2869 11883 2927 11889
rect 2869 11849 2881 11883
rect 2915 11880 2927 11883
rect 2958 11880 2964 11892
rect 2915 11852 2964 11880
rect 2915 11849 2927 11852
rect 2869 11843 2927 11849
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 4522 11880 4528 11892
rect 4483 11852 4528 11880
rect 4522 11840 4528 11852
rect 4580 11840 4586 11892
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 5169 11883 5227 11889
rect 5169 11880 5181 11883
rect 5132 11852 5181 11880
rect 5132 11840 5138 11852
rect 5169 11849 5181 11852
rect 5215 11849 5227 11883
rect 5169 11843 5227 11849
rect 5534 11840 5540 11892
rect 5592 11880 5598 11892
rect 6546 11880 6552 11892
rect 5592 11852 6552 11880
rect 5592 11840 5598 11852
rect 6546 11840 6552 11852
rect 6604 11880 6610 11892
rect 7466 11880 7472 11892
rect 6604 11852 7472 11880
rect 6604 11840 6610 11852
rect 2038 11812 2044 11824
rect 1596 11784 2044 11812
rect 1596 11753 1624 11784
rect 2038 11772 2044 11784
rect 2096 11772 2102 11824
rect 2225 11815 2283 11821
rect 2225 11781 2237 11815
rect 2271 11781 2283 11815
rect 2225 11775 2283 11781
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11713 1639 11747
rect 1762 11744 1768 11756
rect 1723 11716 1768 11744
rect 1581 11707 1639 11713
rect 1762 11704 1768 11716
rect 1820 11704 1826 11756
rect 2240 11744 2268 11775
rect 3329 11747 3387 11753
rect 3329 11744 3341 11747
rect 2240 11716 3341 11744
rect 2332 11685 2360 11716
rect 3329 11713 3341 11716
rect 3375 11713 3387 11747
rect 3329 11707 3387 11713
rect 4801 11747 4859 11753
rect 4801 11713 4813 11747
rect 4847 11744 4859 11747
rect 5074 11744 5080 11756
rect 4847 11716 5080 11744
rect 4847 11713 4859 11716
rect 4801 11707 4859 11713
rect 5074 11704 5080 11716
rect 5132 11704 5138 11756
rect 5442 11744 5448 11756
rect 5276 11716 5448 11744
rect 2317 11679 2375 11685
rect 2317 11645 2329 11679
rect 2363 11645 2375 11679
rect 2866 11676 2872 11688
rect 2827 11648 2872 11676
rect 2317 11639 2375 11645
rect 2866 11636 2872 11648
rect 2924 11636 2930 11688
rect 2958 11636 2964 11688
rect 3016 11676 3022 11688
rect 4709 11679 4767 11685
rect 3016 11648 3061 11676
rect 3016 11636 3022 11648
rect 4709 11645 4721 11679
rect 4755 11645 4767 11679
rect 4709 11639 4767 11645
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11645 4951 11679
rect 4893 11639 4951 11645
rect 4985 11679 5043 11685
rect 4985 11645 4997 11679
rect 5031 11676 5043 11679
rect 5276 11676 5304 11716
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 6656 11753 6684 11852
rect 7466 11840 7472 11852
rect 7524 11840 7530 11892
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 9861 11883 9919 11889
rect 9861 11880 9873 11883
rect 9824 11852 9873 11880
rect 9824 11840 9830 11852
rect 9861 11849 9873 11852
rect 9907 11849 9919 11883
rect 9861 11843 9919 11849
rect 12802 11840 12808 11892
rect 12860 11880 12866 11892
rect 14093 11883 14151 11889
rect 14093 11880 14105 11883
rect 12860 11852 14105 11880
rect 12860 11840 12866 11852
rect 14093 11849 14105 11852
rect 14139 11849 14151 11883
rect 14093 11843 14151 11849
rect 18141 11883 18199 11889
rect 18141 11849 18153 11883
rect 18187 11880 18199 11883
rect 18230 11880 18236 11892
rect 18187 11852 18236 11880
rect 18187 11849 18199 11852
rect 18141 11843 18199 11849
rect 18230 11840 18236 11852
rect 18288 11840 18294 11892
rect 9401 11815 9459 11821
rect 9401 11781 9413 11815
rect 9447 11812 9459 11815
rect 9490 11812 9496 11824
rect 9447 11784 9496 11812
rect 9447 11781 9459 11784
rect 9401 11775 9459 11781
rect 9490 11772 9496 11784
rect 9548 11772 9554 11824
rect 6641 11747 6699 11753
rect 6641 11713 6653 11747
rect 6687 11713 6699 11747
rect 6914 11744 6920 11756
rect 6875 11716 6920 11744
rect 6641 11707 6699 11713
rect 6914 11704 6920 11716
rect 6972 11704 6978 11756
rect 8294 11704 8300 11756
rect 8352 11744 8358 11756
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 8352 11716 9321 11744
rect 8352 11704 8358 11716
rect 9309 11713 9321 11716
rect 9355 11713 9367 11747
rect 12618 11744 12624 11756
rect 12579 11716 12624 11744
rect 9309 11707 9367 11713
rect 5031 11648 5304 11676
rect 5353 11679 5411 11685
rect 5031 11645 5043 11648
rect 4985 11639 5043 11645
rect 5353 11645 5365 11679
rect 5399 11676 5411 11679
rect 5399 11648 6684 11676
rect 5399 11645 5411 11648
rect 5353 11639 5411 11645
rect 1857 11611 1915 11617
rect 1857 11577 1869 11611
rect 1903 11608 1915 11611
rect 4154 11608 4160 11620
rect 1903 11580 4160 11608
rect 1903 11577 1915 11580
rect 1857 11571 1915 11577
rect 4154 11568 4160 11580
rect 4212 11568 4218 11620
rect 4724 11608 4752 11639
rect 4798 11608 4804 11620
rect 4724 11580 4804 11608
rect 4798 11568 4804 11580
rect 4856 11568 4862 11620
rect 4908 11608 4936 11639
rect 6362 11608 6368 11620
rect 4908 11580 6368 11608
rect 6362 11568 6368 11580
rect 6420 11568 6426 11620
rect 6656 11608 6684 11648
rect 8202 11636 8208 11688
rect 8260 11676 8266 11688
rect 8662 11676 8668 11688
rect 8260 11648 8668 11676
rect 8260 11636 8266 11648
rect 8662 11636 8668 11648
rect 8720 11676 8726 11688
rect 9125 11679 9183 11685
rect 9125 11676 9137 11679
rect 8720 11648 9137 11676
rect 8720 11636 8726 11648
rect 9125 11645 9137 11648
rect 9171 11645 9183 11679
rect 9324 11676 9352 11707
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 14182 11744 14188 11756
rect 14143 11716 14188 11744
rect 14182 11704 14188 11716
rect 14240 11704 14246 11756
rect 15286 11704 15292 11756
rect 15344 11744 15350 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15344 11716 15945 11744
rect 15344 11704 15350 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 9398 11676 9404 11688
rect 9324 11648 9404 11676
rect 9125 11639 9183 11645
rect 9398 11636 9404 11648
rect 9456 11636 9462 11688
rect 9493 11679 9551 11685
rect 9493 11645 9505 11679
rect 9539 11645 9551 11679
rect 9493 11639 9551 11645
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11676 9643 11679
rect 9766 11676 9772 11688
rect 9631 11648 9772 11676
rect 9631 11645 9643 11648
rect 9585 11639 9643 11645
rect 7006 11608 7012 11620
rect 6656 11580 7012 11608
rect 7006 11568 7012 11580
rect 7064 11568 7070 11620
rect 7650 11568 7656 11620
rect 7708 11568 7714 11620
rect 8312 11580 8616 11608
rect 4706 11500 4712 11552
rect 4764 11540 4770 11552
rect 8312 11540 8340 11580
rect 4764 11512 8340 11540
rect 8389 11543 8447 11549
rect 4764 11500 4770 11512
rect 8389 11509 8401 11543
rect 8435 11540 8447 11543
rect 8478 11540 8484 11552
rect 8435 11512 8484 11540
rect 8435 11509 8447 11512
rect 8389 11503 8447 11509
rect 8478 11500 8484 11512
rect 8536 11500 8542 11552
rect 8588 11540 8616 11580
rect 9306 11568 9312 11620
rect 9364 11608 9370 11620
rect 9508 11608 9536 11639
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 12345 11679 12403 11685
rect 12345 11676 12357 11679
rect 12268 11648 12357 11676
rect 9364 11580 9536 11608
rect 9364 11568 9370 11580
rect 10410 11568 10416 11620
rect 10468 11608 10474 11620
rect 12268 11608 12296 11648
rect 12345 11645 12357 11648
rect 12391 11645 12403 11679
rect 16209 11679 16267 11685
rect 12345 11639 12403 11645
rect 13924 11648 14320 11676
rect 12526 11608 12532 11620
rect 10468 11580 12532 11608
rect 10468 11568 10474 11580
rect 12526 11568 12532 11580
rect 12584 11568 12590 11620
rect 13630 11568 13636 11620
rect 13688 11568 13694 11620
rect 13924 11540 13952 11648
rect 8588 11512 13952 11540
rect 14292 11540 14320 11648
rect 16209 11645 16221 11679
rect 16255 11676 16267 11679
rect 16298 11676 16304 11688
rect 16255 11648 16304 11676
rect 16255 11645 16267 11648
rect 16209 11639 16267 11645
rect 14918 11568 14924 11620
rect 14976 11568 14982 11620
rect 16022 11568 16028 11620
rect 16080 11608 16086 11620
rect 16224 11608 16252 11639
rect 16298 11636 16304 11648
rect 16356 11636 16362 11688
rect 16850 11636 16856 11688
rect 16908 11676 16914 11688
rect 17037 11679 17095 11685
rect 17037 11676 17049 11679
rect 16908 11648 17049 11676
rect 16908 11636 16914 11648
rect 17037 11645 17049 11648
rect 17083 11676 17095 11679
rect 17957 11679 18015 11685
rect 17957 11676 17969 11679
rect 17083 11648 17969 11676
rect 17083 11645 17095 11648
rect 17037 11639 17095 11645
rect 17957 11645 17969 11648
rect 18003 11645 18015 11679
rect 18690 11676 18696 11688
rect 18651 11648 18696 11676
rect 17957 11639 18015 11645
rect 18690 11636 18696 11648
rect 18748 11636 18754 11688
rect 16080 11580 16252 11608
rect 16546 11580 18552 11608
rect 16080 11568 16086 11580
rect 16546 11540 16574 11580
rect 14292 11512 16574 11540
rect 17126 11500 17132 11552
rect 17184 11540 17190 11552
rect 18524 11549 18552 11580
rect 17221 11543 17279 11549
rect 17221 11540 17233 11543
rect 17184 11512 17233 11540
rect 17184 11500 17190 11512
rect 17221 11509 17233 11512
rect 17267 11509 17279 11543
rect 17221 11503 17279 11509
rect 18509 11543 18567 11549
rect 18509 11509 18521 11543
rect 18555 11509 18567 11543
rect 18509 11503 18567 11509
rect 1104 11450 19044 11472
rect 1104 11398 6962 11450
rect 7014 11398 7026 11450
rect 7078 11398 7090 11450
rect 7142 11398 7154 11450
rect 7206 11398 12942 11450
rect 12994 11398 13006 11450
rect 13058 11398 13070 11450
rect 13122 11398 13134 11450
rect 13186 11398 19044 11450
rect 1104 11376 19044 11398
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 2958 11336 2964 11348
rect 2915 11308 2964 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 4154 11336 4160 11348
rect 4115 11308 4160 11336
rect 4154 11296 4160 11308
rect 4212 11296 4218 11348
rect 4982 11296 4988 11348
rect 5040 11336 5046 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 5040 11308 5181 11336
rect 5040 11296 5046 11308
rect 5169 11305 5181 11308
rect 5215 11336 5227 11339
rect 8202 11336 8208 11348
rect 5215 11308 6132 11336
rect 8163 11308 8208 11336
rect 5215 11305 5227 11308
rect 5169 11299 5227 11305
rect 3694 11228 3700 11280
rect 3752 11268 3758 11280
rect 6104 11277 6132 11308
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 12526 11296 12532 11348
rect 12584 11336 12590 11348
rect 13722 11336 13728 11348
rect 12584 11308 13728 11336
rect 12584 11296 12590 11308
rect 13722 11296 13728 11308
rect 13780 11296 13786 11348
rect 17310 11296 17316 11348
rect 17368 11336 17374 11348
rect 17865 11339 17923 11345
rect 17865 11336 17877 11339
rect 17368 11308 17877 11336
rect 17368 11296 17374 11308
rect 17865 11305 17877 11308
rect 17911 11305 17923 11339
rect 17865 11299 17923 11305
rect 6089 11271 6147 11277
rect 3752 11240 6040 11268
rect 3752 11228 3758 11240
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 4525 11203 4583 11209
rect 2832 11172 2877 11200
rect 2832 11160 2838 11172
rect 4525 11169 4537 11203
rect 4571 11200 4583 11203
rect 4614 11200 4620 11212
rect 4571 11172 4620 11200
rect 4571 11169 4583 11172
rect 4525 11163 4583 11169
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 5166 11200 5172 11212
rect 5123 11172 5172 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 5166 11160 5172 11172
rect 5224 11160 5230 11212
rect 6012 11200 6040 11240
rect 6089 11237 6101 11271
rect 6135 11237 6147 11271
rect 6270 11268 6276 11280
rect 6231 11240 6276 11268
rect 6089 11231 6147 11237
rect 6270 11228 6276 11240
rect 6328 11228 6334 11280
rect 11333 11271 11391 11277
rect 11333 11268 11345 11271
rect 7576 11240 11345 11268
rect 7576 11200 7604 11240
rect 11333 11237 11345 11240
rect 11379 11237 11391 11271
rect 16390 11268 16396 11280
rect 16351 11240 16396 11268
rect 11333 11231 11391 11237
rect 16390 11228 16396 11240
rect 16448 11228 16454 11280
rect 17126 11228 17132 11280
rect 17184 11228 17190 11280
rect 6012 11172 7604 11200
rect 8113 11203 8171 11209
rect 8113 11169 8125 11203
rect 8159 11200 8171 11203
rect 8478 11200 8484 11212
rect 8159 11172 8484 11200
rect 8159 11169 8171 11172
rect 8113 11163 8171 11169
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11132 4491 11135
rect 5442 11132 5448 11144
rect 4479 11104 5448 11132
rect 4479 11101 4491 11104
rect 4433 11095 4491 11101
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 6362 11092 6368 11144
rect 6420 11132 6426 11144
rect 7558 11132 7564 11144
rect 6420 11104 7564 11132
rect 6420 11092 6426 11104
rect 7558 11092 7564 11104
rect 7616 11132 7622 11144
rect 8128 11132 8156 11163
rect 8478 11160 8484 11172
rect 8536 11200 8542 11212
rect 9214 11200 9220 11212
rect 8536 11172 9220 11200
rect 8536 11160 8542 11172
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 10413 11203 10471 11209
rect 10413 11200 10425 11203
rect 9324 11172 10425 11200
rect 7616 11104 8156 11132
rect 7616 11092 7622 11104
rect 8938 11092 8944 11144
rect 8996 11132 9002 11144
rect 9324 11132 9352 11172
rect 10413 11169 10425 11172
rect 10459 11169 10471 11203
rect 10413 11163 10471 11169
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11169 10655 11203
rect 11422 11200 11428 11212
rect 11383 11172 11428 11200
rect 10597 11163 10655 11169
rect 8996 11104 9352 11132
rect 8996 11092 9002 11104
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 10612 11132 10640 11163
rect 11422 11160 11428 11172
rect 11480 11160 11486 11212
rect 13722 11160 13728 11212
rect 13780 11200 13786 11212
rect 16022 11200 16028 11212
rect 13780 11172 16028 11200
rect 13780 11160 13786 11172
rect 16022 11160 16028 11172
rect 16080 11200 16086 11212
rect 16117 11203 16175 11209
rect 16117 11200 16129 11203
rect 16080 11172 16129 11200
rect 16080 11160 16086 11172
rect 16117 11169 16129 11172
rect 16163 11169 16175 11203
rect 16117 11163 16175 11169
rect 9732 11104 10640 11132
rect 11241 11135 11299 11141
rect 9732 11092 9738 11104
rect 11241 11101 11253 11135
rect 11287 11132 11299 11135
rect 11330 11132 11336 11144
rect 11287 11104 11336 11132
rect 11287 11101 11299 11104
rect 11241 11095 11299 11101
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 6457 11067 6515 11073
rect 6457 11033 6469 11067
rect 6503 11064 6515 11067
rect 8478 11064 8484 11076
rect 6503 11036 8484 11064
rect 6503 11033 6515 11036
rect 6457 11027 6515 11033
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 10781 11067 10839 11073
rect 10781 11033 10793 11067
rect 10827 11064 10839 11067
rect 11054 11064 11060 11076
rect 10827 11036 11060 11064
rect 10827 11033 10839 11036
rect 10781 11027 10839 11033
rect 11054 11024 11060 11036
rect 11112 11024 11118 11076
rect 11793 11067 11851 11073
rect 11793 11033 11805 11067
rect 11839 11064 11851 11067
rect 12618 11064 12624 11076
rect 11839 11036 12624 11064
rect 11839 11033 11851 11036
rect 11793 11027 11851 11033
rect 12618 11024 12624 11036
rect 12676 11024 12682 11076
rect 4525 10999 4583 11005
rect 4525 10965 4537 10999
rect 4571 10996 4583 10999
rect 5350 10996 5356 11008
rect 4571 10968 5356 10996
rect 4571 10965 4583 10968
rect 4525 10959 4583 10965
rect 5350 10956 5356 10968
rect 5408 10956 5414 11008
rect 10318 10956 10324 11008
rect 10376 10996 10382 11008
rect 15470 10996 15476 11008
rect 10376 10968 15476 10996
rect 10376 10956 10382 10968
rect 15470 10956 15476 10968
rect 15528 10956 15534 11008
rect 1104 10906 19044 10928
rect 1104 10854 3972 10906
rect 4024 10854 4036 10906
rect 4088 10854 4100 10906
rect 4152 10854 4164 10906
rect 4216 10854 9952 10906
rect 10004 10854 10016 10906
rect 10068 10854 10080 10906
rect 10132 10854 10144 10906
rect 10196 10854 15932 10906
rect 15984 10854 15996 10906
rect 16048 10854 16060 10906
rect 16112 10854 16124 10906
rect 16176 10854 19044 10906
rect 1104 10832 19044 10854
rect 4798 10752 4804 10804
rect 4856 10792 4862 10804
rect 4893 10795 4951 10801
rect 4893 10792 4905 10795
rect 4856 10764 4905 10792
rect 4856 10752 4862 10764
rect 4893 10761 4905 10764
rect 4939 10761 4951 10795
rect 6178 10792 6184 10804
rect 6139 10764 6184 10792
rect 4893 10755 4951 10761
rect 6178 10752 6184 10764
rect 6236 10752 6242 10804
rect 6733 10795 6791 10801
rect 6733 10761 6745 10795
rect 6779 10761 6791 10795
rect 7282 10792 7288 10804
rect 7243 10764 7288 10792
rect 6733 10755 6791 10761
rect 4614 10684 4620 10736
rect 4672 10724 4678 10736
rect 6748 10724 6776 10755
rect 7282 10752 7288 10764
rect 7340 10792 7346 10804
rect 8481 10795 8539 10801
rect 8481 10792 8493 10795
rect 7340 10764 8493 10792
rect 7340 10752 7346 10764
rect 8481 10761 8493 10764
rect 8527 10761 8539 10795
rect 9585 10795 9643 10801
rect 9585 10792 9597 10795
rect 8481 10755 8539 10761
rect 8588 10764 9597 10792
rect 8588 10724 8616 10764
rect 9585 10761 9597 10764
rect 9631 10792 9643 10795
rect 9674 10792 9680 10804
rect 9631 10764 9680 10792
rect 9631 10761 9643 10764
rect 9585 10755 9643 10761
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 9953 10795 10011 10801
rect 9953 10761 9965 10795
rect 9999 10792 10011 10795
rect 10318 10792 10324 10804
rect 9999 10764 10324 10792
rect 9999 10761 10011 10764
rect 9953 10755 10011 10761
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 11422 10752 11428 10804
rect 11480 10792 11486 10804
rect 11701 10795 11759 10801
rect 11701 10792 11713 10795
rect 11480 10764 11713 10792
rect 11480 10752 11486 10764
rect 11701 10761 11713 10764
rect 11747 10761 11759 10795
rect 11701 10755 11759 10761
rect 4672 10696 6776 10724
rect 7944 10696 8616 10724
rect 8849 10727 8907 10733
rect 4672 10684 4678 10696
rect 4798 10616 4804 10668
rect 4856 10656 4862 10668
rect 7944 10656 7972 10696
rect 8849 10693 8861 10727
rect 8895 10724 8907 10727
rect 11146 10724 11152 10736
rect 8895 10696 10732 10724
rect 8895 10693 8907 10696
rect 8849 10687 8907 10693
rect 9398 10656 9404 10668
rect 4856 10628 7972 10656
rect 8680 10628 9260 10656
rect 9359 10628 9404 10656
rect 4856 10616 4862 10628
rect 4617 10591 4675 10597
rect 4617 10557 4629 10591
rect 4663 10588 4675 10591
rect 5166 10588 5172 10600
rect 4663 10560 5172 10588
rect 4663 10557 4675 10560
rect 4617 10551 4675 10557
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 6104 10597 6132 10628
rect 8680 10600 8708 10628
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10557 6147 10591
rect 6089 10551 6147 10557
rect 6362 10548 6368 10600
rect 6420 10588 6426 10600
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 6420 10560 6653 10588
rect 6420 10548 6426 10560
rect 6641 10557 6653 10560
rect 6687 10588 6699 10591
rect 6730 10588 6736 10600
rect 6687 10560 6736 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 6730 10548 6736 10560
rect 6788 10548 6794 10600
rect 7193 10591 7251 10597
rect 7193 10557 7205 10591
rect 7239 10557 7251 10591
rect 7193 10551 7251 10557
rect 4801 10523 4859 10529
rect 4801 10489 4813 10523
rect 4847 10489 4859 10523
rect 4801 10483 4859 10489
rect 4816 10452 4844 10483
rect 5074 10480 5080 10532
rect 5132 10520 5138 10532
rect 6457 10523 6515 10529
rect 6457 10520 6469 10523
rect 5132 10492 6469 10520
rect 5132 10480 5138 10492
rect 6457 10489 6469 10492
rect 6503 10520 6515 10523
rect 7208 10520 7236 10551
rect 7834 10548 7840 10600
rect 7892 10588 7898 10600
rect 8113 10591 8171 10597
rect 8113 10588 8125 10591
rect 7892 10560 8125 10588
rect 7892 10548 7898 10560
rect 8113 10557 8125 10560
rect 8159 10557 8171 10591
rect 8294 10588 8300 10600
rect 8255 10560 8300 10588
rect 8113 10551 8171 10557
rect 8018 10520 8024 10532
rect 6503 10492 8024 10520
rect 6503 10489 6515 10492
rect 6457 10483 6515 10489
rect 8018 10480 8024 10492
rect 8076 10480 8082 10532
rect 8128 10520 8156 10551
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 8478 10588 8484 10600
rect 8439 10560 8484 10588
rect 8478 10548 8484 10560
rect 8536 10548 8542 10600
rect 8662 10588 8668 10600
rect 8623 10560 8668 10588
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 8938 10548 8944 10600
rect 8996 10588 9002 10600
rect 9232 10597 9260 10628
rect 9398 10616 9404 10628
rect 9456 10616 9462 10668
rect 9125 10591 9183 10597
rect 9125 10588 9137 10591
rect 8996 10560 9137 10588
rect 8996 10548 9002 10560
rect 9125 10557 9137 10560
rect 9171 10557 9183 10591
rect 9125 10551 9183 10557
rect 9217 10591 9275 10597
rect 9217 10557 9229 10591
rect 9263 10557 9275 10591
rect 9217 10551 9275 10557
rect 9490 10548 9496 10600
rect 9548 10588 9554 10600
rect 9677 10591 9735 10597
rect 9548 10560 9593 10588
rect 9548 10548 9554 10560
rect 9677 10557 9689 10591
rect 9723 10588 9735 10591
rect 9766 10588 9772 10600
rect 9723 10560 9772 10588
rect 9723 10557 9735 10560
rect 9677 10551 9735 10557
rect 9766 10548 9772 10560
rect 9824 10548 9830 10600
rect 10704 10597 10732 10696
rect 10888 10696 11152 10724
rect 10888 10665 10916 10696
rect 11146 10684 11152 10696
rect 11204 10684 11210 10736
rect 11517 10727 11575 10733
rect 11517 10693 11529 10727
rect 11563 10724 11575 10727
rect 14366 10724 14372 10736
rect 11563 10696 12112 10724
rect 11563 10693 11575 10696
rect 11517 10687 11575 10693
rect 10873 10659 10931 10665
rect 10873 10625 10885 10659
rect 10919 10625 10931 10659
rect 11054 10656 11060 10668
rect 11015 10628 11060 10656
rect 10873 10619 10931 10625
rect 11054 10616 11060 10628
rect 11112 10656 11118 10668
rect 12084 10665 12112 10696
rect 13464 10696 14372 10724
rect 13464 10665 13492 10696
rect 14366 10684 14372 10696
rect 14424 10684 14430 10736
rect 12069 10659 12127 10665
rect 11112 10628 12020 10656
rect 11112 10616 11118 10628
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10557 10563 10591
rect 10505 10551 10563 10557
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10588 10747 10591
rect 11149 10591 11207 10597
rect 11149 10588 11161 10591
rect 10735 10560 11161 10588
rect 10735 10557 10747 10560
rect 10689 10551 10747 10557
rect 11149 10557 11161 10560
rect 11195 10557 11207 10591
rect 11149 10551 11207 10557
rect 11885 10591 11943 10597
rect 11885 10557 11897 10591
rect 11931 10557 11943 10591
rect 11992 10588 12020 10628
rect 12069 10625 12081 10659
rect 12115 10625 12127 10659
rect 12069 10619 12127 10625
rect 13449 10659 13507 10665
rect 13449 10625 13461 10659
rect 13495 10625 13507 10659
rect 13630 10656 13636 10668
rect 13591 10628 13636 10656
rect 13449 10619 13507 10625
rect 13630 10616 13636 10628
rect 13688 10616 13694 10668
rect 12437 10591 12495 10597
rect 12437 10588 12449 10591
rect 11992 10560 12449 10588
rect 11885 10551 11943 10557
rect 12437 10557 12449 10560
rect 12483 10557 12495 10591
rect 12437 10551 12495 10557
rect 9033 10523 9091 10529
rect 9033 10520 9045 10523
rect 8128 10492 9045 10520
rect 9033 10489 9045 10492
rect 9079 10489 9091 10523
rect 9508 10520 9536 10548
rect 10520 10520 10548 10551
rect 11900 10520 11928 10551
rect 12710 10548 12716 10600
rect 12768 10588 12774 10600
rect 15013 10591 15071 10597
rect 12768 10560 13952 10588
rect 12768 10548 12774 10560
rect 9508 10492 10548 10520
rect 10612 10492 11928 10520
rect 12621 10523 12679 10529
rect 9033 10483 9091 10489
rect 10612 10464 10640 10492
rect 12621 10489 12633 10523
rect 12667 10489 12679 10523
rect 12621 10483 12679 10489
rect 12805 10523 12863 10529
rect 12805 10489 12817 10523
rect 12851 10520 12863 10523
rect 13357 10523 13415 10529
rect 13357 10520 13369 10523
rect 12851 10492 13369 10520
rect 12851 10489 12863 10492
rect 12805 10483 12863 10489
rect 13357 10489 13369 10492
rect 13403 10489 13415 10523
rect 13924 10520 13952 10560
rect 15013 10557 15025 10591
rect 15059 10588 15071 10591
rect 15102 10588 15108 10600
rect 15059 10560 15108 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 15378 10588 15384 10600
rect 15339 10560 15384 10588
rect 15378 10548 15384 10560
rect 15436 10548 15442 10600
rect 18506 10520 18512 10532
rect 13924 10492 18512 10520
rect 13357 10483 13415 10489
rect 5350 10452 5356 10464
rect 4816 10424 5356 10452
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 8113 10455 8171 10461
rect 8113 10421 8125 10455
rect 8159 10452 8171 10455
rect 8202 10452 8208 10464
rect 8159 10424 8208 10452
rect 8159 10421 8171 10424
rect 8113 10415 8171 10421
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 10594 10452 10600 10464
rect 10555 10424 10600 10452
rect 10594 10412 10600 10424
rect 10652 10412 10658 10464
rect 11146 10412 11152 10464
rect 11204 10452 11210 10464
rect 12342 10452 12348 10464
rect 11204 10424 12348 10452
rect 11204 10412 11210 10424
rect 12342 10412 12348 10424
rect 12400 10452 12406 10464
rect 12636 10452 12664 10483
rect 18506 10480 18512 10492
rect 18564 10480 18570 10532
rect 12400 10424 12664 10452
rect 12989 10455 13047 10461
rect 12400 10412 12406 10424
rect 12989 10421 13001 10455
rect 13035 10452 13047 10455
rect 13262 10452 13268 10464
rect 13035 10424 13268 10452
rect 13035 10421 13047 10424
rect 12989 10415 13047 10421
rect 13262 10412 13268 10424
rect 13320 10412 13326 10464
rect 15381 10455 15439 10461
rect 15381 10421 15393 10455
rect 15427 10452 15439 10455
rect 15746 10452 15752 10464
rect 15427 10424 15752 10452
rect 15427 10421 15439 10424
rect 15381 10415 15439 10421
rect 15746 10412 15752 10424
rect 15804 10412 15810 10464
rect 1104 10362 19044 10384
rect 1104 10310 6962 10362
rect 7014 10310 7026 10362
rect 7078 10310 7090 10362
rect 7142 10310 7154 10362
rect 7206 10310 12942 10362
rect 12994 10310 13006 10362
rect 13058 10310 13070 10362
rect 13122 10310 13134 10362
rect 13186 10310 19044 10362
rect 1104 10288 19044 10310
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 3237 10251 3295 10257
rect 3237 10248 3249 10251
rect 2832 10220 3249 10248
rect 2832 10208 2838 10220
rect 3237 10217 3249 10220
rect 3283 10217 3295 10251
rect 4706 10248 4712 10260
rect 4667 10220 4712 10248
rect 3237 10211 3295 10217
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 6546 10208 6552 10260
rect 6604 10248 6610 10260
rect 6825 10251 6883 10257
rect 6825 10248 6837 10251
rect 6604 10220 6837 10248
rect 6604 10208 6610 10220
rect 6825 10217 6837 10220
rect 6871 10217 6883 10251
rect 10855 10251 10913 10257
rect 10855 10248 10867 10251
rect 6825 10211 6883 10217
rect 6932 10220 10867 10248
rect 6932 10180 6960 10220
rect 10855 10217 10867 10220
rect 10901 10217 10913 10251
rect 10855 10211 10913 10217
rect 11333 10251 11391 10257
rect 11333 10217 11345 10251
rect 11379 10248 11391 10251
rect 12710 10248 12716 10260
rect 11379 10220 12716 10248
rect 11379 10217 11391 10220
rect 11333 10211 11391 10217
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 12805 10251 12863 10257
rect 12805 10217 12817 10251
rect 12851 10248 12863 10251
rect 13449 10251 13507 10257
rect 12851 10220 13308 10248
rect 12851 10217 12863 10220
rect 12805 10211 12863 10217
rect 4448 10152 6960 10180
rect 2225 10115 2283 10121
rect 2225 10081 2237 10115
rect 2271 10081 2283 10115
rect 2225 10075 2283 10081
rect 2777 10115 2835 10121
rect 2777 10081 2789 10115
rect 2823 10112 2835 10115
rect 2958 10112 2964 10124
rect 2823 10084 2964 10112
rect 2823 10081 2835 10084
rect 2777 10075 2835 10081
rect 2240 10044 2268 10075
rect 2958 10072 2964 10084
rect 3016 10112 3022 10124
rect 3510 10112 3516 10124
rect 3016 10084 3516 10112
rect 3016 10072 3022 10084
rect 3510 10072 3516 10084
rect 3568 10072 3574 10124
rect 2869 10047 2927 10053
rect 2869 10044 2881 10047
rect 2240 10016 2881 10044
rect 2869 10013 2881 10016
rect 2915 10044 2927 10047
rect 4448 10044 4476 10152
rect 8202 10140 8208 10192
rect 8260 10180 8266 10192
rect 8260 10152 10272 10180
rect 8260 10140 8266 10152
rect 4522 10072 4528 10124
rect 4580 10112 4586 10124
rect 4801 10115 4859 10121
rect 4801 10112 4813 10115
rect 4580 10084 4813 10112
rect 4580 10072 4586 10084
rect 4801 10081 4813 10084
rect 4847 10081 4859 10115
rect 4801 10075 4859 10081
rect 4982 10072 4988 10124
rect 5040 10112 5046 10124
rect 5445 10115 5503 10121
rect 5445 10112 5457 10115
rect 5040 10084 5457 10112
rect 5040 10072 5046 10084
rect 5445 10081 5457 10084
rect 5491 10081 5503 10115
rect 5445 10075 5503 10081
rect 6178 10072 6184 10124
rect 6236 10112 6242 10124
rect 6549 10115 6607 10121
rect 6549 10112 6561 10115
rect 6236 10084 6561 10112
rect 6236 10072 6242 10084
rect 6549 10081 6561 10084
rect 6595 10081 6607 10115
rect 6549 10075 6607 10081
rect 7282 10072 7288 10124
rect 7340 10112 7346 10124
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 7340 10084 9137 10112
rect 7340 10072 7346 10084
rect 9125 10081 9137 10084
rect 9171 10081 9183 10115
rect 9125 10075 9183 10081
rect 9214 10072 9220 10124
rect 9272 10112 9278 10124
rect 9401 10115 9459 10121
rect 9272 10084 9317 10112
rect 9272 10072 9278 10084
rect 9401 10081 9413 10115
rect 9447 10112 9459 10115
rect 9490 10112 9496 10124
rect 9447 10084 9496 10112
rect 9447 10081 9459 10084
rect 9401 10075 9459 10081
rect 2915 10016 4476 10044
rect 4709 10047 4767 10053
rect 2915 10013 2927 10016
rect 2869 10007 2927 10013
rect 4709 10013 4721 10047
rect 4755 10013 4767 10047
rect 4709 10007 4767 10013
rect 2774 9936 2780 9988
rect 2832 9976 2838 9988
rect 3237 9979 3295 9985
rect 2832 9948 2877 9976
rect 2832 9936 2838 9948
rect 3237 9945 3249 9979
rect 3283 9976 3295 9979
rect 3329 9979 3387 9985
rect 3329 9976 3341 9979
rect 3283 9948 3341 9976
rect 3283 9945 3295 9948
rect 3237 9939 3295 9945
rect 3329 9945 3341 9948
rect 3375 9945 3387 9979
rect 4724 9976 4752 10007
rect 5074 10004 5080 10056
rect 5132 10044 5138 10056
rect 5169 10047 5227 10053
rect 5169 10044 5181 10047
rect 5132 10016 5181 10044
rect 5132 10004 5138 10016
rect 5169 10013 5181 10016
rect 5215 10013 5227 10047
rect 5169 10007 5227 10013
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10013 5319 10047
rect 5261 10007 5319 10013
rect 4985 9979 5043 9985
rect 4985 9976 4997 9979
rect 4724 9948 4997 9976
rect 3329 9939 3387 9945
rect 4985 9945 4997 9948
rect 5031 9945 5043 9979
rect 5276 9976 5304 10007
rect 5350 10004 5356 10056
rect 5408 10044 5414 10056
rect 6825 10047 6883 10053
rect 5408 10016 5453 10044
rect 5408 10004 5414 10016
rect 6825 10013 6837 10047
rect 6871 10044 6883 10047
rect 7650 10044 7656 10056
rect 6871 10016 7656 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 8294 10004 8300 10056
rect 8352 10044 8358 10056
rect 9416 10044 9444 10075
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 9674 10072 9680 10124
rect 9732 10112 9738 10124
rect 10244 10121 10272 10152
rect 10594 10140 10600 10192
rect 10652 10180 10658 10192
rect 13280 10189 13308 10220
rect 13449 10217 13461 10251
rect 13495 10248 13507 10251
rect 13538 10248 13544 10260
rect 13495 10220 13544 10248
rect 13495 10217 13507 10220
rect 13449 10211 13507 10217
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 15102 10248 15108 10260
rect 15063 10220 15108 10248
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 15470 10248 15476 10260
rect 15431 10220 15476 10248
rect 15470 10208 15476 10220
rect 15528 10208 15534 10260
rect 15565 10251 15623 10257
rect 15565 10217 15577 10251
rect 15611 10248 15623 10251
rect 16574 10248 16580 10260
rect 15611 10220 16580 10248
rect 15611 10217 15623 10220
rect 15565 10211 15623 10217
rect 16574 10208 16580 10220
rect 16632 10208 16638 10260
rect 17037 10251 17095 10257
rect 17037 10217 17049 10251
rect 17083 10248 17095 10251
rect 17954 10248 17960 10260
rect 17083 10220 17960 10248
rect 17083 10217 17095 10220
rect 17037 10211 17095 10217
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 11149 10183 11207 10189
rect 11149 10180 11161 10183
rect 10652 10152 11161 10180
rect 10652 10140 10658 10152
rect 11149 10149 11161 10152
rect 11195 10149 11207 10183
rect 13265 10183 13323 10189
rect 11149 10143 11207 10149
rect 11440 10152 12940 10180
rect 9861 10115 9919 10121
rect 9861 10112 9873 10115
rect 9732 10084 9873 10112
rect 9732 10072 9738 10084
rect 9861 10081 9873 10084
rect 9907 10112 9919 10115
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 9907 10084 10057 10112
rect 9907 10081 9919 10084
rect 9861 10075 9919 10081
rect 10045 10081 10057 10084
rect 10091 10081 10103 10115
rect 10045 10075 10103 10081
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10081 10287 10115
rect 10229 10075 10287 10081
rect 11440 10056 11468 10152
rect 12342 10072 12348 10124
rect 12400 10112 12406 10124
rect 12621 10115 12679 10121
rect 12621 10112 12633 10115
rect 12400 10084 12633 10112
rect 12400 10072 12406 10084
rect 12621 10081 12633 10084
rect 12667 10081 12679 10115
rect 12912 10112 12940 10152
rect 13265 10149 13277 10183
rect 13311 10149 13323 10183
rect 13265 10143 13323 10149
rect 13541 10115 13599 10121
rect 13541 10112 13553 10115
rect 12912 10084 13553 10112
rect 12621 10075 12679 10081
rect 13541 10081 13553 10084
rect 13587 10112 13599 10115
rect 13630 10112 13636 10124
rect 13587 10084 13636 10112
rect 13587 10081 13599 10084
rect 13541 10075 13599 10081
rect 13630 10072 13636 10084
rect 13688 10072 13694 10124
rect 14461 10115 14519 10121
rect 14461 10081 14473 10115
rect 14507 10112 14519 10115
rect 14550 10112 14556 10124
rect 14507 10084 14556 10112
rect 14507 10081 14519 10084
rect 14461 10075 14519 10081
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 15013 10115 15071 10121
rect 15013 10081 15025 10115
rect 15059 10112 15071 10115
rect 15102 10112 15108 10124
rect 15059 10084 15108 10112
rect 15059 10081 15071 10084
rect 15013 10075 15071 10081
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 17129 10115 17187 10121
rect 17129 10081 17141 10115
rect 17175 10081 17187 10115
rect 17129 10075 17187 10081
rect 8352 10016 9444 10044
rect 8352 10004 8358 10016
rect 9582 10004 9588 10056
rect 9640 10044 9646 10056
rect 9953 10047 10011 10053
rect 9953 10044 9965 10047
rect 9640 10016 9965 10044
rect 9640 10004 9646 10016
rect 9953 10013 9965 10016
rect 9999 10013 10011 10047
rect 11422 10044 11428 10056
rect 11383 10016 11428 10044
rect 9953 10007 10011 10013
rect 11422 10004 11428 10016
rect 11480 10004 11486 10056
rect 13648 10044 13676 10072
rect 15657 10047 15715 10053
rect 15657 10044 15669 10047
rect 13648 10016 15669 10044
rect 15657 10013 15669 10016
rect 15703 10044 15715 10047
rect 16853 10047 16911 10053
rect 16853 10044 16865 10047
rect 15703 10016 16865 10044
rect 15703 10013 15715 10016
rect 15657 10007 15715 10013
rect 16853 10013 16865 10016
rect 16899 10013 16911 10047
rect 16853 10007 16911 10013
rect 4985 9939 5043 9945
rect 5184 9948 5304 9976
rect 10413 9979 10471 9985
rect 5184 9920 5212 9948
rect 10413 9945 10425 9979
rect 10459 9976 10471 9979
rect 10459 9948 16574 9976
rect 10459 9945 10471 9948
rect 10413 9939 10471 9945
rect 4249 9911 4307 9917
rect 4249 9877 4261 9911
rect 4295 9908 4307 9911
rect 4430 9908 4436 9920
rect 4295 9880 4436 9908
rect 4295 9877 4307 9880
rect 4249 9871 4307 9877
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 5166 9868 5172 9920
rect 5224 9868 5230 9920
rect 6638 9908 6644 9920
rect 6599 9880 6644 9908
rect 6638 9868 6644 9880
rect 6696 9868 6702 9920
rect 12802 9868 12808 9920
rect 12860 9908 12866 9920
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 12860 9880 13001 9908
rect 12860 9868 12866 9880
rect 12989 9877 13001 9880
rect 13035 9877 13047 9911
rect 12989 9871 13047 9877
rect 14461 9911 14519 9917
rect 14461 9877 14473 9911
rect 14507 9908 14519 9911
rect 15746 9908 15752 9920
rect 14507 9880 15752 9908
rect 14507 9877 14519 9880
rect 14461 9871 14519 9877
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 16546 9908 16574 9948
rect 17144 9908 17172 10075
rect 17494 9908 17500 9920
rect 16546 9880 17172 9908
rect 17455 9880 17500 9908
rect 17494 9868 17500 9880
rect 17552 9868 17558 9920
rect 1104 9818 19044 9840
rect 1104 9766 3972 9818
rect 4024 9766 4036 9818
rect 4088 9766 4100 9818
rect 4152 9766 4164 9818
rect 4216 9766 9952 9818
rect 10004 9766 10016 9818
rect 10068 9766 10080 9818
rect 10132 9766 10144 9818
rect 10196 9766 15932 9818
rect 15984 9766 15996 9818
rect 16048 9766 16060 9818
rect 16112 9766 16124 9818
rect 16176 9766 19044 9818
rect 1104 9744 19044 9766
rect 4614 9664 4620 9716
rect 4672 9704 4678 9716
rect 8938 9704 8944 9716
rect 4672 9676 8944 9704
rect 4672 9664 4678 9676
rect 8938 9664 8944 9676
rect 8996 9664 9002 9716
rect 15378 9664 15384 9716
rect 15436 9704 15442 9716
rect 15473 9707 15531 9713
rect 15473 9704 15485 9707
rect 15436 9676 15485 9704
rect 15436 9664 15442 9676
rect 15473 9673 15485 9676
rect 15519 9673 15531 9707
rect 15473 9667 15531 9673
rect 4522 9636 4528 9648
rect 2056 9608 4528 9636
rect 2056 9580 2084 9608
rect 4522 9596 4528 9608
rect 4580 9596 4586 9648
rect 5258 9636 5264 9648
rect 4724 9608 5264 9636
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9568 1731 9571
rect 2038 9568 2044 9580
rect 1719 9540 2044 9568
rect 1719 9537 1731 9540
rect 1673 9531 1731 9537
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 4724 9577 4752 9608
rect 5258 9596 5264 9608
rect 5316 9596 5322 9648
rect 6270 9596 6276 9648
rect 6328 9636 6334 9648
rect 6733 9639 6791 9645
rect 6733 9636 6745 9639
rect 6328 9608 6745 9636
rect 6328 9596 6334 9608
rect 6733 9605 6745 9608
rect 6779 9605 6791 9639
rect 6733 9599 6791 9605
rect 6917 9639 6975 9645
rect 6917 9605 6929 9639
rect 6963 9636 6975 9639
rect 7282 9636 7288 9648
rect 6963 9608 7288 9636
rect 6963 9605 6975 9608
rect 6917 9599 6975 9605
rect 7282 9596 7288 9608
rect 7340 9636 7346 9648
rect 7650 9636 7656 9648
rect 7340 9608 7420 9636
rect 7611 9608 7656 9636
rect 7340 9596 7346 9608
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9537 4767 9571
rect 4709 9531 4767 9537
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9568 4859 9571
rect 5074 9568 5080 9580
rect 4847 9540 5080 9568
rect 4847 9537 4859 9540
rect 4801 9531 4859 9537
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9568 6239 9571
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6227 9540 6561 9568
rect 6227 9537 6239 9540
rect 6181 9531 6239 9537
rect 6549 9537 6561 9540
rect 6595 9568 6607 9571
rect 6638 9568 6644 9580
rect 6595 9540 6644 9568
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 6638 9528 6644 9540
rect 6696 9568 6702 9580
rect 7392 9577 7420 9608
rect 7650 9596 7656 9608
rect 7708 9596 7714 9648
rect 18506 9636 18512 9648
rect 18467 9608 18512 9636
rect 18506 9596 18512 9608
rect 18564 9596 18570 9648
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 6696 9540 7205 9568
rect 6696 9528 6702 9540
rect 7193 9537 7205 9540
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 8294 9568 8300 9580
rect 7515 9540 8300 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 8294 9528 8300 9540
rect 8352 9528 8358 9580
rect 4617 9503 4675 9509
rect 4617 9469 4629 9503
rect 4663 9469 4675 9503
rect 4890 9500 4896 9512
rect 4851 9472 4896 9500
rect 4617 9463 4675 9469
rect 1578 9392 1584 9444
rect 1636 9432 1642 9444
rect 1765 9435 1823 9441
rect 1765 9432 1777 9435
rect 1636 9404 1777 9432
rect 1636 9392 1642 9404
rect 1765 9401 1777 9404
rect 1811 9401 1823 9435
rect 1765 9395 1823 9401
rect 1854 9364 1860 9376
rect 1815 9336 1860 9364
rect 1854 9324 1860 9336
rect 1912 9324 1918 9376
rect 2225 9367 2283 9373
rect 2225 9333 2237 9367
rect 2271 9364 2283 9367
rect 2314 9364 2320 9376
rect 2271 9336 2320 9364
rect 2271 9333 2283 9336
rect 2225 9327 2283 9333
rect 2314 9324 2320 9336
rect 2372 9324 2378 9376
rect 4338 9324 4344 9376
rect 4396 9364 4402 9376
rect 4433 9367 4491 9373
rect 4433 9364 4445 9367
rect 4396 9336 4445 9364
rect 4396 9324 4402 9336
rect 4433 9333 4445 9336
rect 4479 9333 4491 9367
rect 4632 9364 4660 9463
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 6089 9503 6147 9509
rect 6089 9500 6101 9503
rect 5092 9472 6101 9500
rect 4982 9392 4988 9444
rect 5040 9432 5046 9444
rect 5092 9441 5120 9472
rect 6089 9469 6101 9472
rect 6135 9469 6147 9503
rect 6089 9463 6147 9469
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 6871 9472 6929 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 6917 9469 6929 9472
rect 6963 9469 6975 9503
rect 6917 9463 6975 9469
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9469 7343 9503
rect 7285 9463 7343 9469
rect 5077 9435 5135 9441
rect 5077 9432 5089 9435
rect 5040 9404 5089 9432
rect 5040 9392 5046 9404
rect 5077 9401 5089 9404
rect 5123 9401 5135 9435
rect 5077 9395 5135 9401
rect 5261 9435 5319 9441
rect 5261 9401 5273 9435
rect 5307 9432 5319 9435
rect 5350 9432 5356 9444
rect 5307 9404 5356 9432
rect 5307 9401 5319 9404
rect 5261 9395 5319 9401
rect 5350 9392 5356 9404
rect 5408 9392 5414 9444
rect 5445 9435 5503 9441
rect 5445 9401 5457 9435
rect 5491 9432 5503 9435
rect 6730 9432 6736 9444
rect 5491 9404 6736 9432
rect 5491 9401 5503 9404
rect 5445 9395 5503 9401
rect 5460 9364 5488 9395
rect 6730 9392 6736 9404
rect 6788 9432 6794 9444
rect 7300 9432 7328 9463
rect 14550 9460 14556 9512
rect 14608 9500 14614 9512
rect 15657 9503 15715 9509
rect 15657 9500 15669 9503
rect 14608 9472 15669 9500
rect 14608 9460 14614 9472
rect 15657 9469 15669 9472
rect 15703 9469 15715 9503
rect 15657 9463 15715 9469
rect 15746 9460 15752 9512
rect 15804 9500 15810 9512
rect 18690 9500 18696 9512
rect 15804 9472 15849 9500
rect 18651 9472 18696 9500
rect 15804 9460 15810 9472
rect 18690 9460 18696 9472
rect 18748 9460 18754 9512
rect 6788 9404 7328 9432
rect 6788 9392 6794 9404
rect 15470 9392 15476 9444
rect 15528 9432 15534 9444
rect 15841 9435 15899 9441
rect 15841 9432 15853 9435
rect 15528 9404 15853 9432
rect 15528 9392 15534 9404
rect 15841 9401 15853 9404
rect 15887 9401 15899 9435
rect 15841 9395 15899 9401
rect 4632 9336 5488 9364
rect 6549 9367 6607 9373
rect 4433 9327 4491 9333
rect 6549 9333 6561 9367
rect 6595 9364 6607 9367
rect 6822 9364 6828 9376
rect 6595 9336 6828 9364
rect 6595 9333 6607 9336
rect 6549 9327 6607 9333
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 1104 9274 19044 9296
rect 1104 9222 6962 9274
rect 7014 9222 7026 9274
rect 7078 9222 7090 9274
rect 7142 9222 7154 9274
rect 7206 9222 12942 9274
rect 12994 9222 13006 9274
rect 13058 9222 13070 9274
rect 13122 9222 13134 9274
rect 13186 9222 19044 9274
rect 1104 9200 19044 9222
rect 1854 9120 1860 9172
rect 1912 9160 1918 9172
rect 3881 9163 3939 9169
rect 3881 9160 3893 9163
rect 1912 9132 3893 9160
rect 1912 9120 1918 9132
rect 3881 9129 3893 9132
rect 3927 9129 3939 9163
rect 4890 9160 4896 9172
rect 3881 9123 3939 9129
rect 4080 9132 4896 9160
rect 2498 9052 2504 9104
rect 2556 9092 2562 9104
rect 2593 9095 2651 9101
rect 2593 9092 2605 9095
rect 2556 9064 2605 9092
rect 2556 9052 2562 9064
rect 2593 9061 2605 9064
rect 2639 9061 2651 9095
rect 2593 9055 2651 9061
rect 1578 9024 1584 9036
rect 1539 8996 1584 9024
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 4080 9033 4108 9132
rect 4890 9120 4896 9132
rect 4948 9160 4954 9172
rect 5350 9160 5356 9172
rect 4948 9132 5356 9160
rect 4948 9120 4954 9132
rect 5350 9120 5356 9132
rect 5408 9160 5414 9172
rect 9122 9160 9128 9172
rect 5408 9132 9128 9160
rect 5408 9120 5414 9132
rect 9122 9120 9128 9132
rect 9180 9160 9186 9172
rect 11241 9163 11299 9169
rect 9180 9132 9444 9160
rect 9180 9120 9186 9132
rect 4522 9052 4528 9104
rect 4580 9092 4586 9104
rect 4706 9092 4712 9104
rect 4580 9064 4712 9092
rect 4580 9052 4586 9064
rect 4706 9052 4712 9064
rect 4764 9052 4770 9104
rect 9416 9101 9444 9132
rect 11241 9129 11253 9163
rect 11287 9160 11299 9163
rect 11606 9160 11612 9172
rect 11287 9132 11612 9160
rect 11287 9129 11299 9132
rect 11241 9123 11299 9129
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 13173 9163 13231 9169
rect 13173 9129 13185 9163
rect 13219 9129 13231 9163
rect 14550 9160 14556 9172
rect 14511 9132 14556 9160
rect 13173 9123 13231 9129
rect 9674 9101 9680 9104
rect 7193 9095 7251 9101
rect 7193 9092 7205 9095
rect 5368 9064 7205 9092
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 8993 4123 9027
rect 4065 8987 4123 8993
rect 4341 9027 4399 9033
rect 4341 8993 4353 9027
rect 4387 9024 4399 9027
rect 5258 9024 5264 9036
rect 4387 8996 5264 9024
rect 4387 8993 4399 8996
rect 4341 8987 4399 8993
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 5368 9033 5396 9064
rect 7193 9061 7205 9064
rect 7239 9092 7251 9095
rect 9401 9095 9459 9101
rect 7239 9064 9260 9092
rect 7239 9061 7251 9064
rect 7193 9055 7251 9061
rect 5353 9027 5411 9033
rect 5353 8993 5365 9027
rect 5399 8993 5411 9027
rect 5353 8987 5411 8993
rect 6270 8984 6276 9036
rect 6328 9024 6334 9036
rect 6641 9027 6699 9033
rect 6641 9024 6653 9027
rect 6328 8996 6653 9024
rect 6328 8984 6334 8996
rect 6641 8993 6653 8996
rect 6687 8993 6699 9027
rect 6641 8987 6699 8993
rect 7285 9027 7343 9033
rect 7285 8993 7297 9027
rect 7331 9024 7343 9027
rect 7650 9024 7656 9036
rect 7331 8996 7656 9024
rect 7331 8993 7343 8996
rect 7285 8987 7343 8993
rect 4982 8916 4988 8968
rect 5040 8956 5046 8968
rect 5077 8959 5135 8965
rect 5077 8956 5089 8959
rect 5040 8928 5089 8956
rect 5040 8916 5046 8928
rect 5077 8925 5089 8928
rect 5123 8925 5135 8959
rect 5077 8919 5135 8925
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 6917 8959 6975 8965
rect 5215 8928 5304 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5276 8900 5304 8928
rect 6917 8925 6929 8959
rect 6963 8956 6975 8959
rect 7300 8956 7328 8987
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 8202 8984 8208 9036
rect 8260 9024 8266 9036
rect 8481 9027 8539 9033
rect 8481 9024 8493 9027
rect 8260 8996 8493 9024
rect 8260 8984 8266 8996
rect 8481 8993 8493 8996
rect 8527 8993 8539 9027
rect 8481 8987 8539 8993
rect 8570 8984 8576 9036
rect 8628 9024 8634 9036
rect 9125 9027 9183 9033
rect 9125 9024 9137 9027
rect 8628 8996 9137 9024
rect 8628 8984 8634 8996
rect 9125 8993 9137 8996
rect 9171 8993 9183 9027
rect 9232 9024 9260 9064
rect 9401 9061 9413 9095
rect 9447 9061 9459 9095
rect 9401 9055 9459 9061
rect 9617 9095 9680 9101
rect 9617 9061 9629 9095
rect 9663 9061 9680 9095
rect 9617 9055 9680 9061
rect 9674 9052 9680 9055
rect 9732 9052 9738 9104
rect 12621 9095 12679 9101
rect 12621 9061 12633 9095
rect 12667 9092 12679 9095
rect 13188 9092 13216 9123
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 14461 9095 14519 9101
rect 14461 9092 14473 9095
rect 12667 9064 14473 9092
rect 12667 9061 12679 9064
rect 12621 9055 12679 9061
rect 14461 9061 14473 9064
rect 14507 9061 14519 9095
rect 14461 9055 14519 9061
rect 11333 9027 11391 9033
rect 11333 9024 11345 9027
rect 9232 8996 11345 9024
rect 9125 8987 9183 8993
rect 11333 8993 11345 8996
rect 11379 8993 11391 9027
rect 11333 8987 11391 8993
rect 12342 8984 12348 9036
rect 12400 9024 12406 9036
rect 12529 9027 12587 9033
rect 12529 9024 12541 9027
rect 12400 8996 12541 9024
rect 12400 8984 12406 8996
rect 12529 8993 12541 8996
rect 12575 8993 12587 9027
rect 12529 8987 12587 8993
rect 13081 9027 13139 9033
rect 13081 8993 13093 9027
rect 13127 9024 13139 9027
rect 13262 9024 13268 9036
rect 13127 8996 13268 9024
rect 13127 8993 13139 8996
rect 13081 8987 13139 8993
rect 13262 8984 13268 8996
rect 13320 9024 13326 9036
rect 13541 9027 13599 9033
rect 13541 9024 13553 9027
rect 13320 8996 13553 9024
rect 13320 8984 13326 8996
rect 13541 8993 13553 8996
rect 13587 8993 13599 9027
rect 13541 8987 13599 8993
rect 6963 8928 7328 8956
rect 8757 8959 8815 8965
rect 6963 8925 6975 8928
rect 6917 8919 6975 8925
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 8846 8956 8852 8968
rect 8803 8928 8852 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 8846 8916 8852 8928
rect 8904 8956 8910 8968
rect 9217 8959 9275 8965
rect 9217 8956 9229 8959
rect 8904 8928 9229 8956
rect 8904 8916 8910 8928
rect 9217 8925 9229 8928
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8956 11207 8959
rect 11422 8956 11428 8968
rect 11195 8928 11428 8956
rect 11195 8925 11207 8928
rect 11149 8919 11207 8925
rect 11422 8916 11428 8928
rect 11480 8956 11486 8968
rect 12158 8956 12164 8968
rect 11480 8928 12164 8956
rect 11480 8916 11486 8928
rect 12158 8916 12164 8928
rect 12216 8916 12222 8968
rect 12894 8916 12900 8968
rect 12952 8956 12958 8968
rect 13173 8959 13231 8965
rect 13173 8956 13185 8959
rect 12952 8928 13185 8956
rect 12952 8916 12958 8928
rect 13173 8925 13185 8928
rect 13219 8925 13231 8959
rect 13173 8919 13231 8925
rect 1394 8888 1400 8900
rect 1355 8860 1400 8888
rect 1394 8848 1400 8860
rect 1452 8848 1458 8900
rect 2774 8848 2780 8900
rect 2832 8888 2838 8900
rect 4249 8891 4307 8897
rect 2832 8860 2877 8888
rect 2832 8848 2838 8860
rect 4249 8857 4261 8891
rect 4295 8888 4307 8891
rect 4614 8888 4620 8900
rect 4295 8860 4620 8888
rect 4295 8857 4307 8860
rect 4249 8851 4307 8857
rect 4614 8848 4620 8860
rect 4672 8848 4678 8900
rect 5258 8848 5264 8900
rect 5316 8848 5322 8900
rect 6638 8848 6644 8900
rect 6696 8888 6702 8900
rect 6733 8891 6791 8897
rect 6733 8888 6745 8891
rect 6696 8860 6745 8888
rect 6696 8848 6702 8860
rect 6733 8857 6745 8860
rect 6779 8857 6791 8891
rect 6733 8851 6791 8857
rect 6825 8891 6883 8897
rect 6825 8857 6837 8891
rect 6871 8888 6883 8891
rect 7374 8888 7380 8900
rect 6871 8860 7380 8888
rect 6871 8857 6883 8860
rect 6825 8851 6883 8857
rect 7374 8848 7380 8860
rect 7432 8848 7438 8900
rect 8665 8891 8723 8897
rect 8665 8857 8677 8891
rect 8711 8888 8723 8891
rect 9674 8888 9680 8900
rect 8711 8860 9680 8888
rect 8711 8857 8723 8860
rect 8665 8851 8723 8857
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 4522 8780 4528 8832
rect 4580 8820 4586 8832
rect 4893 8823 4951 8829
rect 4893 8820 4905 8823
rect 4580 8792 4905 8820
rect 4580 8780 4586 8792
rect 4893 8789 4905 8792
rect 4939 8789 4951 8823
rect 8294 8820 8300 8832
rect 8255 8792 8300 8820
rect 4893 8783 4951 8789
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 8938 8780 8944 8832
rect 8996 8820 9002 8832
rect 9585 8823 9643 8829
rect 9585 8820 9597 8823
rect 8996 8792 9597 8820
rect 8996 8780 9002 8792
rect 9585 8789 9597 8792
rect 9631 8789 9643 8823
rect 9585 8783 9643 8789
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 10318 8820 10324 8832
rect 9824 8792 10324 8820
rect 9824 8780 9830 8792
rect 10318 8780 10324 8792
rect 10376 8780 10382 8832
rect 11701 8823 11759 8829
rect 11701 8789 11713 8823
rect 11747 8820 11759 8823
rect 14458 8820 14464 8832
rect 11747 8792 14464 8820
rect 11747 8789 11759 8792
rect 11701 8783 11759 8789
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 1104 8730 19044 8752
rect 1104 8678 3972 8730
rect 4024 8678 4036 8730
rect 4088 8678 4100 8730
rect 4152 8678 4164 8730
rect 4216 8678 9952 8730
rect 10004 8678 10016 8730
rect 10068 8678 10080 8730
rect 10132 8678 10144 8730
rect 10196 8678 15932 8730
rect 15984 8678 15996 8730
rect 16048 8678 16060 8730
rect 16112 8678 16124 8730
rect 16176 8678 19044 8730
rect 1104 8656 19044 8678
rect 8570 8576 8576 8628
rect 8628 8616 8634 8628
rect 8849 8619 8907 8625
rect 8849 8616 8861 8619
rect 8628 8588 8861 8616
rect 8628 8576 8634 8588
rect 8849 8585 8861 8588
rect 8895 8585 8907 8619
rect 8849 8579 8907 8585
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 9674 8616 9680 8628
rect 9355 8588 9680 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 12894 8616 12900 8628
rect 12855 8588 12900 8616
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 15013 8619 15071 8625
rect 15013 8585 15025 8619
rect 15059 8616 15071 8619
rect 15473 8619 15531 8625
rect 15473 8616 15485 8619
rect 15059 8588 15485 8616
rect 15059 8585 15071 8588
rect 15013 8579 15071 8585
rect 15473 8585 15485 8588
rect 15519 8585 15531 8619
rect 15473 8579 15531 8585
rect 2685 8551 2743 8557
rect 2685 8517 2697 8551
rect 2731 8548 2743 8551
rect 2777 8551 2835 8557
rect 2777 8548 2789 8551
rect 2731 8520 2789 8548
rect 2731 8517 2743 8520
rect 2685 8511 2743 8517
rect 2777 8517 2789 8520
rect 2823 8517 2835 8551
rect 2777 8511 2835 8517
rect 4433 8551 4491 8557
rect 4433 8517 4445 8551
rect 4479 8548 4491 8551
rect 12069 8551 12127 8557
rect 4479 8520 10916 8548
rect 4479 8517 4491 8520
rect 4433 8511 4491 8517
rect 2314 8480 2320 8492
rect 1688 8452 2320 8480
rect 1688 8421 1716 8452
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8480 4123 8483
rect 4338 8480 4344 8492
rect 4111 8452 4344 8480
rect 4111 8449 4123 8452
rect 4065 8443 4123 8449
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 4706 8440 4712 8492
rect 4764 8480 4770 8492
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 4764 8452 5917 8480
rect 4764 8440 4770 8452
rect 5905 8449 5917 8452
rect 5951 8480 5963 8483
rect 7282 8480 7288 8492
rect 5951 8452 7288 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 7282 8440 7288 8452
rect 7340 8480 7346 8492
rect 8205 8483 8263 8489
rect 8205 8480 8217 8483
rect 7340 8452 8217 8480
rect 7340 8440 7346 8452
rect 8205 8449 8217 8452
rect 8251 8449 8263 8483
rect 8386 8480 8392 8492
rect 8347 8452 8392 8480
rect 8205 8443 8263 8449
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8480 9275 8483
rect 9306 8480 9312 8492
rect 9263 8452 9312 8480
rect 9263 8449 9275 8452
rect 9217 8443 9275 8449
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 10888 8480 10916 8520
rect 12069 8517 12081 8551
rect 12115 8548 12127 8551
rect 12161 8551 12219 8557
rect 12161 8548 12173 8551
rect 12115 8520 12173 8548
rect 12115 8517 12127 8520
rect 12069 8511 12127 8517
rect 12161 8517 12173 8520
rect 12207 8517 12219 8551
rect 12161 8511 12219 8517
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 10888 8452 11713 8480
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8381 1731 8415
rect 1673 8375 1731 8381
rect 2225 8415 2283 8421
rect 2225 8381 2237 8415
rect 2271 8412 2283 8415
rect 2774 8412 2780 8424
rect 2271 8384 2780 8412
rect 2271 8381 2283 8384
rect 2225 8375 2283 8381
rect 2774 8372 2780 8384
rect 2832 8412 2838 8424
rect 2961 8415 3019 8421
rect 2961 8412 2973 8415
rect 2832 8384 2973 8412
rect 2832 8372 2838 8384
rect 2961 8381 2973 8384
rect 3007 8412 3019 8415
rect 3142 8412 3148 8424
rect 3007 8384 3148 8412
rect 3007 8381 3019 8384
rect 2961 8375 3019 8381
rect 3142 8372 3148 8384
rect 3200 8372 3206 8424
rect 3418 8372 3424 8424
rect 3476 8412 3482 8424
rect 5813 8415 5871 8421
rect 3476 8384 4016 8412
rect 3476 8372 3482 8384
rect 2133 8347 2191 8353
rect 2133 8313 2145 8347
rect 2179 8344 2191 8347
rect 2498 8344 2504 8356
rect 2179 8316 2504 8344
rect 2179 8313 2191 8316
rect 2133 8307 2191 8313
rect 2498 8304 2504 8316
rect 2556 8344 2562 8356
rect 3988 8353 4016 8384
rect 5813 8381 5825 8415
rect 5859 8412 5871 8415
rect 5994 8412 6000 8424
rect 5859 8384 6000 8412
rect 5859 8381 5871 8384
rect 5813 8375 5871 8381
rect 5994 8372 6000 8384
rect 6052 8372 6058 8424
rect 10888 8421 10916 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 15105 8483 15163 8489
rect 15105 8480 15117 8483
rect 11701 8443 11759 8449
rect 14476 8452 15117 8480
rect 14476 8424 14504 8452
rect 15105 8449 15117 8452
rect 15151 8449 15163 8483
rect 15488 8480 15516 8579
rect 18049 8551 18107 8557
rect 18049 8517 18061 8551
rect 18095 8548 18107 8551
rect 18141 8551 18199 8557
rect 18141 8548 18153 8551
rect 18095 8520 18153 8548
rect 18095 8517 18107 8520
rect 18049 8511 18107 8517
rect 18141 8517 18153 8520
rect 18187 8517 18199 8551
rect 18141 8511 18199 8517
rect 15488 8452 16528 8480
rect 15105 8443 15163 8449
rect 9493 8415 9551 8421
rect 9493 8381 9505 8415
rect 9539 8381 9551 8415
rect 9493 8375 9551 8381
rect 10873 8415 10931 8421
rect 10873 8381 10885 8415
rect 10919 8381 10931 8415
rect 10873 8375 10931 8381
rect 3881 8347 3939 8353
rect 2556 8316 2728 8344
rect 2556 8304 2562 8316
rect 2700 8285 2728 8316
rect 3881 8313 3893 8347
rect 3927 8313 3939 8347
rect 3881 8307 3939 8313
rect 3973 8347 4031 8353
rect 3973 8313 3985 8347
rect 4019 8313 4031 8347
rect 3973 8307 4031 8313
rect 5721 8347 5779 8353
rect 5721 8313 5733 8347
rect 5767 8344 5779 8347
rect 8202 8344 8208 8356
rect 5767 8316 8208 8344
rect 5767 8313 5779 8316
rect 5721 8307 5779 8313
rect 2685 8279 2743 8285
rect 2685 8245 2697 8279
rect 2731 8245 2743 8279
rect 3896 8276 3924 8307
rect 8202 8304 8208 8316
rect 8260 8344 8266 8356
rect 9508 8344 9536 8375
rect 11054 8372 11060 8424
rect 11112 8412 11118 8424
rect 11425 8415 11483 8421
rect 11425 8412 11437 8415
rect 11112 8384 11437 8412
rect 11112 8372 11118 8384
rect 11425 8381 11437 8384
rect 11471 8412 11483 8415
rect 12342 8412 12348 8424
rect 11471 8384 12348 8412
rect 11471 8381 11483 8384
rect 11425 8375 11483 8381
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 14458 8412 14464 8424
rect 14419 8384 14464 8412
rect 14458 8372 14464 8384
rect 14516 8372 14522 8424
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 15013 8415 15071 8421
rect 15013 8412 15025 8415
rect 14608 8384 15025 8412
rect 14608 8372 14614 8384
rect 15013 8381 15025 8384
rect 15059 8381 15071 8415
rect 15470 8412 15476 8424
rect 15431 8384 15476 8412
rect 15013 8375 15071 8381
rect 15470 8372 15476 8384
rect 15528 8372 15534 8424
rect 16500 8421 16528 8452
rect 17052 8452 18368 8480
rect 16485 8415 16543 8421
rect 16485 8381 16497 8415
rect 16531 8381 16543 8415
rect 16666 8412 16672 8424
rect 16579 8384 16672 8412
rect 16485 8375 16543 8381
rect 16666 8372 16672 8384
rect 16724 8412 16730 8424
rect 17052 8421 17080 8452
rect 17037 8415 17095 8421
rect 17037 8412 17049 8415
rect 16724 8384 17049 8412
rect 16724 8372 16730 8384
rect 17037 8381 17049 8384
rect 17083 8381 17095 8415
rect 17037 8375 17095 8381
rect 17494 8372 17500 8424
rect 17552 8412 17558 8424
rect 18340 8421 18368 8452
rect 17589 8415 17647 8421
rect 17589 8412 17601 8415
rect 17552 8384 17601 8412
rect 17552 8372 17558 8384
rect 17589 8381 17601 8384
rect 17635 8412 17647 8415
rect 17681 8415 17739 8421
rect 17681 8412 17693 8415
rect 17635 8384 17693 8412
rect 17635 8381 17647 8384
rect 17589 8375 17647 8381
rect 17681 8381 17693 8384
rect 17727 8381 17739 8415
rect 17681 8375 17739 8381
rect 18325 8415 18383 8421
rect 18325 8381 18337 8415
rect 18371 8381 18383 8415
rect 18325 8375 18383 8381
rect 8260 8316 9536 8344
rect 9677 8347 9735 8353
rect 8260 8304 8266 8316
rect 9677 8313 9689 8347
rect 9723 8344 9735 8347
rect 11238 8344 11244 8356
rect 9723 8316 11244 8344
rect 9723 8313 9735 8316
rect 9677 8307 9735 8313
rect 11238 8304 11244 8316
rect 11296 8304 11302 8356
rect 11333 8347 11391 8353
rect 11333 8313 11345 8347
rect 11379 8344 11391 8347
rect 12805 8347 12863 8353
rect 12805 8344 12817 8347
rect 11379 8316 12817 8344
rect 11379 8313 11391 8316
rect 11333 8307 11391 8313
rect 4706 8276 4712 8288
rect 3896 8248 4712 8276
rect 2685 8239 2743 8245
rect 4706 8236 4712 8248
rect 4764 8236 4770 8288
rect 5350 8276 5356 8288
rect 5311 8248 5356 8276
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 8478 8236 8484 8288
rect 8536 8276 8542 8288
rect 12084 8285 12112 8316
rect 12805 8313 12817 8316
rect 12851 8313 12863 8347
rect 17126 8344 17132 8356
rect 17087 8316 17132 8344
rect 12805 8307 12863 8313
rect 17126 8304 17132 8316
rect 17184 8344 17190 8356
rect 17184 8316 18092 8344
rect 17184 8304 17190 8316
rect 18064 8285 18092 8316
rect 12069 8279 12127 8285
rect 8536 8248 8581 8276
rect 8536 8236 8542 8248
rect 12069 8245 12081 8279
rect 12115 8245 12127 8279
rect 12069 8239 12127 8245
rect 18049 8279 18107 8285
rect 18049 8245 18061 8279
rect 18095 8245 18107 8279
rect 18049 8239 18107 8245
rect 1104 8186 19044 8208
rect 1104 8134 6962 8186
rect 7014 8134 7026 8186
rect 7078 8134 7090 8186
rect 7142 8134 7154 8186
rect 7206 8134 12942 8186
rect 12994 8134 13006 8186
rect 13058 8134 13070 8186
rect 13122 8134 13134 8186
rect 13186 8134 19044 8186
rect 1104 8112 19044 8134
rect 2498 8072 2504 8084
rect 2459 8044 2504 8072
rect 2498 8032 2504 8044
rect 2556 8032 2562 8084
rect 2682 8032 2688 8084
rect 2740 8072 2746 8084
rect 4341 8075 4399 8081
rect 4341 8072 4353 8075
rect 2740 8044 4353 8072
rect 2740 8032 2746 8044
rect 4341 8041 4353 8044
rect 4387 8041 4399 8075
rect 8478 8072 8484 8084
rect 8439 8044 8484 8072
rect 4341 8035 4399 8041
rect 8478 8032 8484 8044
rect 8536 8032 8542 8084
rect 8662 8032 8668 8084
rect 8720 8072 8726 8084
rect 9122 8072 9128 8084
rect 8720 8044 9128 8072
rect 8720 8032 8726 8044
rect 9122 8032 9128 8044
rect 9180 8032 9186 8084
rect 17126 8032 17132 8084
rect 17184 8072 17190 8084
rect 17589 8075 17647 8081
rect 17589 8072 17601 8075
rect 17184 8044 17601 8072
rect 17184 8032 17190 8044
rect 17589 8041 17601 8044
rect 17635 8041 17647 8075
rect 17589 8035 17647 8041
rect 4522 8004 4528 8016
rect 4483 7976 4528 8004
rect 4522 7964 4528 7976
rect 4580 7964 4586 8016
rect 7466 8004 7472 8016
rect 7427 7976 7472 8004
rect 7466 7964 7472 7976
rect 7524 7964 7530 8016
rect 10873 8007 10931 8013
rect 10873 8004 10885 8007
rect 7852 7976 10885 8004
rect 7852 7948 7880 7976
rect 10873 7973 10885 7976
rect 10919 7973 10931 8007
rect 11054 8004 11060 8016
rect 11015 7976 11060 8004
rect 10873 7967 10931 7973
rect 11054 7964 11060 7976
rect 11112 7964 11118 8016
rect 7377 7939 7435 7945
rect 7377 7905 7389 7939
rect 7423 7936 7435 7939
rect 7561 7939 7619 7945
rect 7561 7936 7573 7939
rect 7423 7908 7573 7936
rect 7423 7905 7435 7908
rect 7377 7899 7435 7905
rect 7561 7905 7573 7908
rect 7607 7905 7619 7939
rect 7834 7936 7840 7948
rect 7747 7908 7840 7936
rect 7561 7899 7619 7905
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 8662 7936 8668 7948
rect 8623 7908 8668 7936
rect 8662 7896 8668 7908
rect 8720 7896 8726 7948
rect 8846 7936 8852 7948
rect 8807 7908 8852 7936
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 8938 7896 8944 7948
rect 8996 7936 9002 7948
rect 9122 7936 9128 7948
rect 8996 7908 9041 7936
rect 9083 7908 9128 7936
rect 8996 7896 9002 7908
rect 9122 7896 9128 7908
rect 9180 7896 9186 7948
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4706 7868 4712 7880
rect 4295 7840 4712 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 8956 7868 8984 7896
rect 9217 7871 9275 7877
rect 9217 7868 9229 7871
rect 8956 7840 9229 7868
rect 9217 7837 9229 7840
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 4801 7803 4859 7809
rect 4801 7769 4813 7803
rect 4847 7800 4859 7803
rect 9766 7800 9772 7812
rect 4847 7772 9772 7800
rect 4847 7769 4859 7772
rect 4801 7763 4859 7769
rect 9766 7760 9772 7772
rect 9824 7760 9830 7812
rect 2498 7692 2504 7744
rect 2556 7732 2562 7744
rect 2593 7735 2651 7741
rect 2593 7732 2605 7735
rect 2556 7704 2605 7732
rect 2556 7692 2562 7704
rect 2593 7701 2605 7704
rect 2639 7701 2651 7735
rect 2593 7695 2651 7701
rect 8846 7692 8852 7744
rect 8904 7732 8910 7744
rect 9125 7735 9183 7741
rect 9125 7732 9137 7735
rect 8904 7704 9137 7732
rect 8904 7692 8910 7704
rect 9125 7701 9137 7704
rect 9171 7701 9183 7735
rect 9125 7695 9183 7701
rect 9493 7735 9551 7741
rect 9493 7701 9505 7735
rect 9539 7732 9551 7735
rect 9582 7732 9588 7744
rect 9539 7704 9588 7732
rect 9539 7701 9551 7704
rect 9493 7695 9551 7701
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 16758 7692 16764 7744
rect 16816 7732 16822 7744
rect 17497 7735 17555 7741
rect 17497 7732 17509 7735
rect 16816 7704 17509 7732
rect 16816 7692 16822 7704
rect 17497 7701 17509 7704
rect 17543 7701 17555 7735
rect 17497 7695 17555 7701
rect 1104 7642 19044 7664
rect 1104 7590 3972 7642
rect 4024 7590 4036 7642
rect 4088 7590 4100 7642
rect 4152 7590 4164 7642
rect 4216 7590 9952 7642
rect 10004 7590 10016 7642
rect 10068 7590 10080 7642
rect 10132 7590 10144 7642
rect 10196 7590 15932 7642
rect 15984 7590 15996 7642
rect 16048 7590 16060 7642
rect 16112 7590 16124 7642
rect 16176 7590 19044 7642
rect 1104 7568 19044 7590
rect 13354 7528 13360 7540
rect 13267 7500 13360 7528
rect 13354 7488 13360 7500
rect 13412 7528 13418 7540
rect 13817 7531 13875 7537
rect 13817 7528 13829 7531
rect 13412 7500 13829 7528
rect 13412 7488 13418 7500
rect 13817 7497 13829 7500
rect 13863 7497 13875 7531
rect 13817 7491 13875 7497
rect 2498 7460 2504 7472
rect 2459 7432 2504 7460
rect 2498 7420 2504 7432
rect 2556 7420 2562 7472
rect 16758 7460 16764 7472
rect 16719 7432 16764 7460
rect 16758 7420 16764 7432
rect 16816 7420 16822 7472
rect 13449 7395 13507 7401
rect 13449 7392 13461 7395
rect 12820 7364 13461 7392
rect 2133 7327 2191 7333
rect 2133 7293 2145 7327
rect 2179 7324 2191 7327
rect 2498 7324 2504 7336
rect 2179 7296 2504 7324
rect 2179 7293 2191 7296
rect 2133 7287 2191 7293
rect 2498 7284 2504 7296
rect 2556 7284 2562 7336
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7293 4031 7327
rect 3973 7287 4031 7293
rect 4249 7327 4307 7333
rect 4249 7293 4261 7327
rect 4295 7324 4307 7327
rect 4614 7324 4620 7336
rect 4295 7296 4620 7324
rect 4295 7293 4307 7296
rect 4249 7287 4307 7293
rect 3988 7256 4016 7287
rect 4614 7284 4620 7296
rect 4672 7284 4678 7336
rect 6638 7324 6644 7336
rect 6599 7296 6644 7324
rect 6638 7284 6644 7296
rect 6696 7284 6702 7336
rect 7282 7324 7288 7336
rect 7243 7296 7288 7324
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 8938 7284 8944 7336
rect 8996 7324 9002 7336
rect 10965 7327 11023 7333
rect 10965 7324 10977 7327
rect 8996 7296 10977 7324
rect 8996 7284 9002 7296
rect 10965 7293 10977 7296
rect 11011 7293 11023 7327
rect 10965 7287 11023 7293
rect 12618 7284 12624 7336
rect 12676 7324 12682 7336
rect 12820 7333 12848 7364
rect 13449 7361 13461 7364
rect 13495 7361 13507 7395
rect 16666 7392 16672 7404
rect 13449 7355 13507 7361
rect 16316 7364 16672 7392
rect 12805 7327 12863 7333
rect 12805 7324 12817 7327
rect 12676 7296 12817 7324
rect 12676 7284 12682 7296
rect 12805 7293 12817 7296
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 13357 7327 13415 7333
rect 13357 7293 13369 7327
rect 13403 7293 13415 7327
rect 13814 7324 13820 7336
rect 13775 7296 13820 7324
rect 13357 7287 13415 7293
rect 6822 7256 6828 7268
rect 3988 7228 6828 7256
rect 6822 7216 6828 7228
rect 6880 7216 6886 7268
rect 9122 7216 9128 7268
rect 9180 7256 9186 7268
rect 11149 7259 11207 7265
rect 11149 7256 11161 7259
rect 9180 7228 11161 7256
rect 9180 7216 9186 7228
rect 11149 7225 11161 7228
rect 11195 7225 11207 7259
rect 13372 7256 13400 7287
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 15746 7324 15752 7336
rect 15707 7296 15752 7324
rect 15746 7284 15752 7296
rect 15804 7284 15810 7336
rect 16316 7333 16344 7364
rect 16666 7352 16672 7364
rect 16724 7352 16730 7404
rect 16295 7327 16353 7333
rect 16295 7293 16307 7327
rect 16341 7293 16353 7327
rect 16295 7287 16353 7293
rect 16390 7284 16396 7336
rect 16448 7324 16454 7336
rect 16448 7296 16493 7324
rect 16448 7284 16454 7296
rect 13630 7256 13636 7268
rect 13372 7228 13636 7256
rect 11149 7219 11207 7225
rect 13630 7216 13636 7228
rect 13688 7216 13694 7268
rect 16209 7259 16267 7265
rect 16209 7225 16221 7259
rect 16255 7256 16267 7259
rect 16255 7228 16574 7256
rect 16255 7225 16267 7228
rect 16209 7219 16267 7225
rect 16546 7200 16574 7228
rect 2501 7191 2559 7197
rect 2501 7157 2513 7191
rect 2547 7188 2559 7191
rect 3326 7188 3332 7200
rect 2547 7160 3332 7188
rect 2547 7157 2559 7160
rect 2501 7151 2559 7157
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 3786 7188 3792 7200
rect 3747 7160 3792 7188
rect 3786 7148 3792 7160
rect 3844 7148 3850 7200
rect 4157 7191 4215 7197
rect 4157 7157 4169 7191
rect 4203 7188 4215 7191
rect 5258 7188 5264 7200
rect 4203 7160 5264 7188
rect 4203 7157 4215 7160
rect 4157 7151 4215 7157
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 7742 7188 7748 7200
rect 7703 7160 7748 7188
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 11333 7191 11391 7197
rect 11333 7157 11345 7191
rect 11379 7188 11391 7191
rect 12066 7188 12072 7200
rect 11379 7160 12072 7188
rect 11379 7157 11391 7160
rect 11333 7151 11391 7157
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 15746 7148 15752 7200
rect 15804 7188 15810 7200
rect 16390 7188 16396 7200
rect 15804 7160 16396 7188
rect 15804 7148 15810 7160
rect 16390 7148 16396 7160
rect 16448 7148 16454 7200
rect 16482 7148 16488 7200
rect 16540 7188 16574 7200
rect 16761 7191 16819 7197
rect 16761 7188 16773 7191
rect 16540 7160 16773 7188
rect 16540 7148 16546 7160
rect 16761 7157 16773 7160
rect 16807 7157 16819 7191
rect 16761 7151 16819 7157
rect 1104 7098 19044 7120
rect 1104 7046 6962 7098
rect 7014 7046 7026 7098
rect 7078 7046 7090 7098
rect 7142 7046 7154 7098
rect 7206 7046 12942 7098
rect 12994 7046 13006 7098
rect 13058 7046 13070 7098
rect 13122 7046 13134 7098
rect 13186 7046 19044 7098
rect 1104 7024 19044 7046
rect 2133 6987 2191 6993
rect 2133 6953 2145 6987
rect 2179 6984 2191 6987
rect 3786 6984 3792 6996
rect 2179 6956 3792 6984
rect 2179 6953 2191 6956
rect 2133 6947 2191 6953
rect 3786 6944 3792 6956
rect 3844 6944 3850 6996
rect 8757 6987 8815 6993
rect 8757 6953 8769 6987
rect 8803 6953 8815 6987
rect 12066 6984 12072 6996
rect 12027 6956 12072 6984
rect 8757 6947 8815 6953
rect 4798 6916 4804 6928
rect 4759 6888 4804 6916
rect 4798 6876 4804 6888
rect 4856 6876 4862 6928
rect 7285 6919 7343 6925
rect 7285 6885 7297 6919
rect 7331 6916 7343 6919
rect 7834 6916 7840 6928
rect 7331 6888 7840 6916
rect 7331 6885 7343 6888
rect 7285 6879 7343 6885
rect 7834 6876 7840 6888
rect 7892 6876 7898 6928
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 1964 6820 2176 6848
rect 1964 6789 1992 6820
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6749 2099 6783
rect 2041 6743 2099 6749
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 2056 6712 2084 6743
rect 1627 6684 2084 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 2148 6644 2176 6820
rect 2498 6808 2504 6860
rect 2556 6848 2562 6860
rect 2593 6851 2651 6857
rect 2593 6848 2605 6851
rect 2556 6820 2605 6848
rect 2556 6808 2562 6820
rect 2593 6817 2605 6820
rect 2639 6817 2651 6851
rect 3142 6848 3148 6860
rect 3103 6820 3148 6848
rect 2593 6811 2651 6817
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 4706 6848 4712 6860
rect 4667 6820 4712 6848
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 4982 6848 4988 6860
rect 4943 6820 4988 6848
rect 4982 6808 4988 6820
rect 5040 6808 5046 6860
rect 5718 6848 5724 6860
rect 5679 6820 5724 6848
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 5902 6848 5908 6860
rect 5863 6820 5908 6848
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 6273 6851 6331 6857
rect 6273 6817 6285 6851
rect 6319 6848 6331 6851
rect 6638 6848 6644 6860
rect 6319 6820 6644 6848
rect 6319 6817 6331 6820
rect 6273 6811 6331 6817
rect 6638 6808 6644 6820
rect 6696 6808 6702 6860
rect 7561 6851 7619 6857
rect 7561 6817 7573 6851
rect 7607 6848 7619 6851
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 7607 6820 7665 6848
rect 7607 6817 7619 6820
rect 7561 6811 7619 6817
rect 7653 6817 7665 6820
rect 7699 6817 7711 6851
rect 7653 6811 7711 6817
rect 8389 6851 8447 6857
rect 8389 6817 8401 6851
rect 8435 6848 8447 6851
rect 8570 6848 8576 6860
rect 8435 6820 8576 6848
rect 8435 6817 8447 6820
rect 8389 6811 8447 6817
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 8772 6848 8800 6947
rect 12066 6944 12072 6956
rect 12124 6944 12130 6996
rect 13354 6984 13360 6996
rect 13315 6956 13360 6984
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 13814 6984 13820 6996
rect 13775 6956 13820 6984
rect 13814 6944 13820 6956
rect 13872 6944 13878 6996
rect 16482 6916 16488 6928
rect 14568 6888 14964 6916
rect 16443 6888 16488 6916
rect 9214 6848 9220 6860
rect 8772 6820 9220 6848
rect 9214 6808 9220 6820
rect 9272 6808 9278 6860
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 9953 6851 10011 6857
rect 9953 6848 9965 6851
rect 9824 6820 9965 6848
rect 9824 6808 9830 6820
rect 9953 6817 9965 6820
rect 9999 6848 10011 6851
rect 10502 6848 10508 6860
rect 9999 6820 10508 6848
rect 9999 6817 10011 6820
rect 9953 6811 10011 6817
rect 10502 6808 10508 6820
rect 10560 6808 10566 6860
rect 10686 6848 10692 6860
rect 10647 6820 10692 6848
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 10873 6851 10931 6857
rect 10873 6817 10885 6851
rect 10919 6817 10931 6851
rect 10873 6811 10931 6817
rect 2516 6721 2544 6808
rect 4724 6780 4752 6808
rect 2746 6752 4752 6780
rect 2501 6715 2559 6721
rect 2501 6681 2513 6715
rect 2547 6681 2559 6715
rect 2501 6675 2559 6681
rect 2746 6644 2774 6752
rect 10594 6740 10600 6792
rect 10652 6780 10658 6792
rect 10888 6780 10916 6811
rect 12618 6808 12624 6860
rect 12676 6848 12682 6860
rect 13630 6848 13636 6860
rect 12676 6820 13636 6848
rect 12676 6808 12682 6820
rect 13630 6808 13636 6820
rect 13688 6848 13694 6860
rect 14568 6848 14596 6888
rect 14734 6848 14740 6860
rect 13688 6820 14596 6848
rect 14695 6820 14740 6848
rect 13688 6808 13694 6820
rect 14734 6808 14740 6820
rect 14792 6808 14798 6860
rect 14936 6848 14964 6888
rect 16482 6876 16488 6888
rect 16540 6876 16546 6928
rect 16301 6851 16359 6857
rect 16301 6848 16313 6851
rect 14936 6820 16313 6848
rect 16301 6817 16313 6820
rect 16347 6817 16359 6851
rect 18690 6848 18696 6860
rect 18651 6820 18696 6848
rect 16301 6811 16359 6817
rect 18690 6808 18696 6820
rect 18748 6808 18754 6860
rect 10652 6752 10916 6780
rect 11885 6783 11943 6789
rect 10652 6740 10658 6752
rect 11885 6749 11897 6783
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6780 12035 6783
rect 12023 6752 12434 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 5261 6715 5319 6721
rect 5261 6681 5273 6715
rect 5307 6712 5319 6715
rect 8662 6712 8668 6724
rect 5307 6684 8668 6712
rect 5307 6681 5319 6684
rect 5261 6675 5319 6681
rect 8662 6672 8668 6684
rect 8720 6672 8726 6724
rect 8757 6715 8815 6721
rect 8757 6681 8769 6715
rect 8803 6712 8815 6715
rect 9766 6712 9772 6724
rect 8803 6684 9772 6712
rect 8803 6681 8815 6684
rect 8757 6675 8815 6681
rect 9766 6672 9772 6684
rect 9824 6672 9830 6724
rect 11900 6712 11928 6743
rect 12158 6712 12164 6724
rect 11900 6684 12164 6712
rect 12158 6672 12164 6684
rect 12216 6672 12222 6724
rect 12406 6712 12434 6752
rect 13722 6740 13728 6792
rect 13780 6780 13786 6792
rect 14829 6783 14887 6789
rect 14829 6780 14841 6783
rect 13780 6752 14841 6780
rect 13780 6740 13786 6752
rect 14829 6749 14841 6752
rect 14875 6749 14887 6783
rect 15010 6780 15016 6792
rect 14971 6752 15016 6780
rect 14829 6743 14887 6749
rect 15010 6740 15016 6752
rect 15068 6740 15074 6792
rect 18509 6715 18567 6721
rect 18509 6712 18521 6715
rect 12406 6684 18521 6712
rect 18509 6681 18521 6684
rect 18555 6681 18567 6715
rect 18509 6675 18567 6681
rect 2148 6616 2774 6644
rect 3145 6647 3203 6653
rect 3145 6613 3157 6647
rect 3191 6644 3203 6647
rect 3326 6644 3332 6656
rect 3191 6616 3332 6644
rect 3191 6613 3203 6616
rect 3145 6607 3203 6613
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 12342 6604 12348 6656
rect 12400 6644 12406 6656
rect 12437 6647 12495 6653
rect 12437 6644 12449 6647
rect 12400 6616 12449 6644
rect 12400 6604 12406 6616
rect 12437 6613 12449 6616
rect 12483 6613 12495 6647
rect 12437 6607 12495 6613
rect 12710 6604 12716 6656
rect 12768 6644 12774 6656
rect 13265 6647 13323 6653
rect 13265 6644 13277 6647
rect 12768 6616 13277 6644
rect 12768 6604 12774 6616
rect 13265 6613 13277 6616
rect 13311 6613 13323 6647
rect 14366 6644 14372 6656
rect 14327 6616 14372 6644
rect 13265 6607 13323 6613
rect 14366 6604 14372 6616
rect 14424 6604 14430 6656
rect 1104 6554 19044 6576
rect 1104 6502 3972 6554
rect 4024 6502 4036 6554
rect 4088 6502 4100 6554
rect 4152 6502 4164 6554
rect 4216 6502 9952 6554
rect 10004 6502 10016 6554
rect 10068 6502 10080 6554
rect 10132 6502 10144 6554
rect 10196 6502 15932 6554
rect 15984 6502 15996 6554
rect 16048 6502 16060 6554
rect 16112 6502 16124 6554
rect 16176 6502 19044 6554
rect 1104 6480 19044 6502
rect 5902 6440 5908 6452
rect 2746 6412 5908 6440
rect 1670 6332 1676 6384
rect 1728 6372 1734 6384
rect 2746 6372 2774 6412
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 9766 6440 9772 6452
rect 9727 6412 9772 6440
rect 9766 6400 9772 6412
rect 9824 6400 9830 6452
rect 14366 6440 14372 6452
rect 12406 6412 14372 6440
rect 12406 6372 12434 6412
rect 14366 6400 14372 6412
rect 14424 6400 14430 6452
rect 15746 6440 15752 6452
rect 14476 6412 15752 6440
rect 12710 6372 12716 6384
rect 1728 6344 2774 6372
rect 4540 6344 12434 6372
rect 12671 6344 12716 6372
rect 1728 6332 1734 6344
rect 1578 6264 1584 6316
rect 1636 6304 1642 6316
rect 4540 6304 4568 6344
rect 12710 6332 12716 6344
rect 12768 6332 12774 6384
rect 1636 6276 4568 6304
rect 6917 6307 6975 6313
rect 1636 6264 1642 6276
rect 6917 6273 6929 6307
rect 6963 6304 6975 6307
rect 6963 6276 8156 6304
rect 6963 6273 6975 6276
rect 6917 6267 6975 6273
rect 6549 6239 6607 6245
rect 6549 6205 6561 6239
rect 6595 6236 6607 6239
rect 6638 6236 6644 6248
rect 6595 6208 6644 6236
rect 6595 6205 6607 6208
rect 6549 6199 6607 6205
rect 6638 6196 6644 6208
rect 6696 6236 6702 6248
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 6696 6208 7021 6236
rect 6696 6196 6702 6208
rect 7009 6205 7021 6208
rect 7055 6205 7067 6239
rect 7926 6236 7932 6248
rect 7887 6208 7932 6236
rect 7009 6199 7067 6205
rect 7926 6196 7932 6208
rect 7984 6196 7990 6248
rect 8128 6245 8156 6276
rect 8662 6264 8668 6316
rect 8720 6304 8726 6316
rect 14476 6304 14504 6412
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 15010 6372 15016 6384
rect 14660 6344 15016 6372
rect 14660 6313 14688 6344
rect 15010 6332 15016 6344
rect 15068 6332 15074 6384
rect 8720 6276 14504 6304
rect 14645 6307 14703 6313
rect 8720 6264 8726 6276
rect 14645 6273 14657 6307
rect 14691 6273 14703 6307
rect 14645 6267 14703 6273
rect 8113 6239 8171 6245
rect 8113 6205 8125 6239
rect 8159 6205 8171 6239
rect 8113 6199 8171 6205
rect 8570 6196 8576 6248
rect 8628 6236 8634 6248
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 8628 6208 9137 6236
rect 8628 6196 8634 6208
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 9125 6199 9183 6205
rect 9677 6239 9735 6245
rect 9677 6205 9689 6239
rect 9723 6236 9735 6239
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 9723 6208 9965 6236
rect 9723 6205 9735 6208
rect 9677 6199 9735 6205
rect 9953 6205 9965 6208
rect 9999 6205 10011 6239
rect 9953 6199 10011 6205
rect 10229 6239 10287 6245
rect 10229 6205 10241 6239
rect 10275 6236 10287 6239
rect 10502 6236 10508 6248
rect 10275 6208 10508 6236
rect 10275 6205 10287 6208
rect 10229 6199 10287 6205
rect 6730 6168 6736 6180
rect 6691 6140 6736 6168
rect 6730 6128 6736 6140
rect 6788 6128 6794 6180
rect 7653 6171 7711 6177
rect 7653 6137 7665 6171
rect 7699 6168 7711 6171
rect 7834 6168 7840 6180
rect 7699 6140 7840 6168
rect 7699 6137 7711 6140
rect 7653 6131 7711 6137
rect 7834 6128 7840 6140
rect 7892 6168 7898 6180
rect 8757 6171 8815 6177
rect 8757 6168 8769 6171
rect 7892 6140 8769 6168
rect 7892 6128 7898 6140
rect 8757 6137 8769 6140
rect 8803 6137 8815 6171
rect 8757 6131 8815 6137
rect 9033 6171 9091 6177
rect 9033 6137 9045 6171
rect 9079 6137 9091 6171
rect 9033 6131 9091 6137
rect 9048 6100 9076 6131
rect 9214 6128 9220 6180
rect 9272 6168 9278 6180
rect 9585 6171 9643 6177
rect 9585 6168 9597 6171
rect 9272 6140 9597 6168
rect 9272 6128 9278 6140
rect 9585 6137 9597 6140
rect 9631 6137 9643 6171
rect 9585 6131 9643 6137
rect 9692 6100 9720 6199
rect 9968 6168 9996 6199
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 10778 6196 10784 6248
rect 10836 6236 10842 6248
rect 10965 6239 11023 6245
rect 10965 6236 10977 6239
rect 10836 6208 10977 6236
rect 10836 6196 10842 6208
rect 10965 6205 10977 6208
rect 11011 6205 11023 6239
rect 12342 6236 12348 6248
rect 12303 6208 12348 6236
rect 10965 6199 11023 6205
rect 12342 6196 12348 6208
rect 12400 6196 12406 6248
rect 14826 6236 14832 6248
rect 14787 6208 14832 6236
rect 14826 6196 14832 6208
rect 14884 6196 14890 6248
rect 15013 6239 15071 6245
rect 15013 6205 15025 6239
rect 15059 6205 15071 6239
rect 15286 6236 15292 6248
rect 15247 6208 15292 6236
rect 15013 6199 15071 6205
rect 10686 6168 10692 6180
rect 9968 6140 10692 6168
rect 10686 6128 10692 6140
rect 10744 6168 10750 6180
rect 10873 6171 10931 6177
rect 10873 6168 10885 6171
rect 10744 6140 10885 6168
rect 10744 6128 10750 6140
rect 10873 6137 10885 6140
rect 10919 6137 10931 6171
rect 15028 6168 15056 6199
rect 15286 6196 15292 6208
rect 15344 6196 15350 6248
rect 15470 6168 15476 6180
rect 15028 6140 15476 6168
rect 10873 6131 10931 6137
rect 15470 6128 15476 6140
rect 15528 6128 15534 6180
rect 12710 6100 12716 6112
rect 9048 6072 9720 6100
rect 12671 6072 12716 6100
rect 12710 6060 12716 6072
rect 12768 6060 12774 6112
rect 14826 6060 14832 6112
rect 14884 6100 14890 6112
rect 16206 6100 16212 6112
rect 14884 6072 16212 6100
rect 14884 6060 14890 6072
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 1104 6010 19044 6032
rect 1104 5958 6962 6010
rect 7014 5958 7026 6010
rect 7078 5958 7090 6010
rect 7142 5958 7154 6010
rect 7206 5958 12942 6010
rect 12994 5958 13006 6010
rect 13058 5958 13070 6010
rect 13122 5958 13134 6010
rect 13186 5958 19044 6010
rect 1104 5936 19044 5958
rect 3145 5899 3203 5905
rect 3145 5865 3157 5899
rect 3191 5896 3203 5899
rect 3510 5896 3516 5908
rect 3191 5868 3516 5896
rect 3191 5865 3203 5868
rect 3145 5859 3203 5865
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 6638 5896 6644 5908
rect 4948 5868 6500 5896
rect 6599 5868 6644 5896
rect 4948 5856 4954 5868
rect 3234 5828 3240 5840
rect 3147 5800 3240 5828
rect 3234 5788 3240 5800
rect 3292 5828 3298 5840
rect 4617 5831 4675 5837
rect 4617 5828 4629 5831
rect 3292 5800 4629 5828
rect 3292 5788 3298 5800
rect 4617 5797 4629 5800
rect 4663 5828 4675 5831
rect 5353 5831 5411 5837
rect 5353 5828 5365 5831
rect 4663 5800 5365 5828
rect 4663 5797 4675 5800
rect 4617 5791 4675 5797
rect 5353 5797 5365 5800
rect 5399 5797 5411 5831
rect 6472 5828 6500 5868
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 6822 5856 6828 5908
rect 6880 5896 6886 5908
rect 7009 5899 7067 5905
rect 7009 5896 7021 5899
rect 6880 5868 7021 5896
rect 6880 5856 6886 5868
rect 7009 5865 7021 5868
rect 7055 5865 7067 5899
rect 7009 5859 7067 5865
rect 7926 5856 7932 5908
rect 7984 5896 7990 5908
rect 8297 5899 8355 5905
rect 8297 5896 8309 5899
rect 7984 5868 8309 5896
rect 7984 5856 7990 5868
rect 8297 5865 8309 5868
rect 8343 5865 8355 5899
rect 8297 5859 8355 5865
rect 8389 5899 8447 5905
rect 8389 5865 8401 5899
rect 8435 5896 8447 5899
rect 9214 5896 9220 5908
rect 8435 5868 9220 5896
rect 8435 5865 8447 5868
rect 8389 5859 8447 5865
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 10778 5896 10784 5908
rect 10739 5868 10784 5896
rect 10778 5856 10784 5868
rect 10836 5856 10842 5908
rect 14645 5899 14703 5905
rect 14645 5896 14657 5899
rect 12406 5868 14657 5896
rect 12406 5828 12434 5868
rect 14645 5865 14657 5868
rect 14691 5865 14703 5899
rect 14645 5859 14703 5865
rect 14734 5856 14740 5908
rect 14792 5896 14798 5908
rect 15105 5899 15163 5905
rect 15105 5896 15117 5899
rect 14792 5868 15117 5896
rect 14792 5856 14798 5868
rect 15105 5865 15117 5868
rect 15151 5865 15163 5899
rect 15105 5859 15163 5865
rect 15289 5899 15347 5905
rect 15289 5865 15301 5899
rect 15335 5865 15347 5899
rect 15289 5859 15347 5865
rect 6472 5800 12434 5828
rect 12529 5831 12587 5837
rect 5353 5791 5411 5797
rect 12529 5797 12541 5831
rect 12575 5828 12587 5831
rect 12710 5828 12716 5840
rect 12575 5800 12716 5828
rect 12575 5797 12587 5800
rect 12529 5791 12587 5797
rect 12710 5788 12716 5800
rect 12768 5788 12774 5840
rect 15304 5828 15332 5859
rect 16301 5831 16359 5837
rect 16301 5828 16313 5831
rect 14568 5800 15332 5828
rect 15672 5800 16313 5828
rect 3881 5763 3939 5769
rect 3881 5729 3893 5763
rect 3927 5760 3939 5763
rect 4430 5760 4436 5772
rect 3927 5732 4436 5760
rect 3927 5729 3939 5732
rect 3881 5723 3939 5729
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 4706 5720 4712 5772
rect 4764 5760 4770 5772
rect 4801 5763 4859 5769
rect 4801 5760 4813 5763
rect 4764 5732 4813 5760
rect 4764 5720 4770 5732
rect 4801 5729 4813 5732
rect 4847 5729 4859 5763
rect 4801 5723 4859 5729
rect 5445 5763 5503 5769
rect 5445 5729 5457 5763
rect 5491 5760 5503 5763
rect 5537 5763 5595 5769
rect 5537 5760 5549 5763
rect 5491 5732 5549 5760
rect 5491 5729 5503 5732
rect 5445 5723 5503 5729
rect 5537 5729 5549 5732
rect 5583 5729 5595 5763
rect 5537 5723 5595 5729
rect 5721 5763 5779 5769
rect 5721 5729 5733 5763
rect 5767 5760 5779 5763
rect 5902 5760 5908 5772
rect 5767 5732 5908 5760
rect 5767 5729 5779 5732
rect 5721 5723 5779 5729
rect 5902 5720 5908 5732
rect 5960 5720 5966 5772
rect 10502 5720 10508 5772
rect 10560 5760 10566 5772
rect 10689 5763 10747 5769
rect 10689 5760 10701 5763
rect 10560 5732 10701 5760
rect 10560 5720 10566 5732
rect 10689 5729 10701 5732
rect 10735 5729 10747 5763
rect 10689 5723 10747 5729
rect 12069 5763 12127 5769
rect 12069 5729 12081 5763
rect 12115 5760 12127 5763
rect 12342 5760 12348 5772
rect 12115 5732 12348 5760
rect 12115 5729 12127 5732
rect 12069 5723 12127 5729
rect 12342 5720 12348 5732
rect 12400 5720 12406 5772
rect 12618 5760 12624 5772
rect 12579 5732 12624 5760
rect 12618 5720 12624 5732
rect 12676 5720 12682 5772
rect 4448 5692 4476 5720
rect 4893 5695 4951 5701
rect 4893 5692 4905 5695
rect 4448 5664 4905 5692
rect 4893 5661 4905 5664
rect 4939 5661 4951 5695
rect 4893 5655 4951 5661
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5661 7159 5695
rect 7282 5692 7288 5704
rect 7243 5664 7288 5692
rect 7101 5655 7159 5661
rect 7116 5556 7144 5655
rect 7282 5652 7288 5664
rect 7340 5652 7346 5704
rect 14568 5701 14596 5800
rect 14734 5760 14740 5772
rect 14695 5732 14740 5760
rect 14734 5720 14740 5732
rect 14792 5720 14798 5772
rect 15286 5760 15292 5772
rect 15199 5732 15292 5760
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 15470 5760 15476 5772
rect 15431 5732 15476 5760
rect 15470 5720 15476 5732
rect 15528 5720 15534 5772
rect 15672 5769 15700 5800
rect 16301 5797 16313 5800
rect 16347 5828 16359 5831
rect 16390 5828 16396 5840
rect 16347 5800 16396 5828
rect 16347 5797 16359 5800
rect 16301 5791 16359 5797
rect 16390 5788 16396 5800
rect 16448 5788 16454 5840
rect 15657 5763 15715 5769
rect 15657 5729 15669 5763
rect 15703 5729 15715 5763
rect 16117 5763 16175 5769
rect 16117 5760 16129 5763
rect 15657 5723 15715 5729
rect 15948 5732 16129 5760
rect 14553 5695 14611 5701
rect 14553 5661 14565 5695
rect 14599 5661 14611 5695
rect 14553 5655 14611 5661
rect 15304 5624 15332 5720
rect 15488 5692 15516 5720
rect 15948 5692 15976 5732
rect 16117 5729 16129 5732
rect 16163 5729 16175 5763
rect 16117 5723 16175 5729
rect 16206 5720 16212 5772
rect 16264 5760 16270 5772
rect 16264 5732 16309 5760
rect 16264 5720 16270 5732
rect 15488 5664 15976 5692
rect 15562 5624 15568 5636
rect 15304 5596 15568 5624
rect 15562 5584 15568 5596
rect 15620 5584 15626 5636
rect 15948 5624 15976 5664
rect 16025 5695 16083 5701
rect 16025 5661 16037 5695
rect 16071 5692 16083 5695
rect 16298 5692 16304 5704
rect 16071 5664 16304 5692
rect 16071 5661 16083 5664
rect 16025 5655 16083 5661
rect 16298 5652 16304 5664
rect 16356 5652 16362 5704
rect 18414 5624 18420 5636
rect 15948 5596 18420 5624
rect 18414 5584 18420 5596
rect 18472 5584 18478 5636
rect 18506 5556 18512 5568
rect 7116 5528 18512 5556
rect 18506 5516 18512 5528
rect 18564 5516 18570 5568
rect 1104 5466 19044 5488
rect 1104 5414 3972 5466
rect 4024 5414 4036 5466
rect 4088 5414 4100 5466
rect 4152 5414 4164 5466
rect 4216 5414 9952 5466
rect 10004 5414 10016 5466
rect 10068 5414 10080 5466
rect 10132 5414 10144 5466
rect 10196 5414 15932 5466
rect 15984 5414 15996 5466
rect 16048 5414 16060 5466
rect 16112 5414 16124 5466
rect 16176 5414 19044 5466
rect 1104 5392 19044 5414
rect 5905 5287 5963 5293
rect 5905 5253 5917 5287
rect 5951 5284 5963 5287
rect 5997 5287 6055 5293
rect 5997 5284 6009 5287
rect 5951 5256 6009 5284
rect 5951 5253 5963 5256
rect 5905 5247 5963 5253
rect 5997 5253 6009 5256
rect 6043 5253 6055 5287
rect 5997 5247 6055 5253
rect 16301 5219 16359 5225
rect 4908 5188 6224 5216
rect 2926 5151 2984 5157
rect 2926 5117 2938 5151
rect 2972 5148 2984 5151
rect 3234 5148 3240 5160
rect 2972 5120 3240 5148
rect 2972 5117 2984 5120
rect 2926 5111 2984 5117
rect 3234 5108 3240 5120
rect 3292 5108 3298 5160
rect 4706 5108 4712 5160
rect 4764 5148 4770 5160
rect 4908 5157 4936 5188
rect 4893 5151 4951 5157
rect 4893 5148 4905 5151
rect 4764 5120 4905 5148
rect 4764 5108 4770 5120
rect 4893 5117 4905 5120
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 5350 5108 5356 5160
rect 5408 5148 5414 5160
rect 6196 5157 6224 5188
rect 16301 5185 16313 5219
rect 16347 5216 16359 5219
rect 16390 5216 16396 5228
rect 16347 5188 16396 5216
rect 16347 5185 16359 5188
rect 16301 5179 16359 5185
rect 16390 5176 16396 5188
rect 16448 5176 16454 5228
rect 5445 5151 5503 5157
rect 5445 5148 5457 5151
rect 5408 5120 5457 5148
rect 5408 5108 5414 5120
rect 5445 5117 5457 5120
rect 5491 5148 5503 5151
rect 5537 5151 5595 5157
rect 5537 5148 5549 5151
rect 5491 5120 5549 5148
rect 5491 5117 5503 5120
rect 5445 5111 5503 5117
rect 5537 5117 5549 5120
rect 5583 5117 5595 5151
rect 5537 5111 5595 5117
rect 6181 5151 6239 5157
rect 6181 5117 6193 5151
rect 6227 5148 6239 5151
rect 6362 5148 6368 5160
rect 6227 5120 6368 5148
rect 6227 5117 6239 5120
rect 6181 5111 6239 5117
rect 6362 5108 6368 5120
rect 6420 5108 6426 5160
rect 12621 5151 12679 5157
rect 12621 5117 12633 5151
rect 12667 5148 12679 5151
rect 12710 5148 12716 5160
rect 12667 5120 12716 5148
rect 12667 5117 12679 5120
rect 12621 5111 12679 5117
rect 12710 5108 12716 5120
rect 12768 5108 12774 5160
rect 14274 5108 14280 5160
rect 14332 5148 14338 5160
rect 14826 5148 14832 5160
rect 14332 5120 14832 5148
rect 14332 5108 14338 5120
rect 14826 5108 14832 5120
rect 14884 5148 14890 5160
rect 15289 5151 15347 5157
rect 15289 5148 15301 5151
rect 14884 5120 15301 5148
rect 14884 5108 14890 5120
rect 15289 5117 15301 5120
rect 15335 5117 15347 5151
rect 15289 5111 15347 5117
rect 15473 5151 15531 5157
rect 15473 5117 15485 5151
rect 15519 5117 15531 5151
rect 15473 5111 15531 5117
rect 4985 5083 5043 5089
rect 4985 5049 4997 5083
rect 5031 5049 5043 5083
rect 12434 5080 12440 5092
rect 12395 5052 12440 5080
rect 4985 5043 5043 5049
rect 2406 4972 2412 5024
rect 2464 5012 2470 5024
rect 2823 5015 2881 5021
rect 2823 5012 2835 5015
rect 2464 4984 2835 5012
rect 2464 4972 2470 4984
rect 2823 4981 2835 4984
rect 2869 4981 2881 5015
rect 5000 5012 5028 5043
rect 12434 5040 12440 5052
rect 12492 5040 12498 5092
rect 15488 5080 15516 5111
rect 15562 5108 15568 5160
rect 15620 5148 15626 5160
rect 15657 5151 15715 5157
rect 15657 5148 15669 5151
rect 15620 5120 15669 5148
rect 15620 5108 15626 5120
rect 15657 5117 15669 5120
rect 15703 5148 15715 5151
rect 15841 5151 15899 5157
rect 15841 5148 15853 5151
rect 15703 5120 15853 5148
rect 15703 5117 15715 5120
rect 15657 5111 15715 5117
rect 15841 5117 15853 5120
rect 15887 5117 15899 5151
rect 16206 5148 16212 5160
rect 16167 5120 16212 5148
rect 15841 5111 15899 5117
rect 16206 5108 16212 5120
rect 16264 5108 16270 5160
rect 16224 5080 16252 5108
rect 15488 5052 16252 5080
rect 5902 5012 5908 5024
rect 5000 4984 5908 5012
rect 2823 4975 2881 4981
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 15654 5012 15660 5024
rect 15615 4984 15660 5012
rect 15654 4972 15660 4984
rect 15712 4972 15718 5024
rect 16393 5015 16451 5021
rect 16393 4981 16405 5015
rect 16439 5012 16451 5015
rect 16482 5012 16488 5024
rect 16439 4984 16488 5012
rect 16439 4981 16451 4984
rect 16393 4975 16451 4981
rect 16482 4972 16488 4984
rect 16540 4972 16546 5024
rect 1104 4922 19044 4944
rect 1104 4870 6962 4922
rect 7014 4870 7026 4922
rect 7078 4870 7090 4922
rect 7142 4870 7154 4922
rect 7206 4870 12942 4922
rect 12994 4870 13006 4922
rect 13058 4870 13070 4922
rect 13122 4870 13134 4922
rect 13186 4870 19044 4922
rect 1104 4848 19044 4870
rect 1486 4808 1492 4820
rect 1447 4780 1492 4808
rect 1486 4768 1492 4780
rect 1544 4768 1550 4820
rect 6362 4808 6368 4820
rect 6323 4780 6368 4808
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 7653 4811 7711 4817
rect 7653 4777 7665 4811
rect 7699 4777 7711 4811
rect 7653 4771 7711 4777
rect 3326 4740 3332 4752
rect 3287 4712 3332 4740
rect 3326 4700 3332 4712
rect 3384 4700 3390 4752
rect 6457 4743 6515 4749
rect 6457 4709 6469 4743
rect 6503 4740 6515 4743
rect 7668 4740 7696 4771
rect 10502 4768 10508 4820
rect 10560 4808 10566 4820
rect 11057 4811 11115 4817
rect 11057 4808 11069 4811
rect 10560 4780 11069 4808
rect 10560 4768 10566 4780
rect 11057 4777 11069 4780
rect 11103 4777 11115 4811
rect 11057 4771 11115 4777
rect 14734 4768 14740 4820
rect 14792 4808 14798 4820
rect 15013 4811 15071 4817
rect 15013 4808 15025 4811
rect 14792 4780 15025 4808
rect 14792 4768 14798 4780
rect 15013 4777 15025 4780
rect 15059 4777 15071 4811
rect 15013 4771 15071 4777
rect 15381 4811 15439 4817
rect 15381 4777 15393 4811
rect 15427 4808 15439 4811
rect 16025 4811 16083 4817
rect 16025 4808 16037 4811
rect 15427 4780 16037 4808
rect 15427 4777 15439 4780
rect 15381 4771 15439 4777
rect 16025 4777 16037 4780
rect 16071 4777 16083 4811
rect 18506 4808 18512 4820
rect 18467 4780 18512 4808
rect 16025 4771 16083 4777
rect 18506 4768 18512 4780
rect 18564 4768 18570 4820
rect 8018 4740 8024 4752
rect 6503 4712 8024 4740
rect 6503 4709 6515 4712
rect 6457 4703 6515 4709
rect 8018 4700 8024 4712
rect 8076 4700 8082 4752
rect 10060 4712 10732 4740
rect 1581 4675 1639 4681
rect 1581 4641 1593 4675
rect 1627 4641 1639 4675
rect 2406 4672 2412 4684
rect 2367 4644 2412 4672
rect 1581 4635 1639 4641
rect 1596 4604 1624 4635
rect 2406 4632 2412 4644
rect 2464 4632 2470 4684
rect 10060 4681 10088 4712
rect 10704 4684 10732 4712
rect 10778 4700 10784 4752
rect 10836 4740 10842 4752
rect 11146 4740 11152 4752
rect 10836 4712 11152 4740
rect 10836 4700 10842 4712
rect 11146 4700 11152 4712
rect 11204 4740 11210 4752
rect 11204 4712 11376 4740
rect 11204 4700 11210 4712
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4641 10103 4675
rect 10594 4672 10600 4684
rect 10555 4644 10600 4672
rect 10045 4635 10103 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 10686 4632 10692 4684
rect 10744 4672 10750 4684
rect 11348 4681 11376 4712
rect 16482 4700 16488 4752
rect 16540 4740 16546 4752
rect 16540 4700 16574 4740
rect 11333 4675 11391 4681
rect 10744 4644 10837 4672
rect 10744 4632 10750 4644
rect 11333 4641 11345 4675
rect 11379 4641 11391 4675
rect 11333 4635 11391 4641
rect 12158 4632 12164 4684
rect 12216 4672 12222 4684
rect 12253 4675 12311 4681
rect 12253 4672 12265 4675
rect 12216 4644 12265 4672
rect 12216 4632 12222 4644
rect 12253 4641 12265 4644
rect 12299 4641 12311 4675
rect 12253 4635 12311 4641
rect 16298 4632 16304 4684
rect 16356 4672 16362 4684
rect 16393 4675 16451 4681
rect 16393 4672 16405 4675
rect 16356 4644 16405 4672
rect 16356 4632 16362 4644
rect 16393 4641 16405 4644
rect 16439 4641 16451 4675
rect 16546 4672 16574 4700
rect 18690 4672 18696 4684
rect 16546 4644 16620 4672
rect 18651 4644 18696 4672
rect 16393 4635 16451 4641
rect 4430 4604 4436 4616
rect 1596 4576 4436 4604
rect 4430 4564 4436 4576
rect 4488 4564 4494 4616
rect 7282 4604 7288 4616
rect 7243 4576 7288 4604
rect 7282 4564 7288 4576
rect 7340 4564 7346 4616
rect 11606 4604 11612 4616
rect 7576 4576 10640 4604
rect 11567 4576 11612 4604
rect 3513 4539 3571 4545
rect 3513 4505 3525 4539
rect 3559 4536 3571 4539
rect 7576 4536 7604 4576
rect 3559 4508 7604 4536
rect 7653 4539 7711 4545
rect 3559 4505 3571 4508
rect 3513 4499 3571 4505
rect 7653 4505 7665 4539
rect 7699 4536 7711 4539
rect 8110 4536 8116 4548
rect 7699 4508 8116 4536
rect 7699 4505 7711 4508
rect 7653 4499 7711 4505
rect 8110 4496 8116 4508
rect 8168 4496 8174 4548
rect 10612 4536 10640 4576
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 15470 4604 15476 4616
rect 15431 4576 15476 4604
rect 15470 4564 15476 4576
rect 15528 4564 15534 4616
rect 15654 4604 15660 4616
rect 15615 4576 15660 4604
rect 15654 4564 15660 4576
rect 15712 4564 15718 4616
rect 16592 4613 16620 4644
rect 18690 4632 18696 4644
rect 18748 4632 18754 4684
rect 16485 4607 16543 4613
rect 16485 4604 16497 4607
rect 16408 4576 16497 4604
rect 16408 4548 16436 4576
rect 16485 4573 16497 4576
rect 16531 4573 16543 4607
rect 16485 4567 16543 4573
rect 16577 4607 16635 4613
rect 16577 4573 16589 4607
rect 16623 4573 16635 4607
rect 16577 4567 16635 4573
rect 11057 4539 11115 4545
rect 10612 4508 10732 4536
rect 2314 4468 2320 4480
rect 2275 4440 2320 4468
rect 2314 4428 2320 4440
rect 2372 4428 2378 4480
rect 10502 4428 10508 4480
rect 10560 4468 10566 4480
rect 10597 4471 10655 4477
rect 10597 4468 10609 4471
rect 10560 4440 10609 4468
rect 10560 4428 10566 4440
rect 10597 4437 10609 4440
rect 10643 4437 10655 4471
rect 10704 4468 10732 4508
rect 11057 4505 11069 4539
rect 11103 4536 11115 4539
rect 11149 4539 11207 4545
rect 11149 4536 11161 4539
rect 11103 4508 11161 4536
rect 11103 4505 11115 4508
rect 11057 4499 11115 4505
rect 11149 4505 11161 4508
rect 11195 4505 11207 4539
rect 11149 4499 11207 4505
rect 16390 4496 16396 4548
rect 16448 4536 16454 4548
rect 17954 4536 17960 4548
rect 16448 4508 17960 4536
rect 16448 4496 16454 4508
rect 17954 4496 17960 4508
rect 18012 4536 18018 4548
rect 18138 4536 18144 4548
rect 18012 4508 18144 4536
rect 18012 4496 18018 4508
rect 18138 4496 18144 4508
rect 18196 4496 18202 4548
rect 13078 4468 13084 4480
rect 10704 4440 13084 4468
rect 10597 4431 10655 4437
rect 13078 4428 13084 4440
rect 13136 4428 13142 4480
rect 1104 4378 19044 4400
rect 1104 4326 3972 4378
rect 4024 4326 4036 4378
rect 4088 4326 4100 4378
rect 4152 4326 4164 4378
rect 4216 4326 9952 4378
rect 10004 4326 10016 4378
rect 10068 4326 10080 4378
rect 10132 4326 10144 4378
rect 10196 4326 15932 4378
rect 15984 4326 15996 4378
rect 16048 4326 16060 4378
rect 16112 4326 16124 4378
rect 16176 4326 19044 4378
rect 1104 4304 19044 4326
rect 7282 4224 7288 4276
rect 7340 4264 7346 4276
rect 7653 4267 7711 4273
rect 7653 4264 7665 4267
rect 7340 4236 7665 4264
rect 7340 4224 7346 4236
rect 7653 4233 7665 4236
rect 7699 4264 7711 4267
rect 7742 4264 7748 4276
rect 7699 4236 7748 4264
rect 7699 4233 7711 4236
rect 7653 4227 7711 4233
rect 7742 4224 7748 4236
rect 7800 4224 7806 4276
rect 10597 4267 10655 4273
rect 10597 4233 10609 4267
rect 10643 4264 10655 4267
rect 10686 4264 10692 4276
rect 10643 4236 10692 4264
rect 10643 4233 10655 4236
rect 10597 4227 10655 4233
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 7190 4196 7196 4208
rect 7103 4168 7196 4196
rect 7116 4137 7144 4168
rect 7190 4156 7196 4168
rect 7248 4196 7254 4208
rect 11606 4196 11612 4208
rect 7248 4168 11612 4196
rect 7248 4156 7254 4168
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4097 7159 4131
rect 7101 4091 7159 4097
rect 8018 4088 8024 4140
rect 8076 4128 8082 4140
rect 9968 4137 9996 4168
rect 11606 4156 11612 4168
rect 11664 4156 11670 4208
rect 8113 4131 8171 4137
rect 8113 4128 8125 4131
rect 8076 4100 8125 4128
rect 8076 4088 8082 4100
rect 8113 4097 8125 4100
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 9953 4131 10011 4137
rect 9953 4097 9965 4131
rect 9999 4097 10011 4131
rect 11885 4131 11943 4137
rect 9953 4091 10011 4097
rect 10060 4100 10456 4128
rect 7285 4063 7343 4069
rect 7285 4029 7297 4063
rect 7331 4060 7343 4063
rect 7374 4060 7380 4072
rect 7331 4032 7380 4060
rect 7331 4029 7343 4032
rect 7285 4023 7343 4029
rect 7374 4020 7380 4032
rect 7432 4020 7438 4072
rect 7742 4060 7748 4072
rect 7703 4032 7748 4060
rect 7742 4020 7748 4032
rect 7800 4020 7806 4072
rect 8297 4063 8355 4069
rect 8297 4029 8309 4063
rect 8343 4060 8355 4063
rect 8570 4060 8576 4072
rect 8343 4032 8576 4060
rect 8343 4029 8355 4032
rect 8297 4023 8355 4029
rect 8570 4020 8576 4032
rect 8628 4060 8634 4072
rect 10060 4060 10088 4100
rect 8628 4032 10088 4060
rect 10229 4063 10287 4069
rect 8628 4020 8634 4032
rect 10229 4029 10241 4063
rect 10275 4060 10287 4063
rect 10318 4060 10324 4072
rect 10275 4032 10324 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 10318 4020 10324 4032
rect 10376 4020 10382 4072
rect 10428 4060 10456 4100
rect 11885 4097 11897 4131
rect 11931 4128 11943 4131
rect 12158 4128 12164 4140
rect 11931 4100 12164 4128
rect 11931 4097 11943 4100
rect 11885 4091 11943 4097
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 12434 4128 12440 4140
rect 12406 4088 12440 4128
rect 12492 4088 12498 4140
rect 13173 4131 13231 4137
rect 13173 4128 13185 4131
rect 12544 4100 13185 4128
rect 12406 4060 12434 4088
rect 12544 4069 12572 4100
rect 13173 4097 13185 4100
rect 13219 4097 13231 4131
rect 13722 4128 13728 4140
rect 13173 4091 13231 4097
rect 13464 4100 13728 4128
rect 10428 4032 12434 4060
rect 12529 4063 12587 4069
rect 12529 4029 12541 4063
rect 12575 4029 12587 4063
rect 13078 4060 13084 4072
rect 13039 4032 13084 4060
rect 12529 4023 12587 4029
rect 6546 3952 6552 4004
rect 6604 3992 6610 4004
rect 10137 3995 10195 4001
rect 6604 3964 10088 3992
rect 6604 3952 6610 3964
rect 7193 3927 7251 3933
rect 7193 3893 7205 3927
rect 7239 3924 7251 3927
rect 9766 3924 9772 3936
rect 7239 3896 9772 3924
rect 7239 3893 7251 3896
rect 7193 3887 7251 3893
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 10060 3924 10088 3964
rect 10137 3961 10149 3995
rect 10183 3992 10195 3995
rect 10594 3992 10600 4004
rect 10183 3964 10600 3992
rect 10183 3961 10195 3964
rect 10137 3955 10195 3961
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 11238 3952 11244 4004
rect 11296 3992 11302 4004
rect 12069 3995 12127 4001
rect 12069 3992 12081 3995
rect 11296 3964 12081 3992
rect 11296 3952 11302 3964
rect 12069 3961 12081 3964
rect 12115 3961 12127 3995
rect 12069 3955 12127 3961
rect 11330 3924 11336 3936
rect 10060 3896 11336 3924
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11974 3924 11980 3936
rect 11935 3896 11980 3924
rect 11974 3884 11980 3896
rect 12032 3884 12038 3936
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3924 12495 3927
rect 12544 3924 12572 4023
rect 13078 4020 13084 4032
rect 13136 4060 13142 4072
rect 13464 4060 13492 4100
rect 13722 4088 13728 4100
rect 13780 4128 13786 4140
rect 13780 4100 13860 4128
rect 13780 4088 13786 4100
rect 13832 4069 13860 4100
rect 13136 4032 13492 4060
rect 13541 4063 13599 4069
rect 13136 4020 13142 4032
rect 13541 4029 13553 4063
rect 13587 4060 13599 4063
rect 13817 4063 13875 4069
rect 13587 4032 13676 4060
rect 13587 4029 13599 4032
rect 13541 4023 13599 4029
rect 12989 3995 13047 4001
rect 12989 3961 13001 3995
rect 13035 3992 13047 3995
rect 13035 3964 13584 3992
rect 13035 3961 13047 3964
rect 12989 3955 13047 3961
rect 13556 3936 13584 3964
rect 13538 3924 13544 3936
rect 12483 3896 12572 3924
rect 13451 3896 13544 3924
rect 12483 3893 12495 3896
rect 12437 3887 12495 3893
rect 13538 3884 13544 3896
rect 13596 3884 13602 3936
rect 13648 3933 13676 4032
rect 13817 4029 13829 4063
rect 13863 4029 13875 4063
rect 13817 4023 13875 4029
rect 13633 3927 13691 3933
rect 13633 3893 13645 3927
rect 13679 3893 13691 3927
rect 13633 3887 13691 3893
rect 1104 3834 19044 3856
rect 1104 3782 6962 3834
rect 7014 3782 7026 3834
rect 7078 3782 7090 3834
rect 7142 3782 7154 3834
rect 7206 3782 12942 3834
rect 12994 3782 13006 3834
rect 13058 3782 13070 3834
rect 13122 3782 13134 3834
rect 13186 3782 19044 3834
rect 1104 3760 19044 3782
rect 11146 3720 11152 3732
rect 5920 3692 8248 3720
rect 11107 3692 11152 3720
rect 5920 3664 5948 3692
rect 5902 3652 5908 3664
rect 5566 3624 5908 3652
rect 5902 3612 5908 3624
rect 5960 3612 5966 3664
rect 5997 3655 6055 3661
rect 5997 3621 6009 3655
rect 6043 3652 6055 3655
rect 8110 3652 8116 3664
rect 6043 3624 6408 3652
rect 8071 3624 8116 3652
rect 6043 3621 6055 3624
rect 5997 3615 6055 3621
rect 6273 3519 6331 3525
rect 6273 3516 6285 3519
rect 4908 3488 6285 3516
rect 4908 3460 4936 3488
rect 6273 3485 6285 3488
rect 6319 3485 6331 3519
rect 6273 3479 6331 3485
rect 6380 3516 6408 3624
rect 8110 3612 8116 3624
rect 8168 3612 8174 3664
rect 8220 3652 8248 3692
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 13538 3680 13544 3732
rect 13596 3720 13602 3732
rect 13909 3723 13967 3729
rect 13909 3720 13921 3723
rect 13596 3692 13921 3720
rect 13596 3680 13602 3692
rect 13909 3689 13921 3692
rect 13955 3689 13967 3723
rect 13909 3683 13967 3689
rect 15378 3652 15384 3664
rect 8220 3624 15384 3652
rect 15378 3612 15384 3624
rect 15436 3652 15442 3664
rect 15436 3624 16330 3652
rect 15436 3612 15442 3624
rect 8297 3587 8355 3593
rect 8297 3553 8309 3587
rect 8343 3584 8355 3587
rect 8386 3584 8392 3596
rect 8343 3556 8392 3584
rect 8343 3553 8355 3556
rect 8297 3547 8355 3553
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 10962 3544 10968 3596
rect 11020 3584 11026 3596
rect 11057 3587 11115 3593
rect 11057 3584 11069 3587
rect 11020 3556 11069 3584
rect 11020 3544 11026 3556
rect 11057 3553 11069 3556
rect 11103 3553 11115 3587
rect 11057 3547 11115 3553
rect 11330 3544 11336 3596
rect 11388 3584 11394 3596
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 11388 3556 14749 3584
rect 11388 3544 11394 3556
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 17589 3587 17647 3593
rect 17589 3553 17601 3587
rect 17635 3584 17647 3587
rect 17862 3584 17868 3596
rect 17635 3556 17868 3584
rect 17635 3553 17647 3556
rect 17589 3547 17647 3553
rect 17862 3544 17868 3556
rect 17920 3544 17926 3596
rect 14826 3516 14832 3528
rect 6380 3488 14688 3516
rect 14787 3488 14832 3516
rect 4890 3408 4896 3460
rect 4948 3408 4954 3460
rect 4265 3383 4323 3389
rect 4265 3349 4277 3383
rect 4311 3380 4323 3383
rect 4430 3380 4436 3392
rect 4311 3352 4436 3380
rect 4311 3349 4323 3352
rect 4265 3343 4323 3349
rect 4430 3340 4436 3352
rect 4488 3380 4494 3392
rect 6380 3380 6408 3488
rect 9766 3408 9772 3460
rect 9824 3448 9830 3460
rect 14660 3448 14688 3488
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 15010 3516 15016 3528
rect 14971 3488 15016 3516
rect 15010 3476 15016 3488
rect 15068 3476 15074 3528
rect 15565 3519 15623 3525
rect 15565 3485 15577 3519
rect 15611 3485 15623 3519
rect 15565 3479 15623 3485
rect 15841 3519 15899 3525
rect 15841 3485 15853 3519
rect 15887 3516 15899 3519
rect 16390 3516 16396 3528
rect 15887 3488 16396 3516
rect 15887 3485 15899 3488
rect 15841 3479 15899 3485
rect 15470 3448 15476 3460
rect 9824 3420 14504 3448
rect 14660 3420 15476 3448
rect 9824 3408 9830 3420
rect 13998 3380 14004 3392
rect 4488 3352 6408 3380
rect 13959 3352 14004 3380
rect 4488 3340 4494 3352
rect 13998 3340 14004 3352
rect 14056 3340 14062 3392
rect 14366 3380 14372 3392
rect 14327 3352 14372 3380
rect 14366 3340 14372 3352
rect 14424 3340 14430 3392
rect 14476 3380 14504 3420
rect 15470 3408 15476 3420
rect 15528 3448 15534 3460
rect 15580 3448 15608 3479
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 15528 3420 15608 3448
rect 15528 3408 15534 3420
rect 18506 3380 18512 3392
rect 14476 3352 18512 3380
rect 18506 3340 18512 3352
rect 18564 3340 18570 3392
rect 1104 3290 19044 3312
rect 1104 3238 3972 3290
rect 4024 3238 4036 3290
rect 4088 3238 4100 3290
rect 4152 3238 4164 3290
rect 4216 3238 9952 3290
rect 10004 3238 10016 3290
rect 10068 3238 10080 3290
rect 10132 3238 10144 3290
rect 10196 3238 15932 3290
rect 15984 3238 15996 3290
rect 16048 3238 16060 3290
rect 16112 3238 16124 3290
rect 16176 3238 19044 3290
rect 1104 3216 19044 3238
rect 5902 3176 5908 3188
rect 5863 3148 5908 3176
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 8386 3176 8392 3188
rect 8347 3148 8392 3176
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 9585 3179 9643 3185
rect 9585 3145 9597 3179
rect 9631 3176 9643 3179
rect 10410 3176 10416 3188
rect 9631 3148 10416 3176
rect 9631 3145 9643 3148
rect 9585 3139 9643 3145
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 10505 3179 10563 3185
rect 10505 3145 10517 3179
rect 10551 3176 10563 3179
rect 10962 3176 10968 3188
rect 10551 3148 10968 3176
rect 10551 3145 10563 3148
rect 10505 3139 10563 3145
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 12069 3179 12127 3185
rect 12069 3176 12081 3179
rect 11992 3148 12081 3176
rect 4890 3108 4896 3120
rect 4356 3080 4896 3108
rect 2314 3000 2320 3052
rect 2372 3040 2378 3052
rect 3053 3043 3111 3049
rect 3053 3040 3065 3043
rect 2372 3012 3065 3040
rect 2372 3000 2378 3012
rect 3053 3009 3065 3012
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3040 3387 3043
rect 4356 3040 4384 3080
rect 4890 3068 4896 3080
rect 4948 3108 4954 3120
rect 5031 3111 5089 3117
rect 5031 3108 5043 3111
rect 4948 3080 5043 3108
rect 4948 3068 4954 3080
rect 5031 3077 5043 3080
rect 5077 3077 5089 3111
rect 5031 3071 5089 3077
rect 5920 3040 5948 3136
rect 8849 3111 8907 3117
rect 8849 3077 8861 3111
rect 8895 3108 8907 3111
rect 8941 3111 8999 3117
rect 8941 3108 8953 3111
rect 8895 3080 8953 3108
rect 8895 3077 8907 3080
rect 8849 3071 8907 3077
rect 8941 3077 8953 3080
rect 8987 3077 8999 3111
rect 8941 3071 8999 3077
rect 8570 3040 8576 3052
rect 3375 3012 4384 3040
rect 4448 3012 5948 3040
rect 8404 3012 8576 3040
rect 3375 3009 3387 3012
rect 3329 3003 3387 3009
rect 1394 2972 1400 2984
rect 1355 2944 1400 2972
rect 1394 2932 1400 2944
rect 1452 2932 1458 2984
rect 4448 2958 4476 3012
rect 5718 2932 5724 2984
rect 5776 2972 5782 2984
rect 8404 2981 8432 3012
rect 8570 3000 8576 3012
rect 8628 3040 8634 3052
rect 10597 3043 10655 3049
rect 10597 3040 10609 3043
rect 8628 3012 9168 3040
rect 8628 3000 8634 3012
rect 9140 2981 9168 3012
rect 9968 3012 10609 3040
rect 9968 2984 9996 3012
rect 10597 3009 10609 3012
rect 10643 3009 10655 3043
rect 10597 3003 10655 3009
rect 5813 2975 5871 2981
rect 5813 2972 5825 2975
rect 5776 2944 5825 2972
rect 5776 2932 5782 2944
rect 5813 2941 5825 2944
rect 5859 2941 5871 2975
rect 5813 2935 5871 2941
rect 7837 2975 7895 2981
rect 7837 2941 7849 2975
rect 7883 2941 7895 2975
rect 7837 2935 7895 2941
rect 8389 2975 8447 2981
rect 8389 2941 8401 2975
rect 8435 2941 8447 2975
rect 8389 2935 8447 2941
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2941 8539 2975
rect 8481 2935 8539 2941
rect 9125 2975 9183 2981
rect 9125 2941 9137 2975
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 7852 2904 7880 2935
rect 8294 2904 8300 2916
rect 5368 2876 6040 2904
rect 7852 2876 8300 2904
rect 1581 2839 1639 2845
rect 1581 2805 1593 2839
rect 1627 2836 1639 2839
rect 5368 2836 5396 2876
rect 1627 2808 5396 2836
rect 6012 2836 6040 2876
rect 8294 2864 8300 2876
rect 8352 2904 8358 2916
rect 8496 2904 8524 2935
rect 9306 2932 9312 2984
rect 9364 2972 9370 2984
rect 9493 2975 9551 2981
rect 9493 2972 9505 2975
rect 9364 2944 9505 2972
rect 9364 2932 9370 2944
rect 9493 2941 9505 2944
rect 9539 2941 9551 2975
rect 9950 2972 9956 2984
rect 9863 2944 9956 2972
rect 9493 2935 9551 2941
rect 9950 2932 9956 2944
rect 10008 2932 10014 2984
rect 11992 2981 12020 3148
rect 12069 3145 12081 3148
rect 12115 3176 12127 3179
rect 13081 3179 13139 3185
rect 13081 3176 13093 3179
rect 12115 3148 13093 3176
rect 12115 3145 12127 3148
rect 12069 3139 12127 3145
rect 13081 3145 13093 3148
rect 13127 3145 13139 3179
rect 13081 3139 13139 3145
rect 14826 3136 14832 3188
rect 14884 3176 14890 3188
rect 18509 3179 18567 3185
rect 18509 3176 18521 3179
rect 14884 3148 18521 3176
rect 14884 3136 14890 3148
rect 18509 3145 18521 3148
rect 18555 3145 18567 3179
rect 18509 3139 18567 3145
rect 12158 3068 12164 3120
rect 12216 3108 12222 3120
rect 15010 3108 15016 3120
rect 12216 3080 15016 3108
rect 12216 3068 12222 3080
rect 15010 3068 15016 3080
rect 15068 3068 15074 3120
rect 12713 3043 12771 3049
rect 12713 3040 12725 3043
rect 12636 3012 12725 3040
rect 12636 2981 12664 3012
rect 12713 3009 12725 3012
rect 12759 3040 12771 3043
rect 12802 3040 12808 3052
rect 12759 3012 12808 3040
rect 12759 3009 12771 3012
rect 12713 3003 12771 3009
rect 12802 3000 12808 3012
rect 12860 3000 12866 3052
rect 16390 3000 16396 3052
rect 16448 3040 16454 3052
rect 16761 3043 16819 3049
rect 16761 3040 16773 3043
rect 16448 3012 16773 3040
rect 16448 3000 16454 3012
rect 16761 3009 16773 3012
rect 16807 3009 16819 3043
rect 16761 3003 16819 3009
rect 10505 2975 10563 2981
rect 10505 2941 10517 2975
rect 10551 2941 10563 2975
rect 10505 2935 10563 2941
rect 10965 2975 11023 2981
rect 10965 2941 10977 2975
rect 11011 2972 11023 2975
rect 11793 2975 11851 2981
rect 11793 2972 11805 2975
rect 11011 2944 11805 2972
rect 11011 2941 11023 2944
rect 10965 2935 11023 2941
rect 11793 2941 11805 2944
rect 11839 2941 11851 2975
rect 11793 2935 11851 2941
rect 11977 2975 12035 2981
rect 11977 2941 11989 2975
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 12069 2975 12127 2981
rect 12069 2941 12081 2975
rect 12115 2972 12127 2975
rect 12621 2975 12679 2981
rect 12115 2944 12434 2972
rect 12115 2941 12127 2944
rect 12069 2935 12127 2941
rect 8352 2876 8524 2904
rect 10520 2904 10548 2935
rect 12084 2904 12112 2935
rect 10520 2876 12112 2904
rect 12406 2904 12434 2944
rect 12621 2941 12633 2975
rect 12667 2941 12679 2975
rect 12621 2935 12679 2941
rect 13081 2975 13139 2981
rect 13081 2941 13093 2975
rect 13127 2972 13139 2975
rect 13262 2972 13268 2984
rect 13127 2944 13268 2972
rect 13127 2941 13139 2944
rect 13081 2935 13139 2941
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 13722 2972 13728 2984
rect 13683 2944 13728 2972
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 14277 2975 14335 2981
rect 14277 2941 14289 2975
rect 14323 2972 14335 2975
rect 14366 2972 14372 2984
rect 14323 2944 14372 2972
rect 14323 2941 14335 2944
rect 14277 2935 14335 2941
rect 14366 2932 14372 2944
rect 14424 2932 14430 2984
rect 15378 2932 15384 2984
rect 15436 2932 15442 2984
rect 18690 2972 18696 2984
rect 18651 2944 18696 2972
rect 18690 2932 18696 2944
rect 18748 2932 18754 2984
rect 13814 2904 13820 2916
rect 12406 2876 12848 2904
rect 13775 2876 13820 2904
rect 8352 2864 8358 2876
rect 12820 2848 12848 2876
rect 13814 2864 13820 2876
rect 13872 2904 13878 2916
rect 14553 2907 14611 2913
rect 14553 2904 14565 2907
rect 13872 2876 14565 2904
rect 13872 2864 13878 2876
rect 14553 2873 14565 2876
rect 14599 2873 14611 2907
rect 14553 2867 14611 2873
rect 16390 2864 16396 2916
rect 16448 2904 16454 2916
rect 16485 2907 16543 2913
rect 16485 2904 16497 2907
rect 16448 2876 16497 2904
rect 16448 2864 16454 2876
rect 16485 2873 16497 2876
rect 16531 2873 16543 2907
rect 16485 2867 16543 2873
rect 7926 2836 7932 2848
rect 6012 2808 7932 2836
rect 1627 2805 1639 2808
rect 1581 2799 1639 2805
rect 7926 2796 7932 2808
rect 7984 2796 7990 2848
rect 8478 2796 8484 2848
rect 8536 2836 8542 2848
rect 8849 2839 8907 2845
rect 8849 2836 8861 2839
rect 8536 2808 8861 2836
rect 8536 2796 8542 2808
rect 8849 2805 8861 2808
rect 8895 2805 8907 2839
rect 8849 2799 8907 2805
rect 12802 2796 12808 2848
rect 12860 2836 12866 2848
rect 14461 2839 14519 2845
rect 14461 2836 14473 2839
rect 12860 2808 14473 2836
rect 12860 2796 12866 2808
rect 14461 2805 14473 2808
rect 14507 2805 14519 2839
rect 14461 2799 14519 2805
rect 14737 2839 14795 2845
rect 14737 2805 14749 2839
rect 14783 2836 14795 2839
rect 16408 2836 16436 2864
rect 14783 2808 16436 2836
rect 14783 2805 14795 2808
rect 14737 2799 14795 2805
rect 1104 2746 19044 2768
rect 1104 2694 6962 2746
rect 7014 2694 7026 2746
rect 7078 2694 7090 2746
rect 7142 2694 7154 2746
rect 7206 2694 12942 2746
rect 12994 2694 13006 2746
rect 13058 2694 13070 2746
rect 13122 2694 13134 2746
rect 13186 2694 19044 2746
rect 1104 2672 19044 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 3418 2632 3424 2644
rect 1627 2604 3280 2632
rect 3379 2604 3424 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 2041 2567 2099 2573
rect 2041 2533 2053 2567
rect 2087 2564 2099 2567
rect 2314 2564 2320 2576
rect 2087 2536 2320 2564
rect 2087 2533 2099 2536
rect 2041 2527 2099 2533
rect 2314 2524 2320 2536
rect 2372 2524 2378 2576
rect 3252 2564 3280 2604
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 4798 2632 4804 2644
rect 4759 2604 4804 2632
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 5718 2592 5724 2644
rect 5776 2632 5782 2644
rect 5997 2635 6055 2641
rect 5997 2632 6009 2635
rect 5776 2604 6009 2632
rect 5776 2592 5782 2604
rect 5997 2601 6009 2604
rect 6043 2601 6055 2635
rect 7926 2632 7932 2644
rect 7887 2604 7932 2632
rect 5997 2595 6055 2601
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 8389 2635 8447 2641
rect 8389 2632 8401 2635
rect 8352 2604 8401 2632
rect 8352 2592 8358 2604
rect 8389 2601 8401 2604
rect 8435 2601 8447 2635
rect 8389 2595 8447 2601
rect 8665 2635 8723 2641
rect 8665 2601 8677 2635
rect 8711 2632 8723 2635
rect 9493 2635 9551 2641
rect 9493 2632 9505 2635
rect 8711 2604 9505 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 9493 2601 9505 2604
rect 9539 2601 9551 2635
rect 9493 2595 9551 2601
rect 9582 2592 9588 2644
rect 9640 2632 9646 2644
rect 9950 2632 9956 2644
rect 9640 2604 9685 2632
rect 9911 2604 9956 2632
rect 9640 2592 9646 2604
rect 9950 2592 9956 2604
rect 10008 2592 10014 2644
rect 10594 2632 10600 2644
rect 10555 2604 10600 2632
rect 10594 2592 10600 2604
rect 10652 2592 10658 2644
rect 11974 2592 11980 2644
rect 12032 2632 12038 2644
rect 12161 2635 12219 2641
rect 12161 2632 12173 2635
rect 12032 2604 12173 2632
rect 12032 2592 12038 2604
rect 12161 2601 12173 2604
rect 12207 2601 12219 2635
rect 12161 2595 12219 2601
rect 12989 2635 13047 2641
rect 12989 2601 13001 2635
rect 13035 2632 13047 2635
rect 13262 2632 13268 2644
rect 13035 2604 13268 2632
rect 13035 2601 13047 2604
rect 12989 2595 13047 2601
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 13814 2592 13820 2644
rect 13872 2632 13878 2644
rect 14001 2635 14059 2641
rect 14001 2632 14013 2635
rect 13872 2604 14013 2632
rect 13872 2592 13878 2604
rect 14001 2601 14013 2604
rect 14047 2601 14059 2635
rect 15562 2632 15568 2644
rect 15523 2604 15568 2632
rect 14001 2595 14059 2601
rect 15562 2592 15568 2604
rect 15620 2592 15626 2644
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 18506 2632 18512 2644
rect 16632 2604 16677 2632
rect 18467 2604 18512 2632
rect 16632 2592 16638 2604
rect 18506 2592 18512 2604
rect 18564 2592 18570 2644
rect 9306 2564 9312 2576
rect 3252 2536 9312 2564
rect 9306 2524 9312 2536
rect 9364 2524 9370 2576
rect 10321 2567 10379 2573
rect 10321 2533 10333 2567
rect 10367 2564 10379 2567
rect 14274 2564 14280 2576
rect 10367 2536 14280 2564
rect 10367 2533 10379 2536
rect 10321 2527 10379 2533
rect 14274 2524 14280 2536
rect 14332 2524 14338 2576
rect 15010 2564 15016 2576
rect 14971 2536 15016 2564
rect 15010 2524 15016 2536
rect 15068 2524 15074 2576
rect 15194 2524 15200 2576
rect 15252 2564 15258 2576
rect 15473 2567 15531 2573
rect 15473 2564 15485 2567
rect 15252 2536 15485 2564
rect 15252 2524 15258 2536
rect 15473 2533 15485 2536
rect 15519 2533 15531 2567
rect 15473 2527 15531 2533
rect 16390 2524 16396 2576
rect 16448 2564 16454 2576
rect 18141 2567 18199 2573
rect 18141 2564 18153 2567
rect 16448 2536 18153 2564
rect 16448 2524 16454 2536
rect 18141 2533 18153 2536
rect 18187 2533 18199 2567
rect 18141 2527 18199 2533
rect 474 2456 480 2508
rect 532 2496 538 2508
rect 1397 2499 1455 2505
rect 1397 2496 1409 2499
rect 532 2468 1409 2496
rect 532 2456 538 2468
rect 1397 2465 1409 2468
rect 1443 2465 1455 2499
rect 3234 2496 3240 2508
rect 3195 2468 3240 2496
rect 1397 2459 1455 2465
rect 3234 2456 3240 2468
rect 3292 2456 3298 2508
rect 4614 2496 4620 2508
rect 4575 2468 4620 2496
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 5994 2456 6000 2508
rect 6052 2496 6058 2508
rect 6181 2499 6239 2505
rect 6181 2496 6193 2499
rect 6052 2468 6193 2496
rect 6052 2456 6058 2468
rect 6181 2465 6193 2468
rect 6227 2465 6239 2499
rect 6181 2459 6239 2465
rect 8021 2499 8079 2505
rect 8021 2465 8033 2499
rect 8067 2496 8079 2499
rect 8386 2496 8392 2508
rect 8067 2468 8392 2496
rect 8067 2465 8079 2468
rect 8021 2459 8079 2465
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 8481 2499 8539 2505
rect 8481 2465 8493 2499
rect 8527 2465 8539 2499
rect 8481 2459 8539 2465
rect 7282 2388 7288 2440
rect 7340 2428 7346 2440
rect 7745 2431 7803 2437
rect 7745 2428 7757 2431
rect 7340 2400 7757 2428
rect 7340 2388 7346 2400
rect 7745 2397 7757 2400
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 1854 2360 1860 2372
rect 1815 2332 1860 2360
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 7760 2360 7788 2391
rect 7834 2388 7840 2440
rect 7892 2428 7898 2440
rect 8496 2428 8524 2459
rect 9214 2456 9220 2508
rect 9272 2496 9278 2508
rect 10137 2499 10195 2505
rect 10137 2496 10149 2499
rect 9272 2468 10149 2496
rect 9272 2456 9278 2468
rect 10137 2465 10149 2468
rect 10183 2465 10195 2499
rect 10137 2459 10195 2465
rect 10594 2456 10600 2508
rect 10652 2496 10658 2508
rect 10781 2499 10839 2505
rect 10781 2496 10793 2499
rect 10652 2468 10793 2496
rect 10652 2456 10658 2468
rect 10781 2465 10793 2468
rect 10827 2465 10839 2499
rect 11974 2496 11980 2508
rect 11935 2468 11980 2496
rect 10781 2459 10839 2465
rect 11974 2456 11980 2468
rect 12032 2456 12038 2508
rect 12802 2496 12808 2508
rect 12763 2468 12808 2496
rect 12802 2456 12808 2468
rect 12860 2456 12866 2508
rect 13998 2496 14004 2508
rect 13959 2468 14004 2496
rect 13998 2456 14004 2468
rect 14056 2456 14062 2508
rect 14366 2496 14372 2508
rect 14327 2468 14372 2496
rect 14366 2456 14372 2468
rect 14424 2456 14430 2508
rect 14645 2499 14703 2505
rect 14645 2465 14657 2499
rect 14691 2465 14703 2499
rect 14645 2459 14703 2465
rect 7892 2400 8524 2428
rect 9309 2431 9367 2437
rect 7892 2388 7898 2400
rect 9309 2397 9321 2431
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 9324 2360 9352 2391
rect 13814 2388 13820 2440
rect 13872 2428 13878 2440
rect 14660 2428 14688 2459
rect 16574 2456 16580 2508
rect 16632 2496 16638 2508
rect 16761 2499 16819 2505
rect 16761 2496 16773 2499
rect 16632 2468 16773 2496
rect 16632 2456 16638 2468
rect 16761 2465 16773 2468
rect 16807 2465 16819 2499
rect 16761 2459 16819 2465
rect 18693 2499 18751 2505
rect 18693 2465 18705 2499
rect 18739 2496 18751 2499
rect 19153 2499 19211 2505
rect 19153 2496 19165 2499
rect 18739 2468 19165 2496
rect 18739 2465 18751 2468
rect 18693 2459 18751 2465
rect 19153 2465 19165 2468
rect 19199 2465 19211 2499
rect 19153 2459 19211 2465
rect 13872 2400 14688 2428
rect 13872 2388 13878 2400
rect 17954 2360 17960 2372
rect 7760 2332 9352 2360
rect 17915 2332 17960 2360
rect 17954 2320 17960 2332
rect 18012 2320 18018 2372
rect 1104 2202 19044 2224
rect 1104 2150 3972 2202
rect 4024 2150 4036 2202
rect 4088 2150 4100 2202
rect 4152 2150 4164 2202
rect 4216 2150 9952 2202
rect 10004 2150 10016 2202
rect 10068 2150 10080 2202
rect 10132 2150 10144 2202
rect 10196 2150 15932 2202
rect 15984 2150 15996 2202
rect 16048 2150 16060 2202
rect 16112 2150 16124 2202
rect 16176 2150 19044 2202
rect 1104 2128 19044 2150
rect 19150 1408 19156 1420
rect 19111 1380 19156 1408
rect 19150 1368 19156 1380
rect 19208 1368 19214 1420
<< via1 >>
rect 6962 20102 7014 20154
rect 7026 20102 7078 20154
rect 7090 20102 7142 20154
rect 7154 20102 7206 20154
rect 12942 20102 12994 20154
rect 13006 20102 13058 20154
rect 13070 20102 13122 20154
rect 13134 20102 13186 20154
rect 1492 20043 1544 20052
rect 1492 20009 1501 20043
rect 1501 20009 1535 20043
rect 1535 20009 1544 20043
rect 1492 20000 1544 20009
rect 940 19932 992 19984
rect 1584 19907 1636 19916
rect 1584 19873 1593 19907
rect 1593 19873 1627 19907
rect 1627 19873 1636 19907
rect 1584 19864 1636 19873
rect 18880 19932 18932 19984
rect 2320 19907 2372 19916
rect 2320 19873 2329 19907
rect 2329 19873 2363 19907
rect 2363 19873 2372 19907
rect 2320 19864 2372 19873
rect 3700 19864 3752 19916
rect 5540 19907 5592 19916
rect 5540 19873 5549 19907
rect 5549 19873 5583 19907
rect 5583 19873 5592 19907
rect 5540 19864 5592 19873
rect 6920 19907 6972 19916
rect 6920 19873 6929 19907
rect 6929 19873 6963 19907
rect 6963 19873 6972 19907
rect 6920 19864 6972 19873
rect 8300 19907 8352 19916
rect 8300 19873 8309 19907
rect 8309 19873 8343 19907
rect 8343 19873 8352 19907
rect 8300 19864 8352 19873
rect 9680 19864 9732 19916
rect 11520 19864 11572 19916
rect 12808 19864 12860 19916
rect 14280 19864 14332 19916
rect 15660 19864 15712 19916
rect 17500 19864 17552 19916
rect 18328 19907 18380 19916
rect 18328 19873 18337 19907
rect 18337 19873 18371 19907
rect 18371 19873 18380 19907
rect 18328 19864 18380 19873
rect 9588 19728 9640 19780
rect 13636 19728 13688 19780
rect 18420 19771 18472 19780
rect 18420 19737 18429 19771
rect 18429 19737 18463 19771
rect 18463 19737 18472 19771
rect 18420 19728 18472 19737
rect 1952 19703 2004 19712
rect 1952 19669 1961 19703
rect 1961 19669 1995 19703
rect 1995 19669 2004 19703
rect 1952 19660 2004 19669
rect 2504 19703 2556 19712
rect 2504 19669 2513 19703
rect 2513 19669 2547 19703
rect 2547 19669 2556 19703
rect 2504 19660 2556 19669
rect 3700 19660 3752 19712
rect 6000 19660 6052 19712
rect 8392 19660 8444 19712
rect 10508 19660 10560 19712
rect 11612 19660 11664 19712
rect 11888 19660 11940 19712
rect 14372 19660 14424 19712
rect 15660 19703 15712 19712
rect 15660 19669 15669 19703
rect 15669 19669 15703 19703
rect 15703 19669 15712 19703
rect 15660 19660 15712 19669
rect 17500 19703 17552 19712
rect 17500 19669 17509 19703
rect 17509 19669 17543 19703
rect 17543 19669 17552 19703
rect 17500 19660 17552 19669
rect 3972 19558 4024 19610
rect 4036 19558 4088 19610
rect 4100 19558 4152 19610
rect 4164 19558 4216 19610
rect 9952 19558 10004 19610
rect 10016 19558 10068 19610
rect 10080 19558 10132 19610
rect 10144 19558 10196 19610
rect 15932 19558 15984 19610
rect 15996 19558 16048 19610
rect 16060 19558 16112 19610
rect 16124 19558 16176 19610
rect 1584 19456 1636 19508
rect 3884 19320 3936 19372
rect 1860 19295 1912 19304
rect 1860 19261 1869 19295
rect 1869 19261 1903 19295
rect 1903 19261 1912 19295
rect 1860 19252 1912 19261
rect 8852 19320 8904 19372
rect 11244 19320 11296 19372
rect 17316 19320 17368 19372
rect 3424 19184 3476 19236
rect 4804 19184 4856 19236
rect 5816 19184 5868 19236
rect 6460 19184 6512 19236
rect 8208 19252 8260 19304
rect 7288 19227 7340 19236
rect 4436 19116 4488 19168
rect 7288 19193 7297 19227
rect 7297 19193 7331 19227
rect 7331 19193 7340 19227
rect 7288 19184 7340 19193
rect 9128 19184 9180 19236
rect 7564 19116 7616 19168
rect 7932 19116 7984 19168
rect 8208 19116 8260 19168
rect 10600 19184 10652 19236
rect 12624 19252 12676 19304
rect 15016 19252 15068 19304
rect 11520 19116 11572 19168
rect 12808 19116 12860 19168
rect 13820 19184 13872 19236
rect 17224 19252 17276 19304
rect 13728 19116 13780 19168
rect 15476 19159 15528 19168
rect 15476 19125 15485 19159
rect 15485 19125 15519 19159
rect 15519 19125 15528 19159
rect 15476 19116 15528 19125
rect 17040 19116 17092 19168
rect 18052 19116 18104 19168
rect 6962 19014 7014 19066
rect 7026 19014 7078 19066
rect 7090 19014 7142 19066
rect 7154 19014 7206 19066
rect 12942 19014 12994 19066
rect 13006 19014 13058 19066
rect 13070 19014 13122 19066
rect 13134 19014 13186 19066
rect 3424 18955 3476 18964
rect 3424 18921 3433 18955
rect 3433 18921 3467 18955
rect 3467 18921 3476 18955
rect 3424 18912 3476 18921
rect 3884 18955 3936 18964
rect 3884 18921 3893 18955
rect 3893 18921 3927 18955
rect 3927 18921 3936 18955
rect 3884 18912 3936 18921
rect 5816 18912 5868 18964
rect 9128 18955 9180 18964
rect 3608 18776 3660 18828
rect 7748 18844 7800 18896
rect 4436 18819 4488 18828
rect 4436 18785 4445 18819
rect 4445 18785 4479 18819
rect 4479 18785 4488 18819
rect 4436 18776 4488 18785
rect 4620 18708 4672 18760
rect 7288 18776 7340 18828
rect 7380 18708 7432 18760
rect 7932 18819 7984 18828
rect 7932 18785 7941 18819
rect 7941 18785 7975 18819
rect 7975 18785 7984 18819
rect 8576 18887 8628 18896
rect 8576 18853 8585 18887
rect 8585 18853 8619 18887
rect 8619 18853 8628 18887
rect 9128 18921 9137 18955
rect 9137 18921 9171 18955
rect 9171 18921 9180 18955
rect 9128 18912 9180 18921
rect 10600 18955 10652 18964
rect 10600 18921 10609 18955
rect 10609 18921 10643 18955
rect 10643 18921 10652 18955
rect 10600 18912 10652 18921
rect 11244 18955 11296 18964
rect 11244 18921 11253 18955
rect 11253 18921 11287 18955
rect 11287 18921 11296 18955
rect 11244 18912 11296 18921
rect 12348 18912 12400 18964
rect 13820 18955 13872 18964
rect 13820 18921 13829 18955
rect 13829 18921 13863 18955
rect 13863 18921 13872 18955
rect 13820 18912 13872 18921
rect 11520 18887 11572 18896
rect 8576 18844 8628 18853
rect 7932 18776 7984 18785
rect 9312 18819 9364 18828
rect 7564 18640 7616 18692
rect 4344 18615 4396 18624
rect 4344 18581 4353 18615
rect 4353 18581 4387 18615
rect 4387 18581 4396 18615
rect 4344 18572 4396 18581
rect 6736 18572 6788 18624
rect 8208 18640 8260 18692
rect 8300 18572 8352 18624
rect 9312 18785 9321 18819
rect 9321 18785 9355 18819
rect 9355 18785 9364 18819
rect 9312 18776 9364 18785
rect 11520 18853 11529 18887
rect 11529 18853 11563 18887
rect 11563 18853 11572 18887
rect 15660 18912 15712 18964
rect 11520 18844 11572 18853
rect 15476 18844 15528 18896
rect 17040 18844 17092 18896
rect 18144 18844 18196 18896
rect 11796 18819 11848 18828
rect 11796 18785 11819 18819
rect 11819 18785 11848 18819
rect 8576 18640 8628 18692
rect 9128 18640 9180 18692
rect 11796 18776 11848 18785
rect 12072 18819 12124 18828
rect 12072 18785 12081 18819
rect 12081 18785 12115 18819
rect 12115 18785 12124 18819
rect 12072 18776 12124 18785
rect 14280 18776 14332 18828
rect 18052 18776 18104 18828
rect 12716 18708 12768 18760
rect 13728 18708 13780 18760
rect 12348 18640 12400 18692
rect 12532 18640 12584 18692
rect 12624 18640 12676 18692
rect 16948 18708 17000 18760
rect 18696 18683 18748 18692
rect 18696 18649 18705 18683
rect 18705 18649 18739 18683
rect 18739 18649 18748 18683
rect 18696 18640 18748 18649
rect 8852 18615 8904 18624
rect 8852 18581 8861 18615
rect 8861 18581 8895 18615
rect 8895 18581 8904 18615
rect 8852 18572 8904 18581
rect 11704 18572 11756 18624
rect 13728 18572 13780 18624
rect 17224 18572 17276 18624
rect 18236 18572 18288 18624
rect 3972 18470 4024 18522
rect 4036 18470 4088 18522
rect 4100 18470 4152 18522
rect 4164 18470 4216 18522
rect 9952 18470 10004 18522
rect 10016 18470 10068 18522
rect 10080 18470 10132 18522
rect 10144 18470 10196 18522
rect 15932 18470 15984 18522
rect 15996 18470 16048 18522
rect 16060 18470 16112 18522
rect 16124 18470 16176 18522
rect 7748 18368 7800 18420
rect 12808 18411 12860 18420
rect 6736 18275 6788 18284
rect 6736 18241 6745 18275
rect 6745 18241 6779 18275
rect 6779 18241 6788 18275
rect 6736 18232 6788 18241
rect 12808 18377 12817 18411
rect 12817 18377 12851 18411
rect 12851 18377 12860 18411
rect 12808 18368 12860 18377
rect 11796 18300 11848 18352
rect 4620 18164 4672 18216
rect 4804 18164 4856 18216
rect 6460 18207 6512 18216
rect 6460 18173 6469 18207
rect 6469 18173 6503 18207
rect 6503 18173 6512 18207
rect 6460 18164 6512 18173
rect 8300 18207 8352 18216
rect 8300 18173 8309 18207
rect 8309 18173 8343 18207
rect 8343 18173 8352 18207
rect 8300 18164 8352 18173
rect 11520 18232 11572 18284
rect 9036 18207 9088 18216
rect 7288 18096 7340 18148
rect 8208 18096 8260 18148
rect 9036 18173 9045 18207
rect 9045 18173 9079 18207
rect 9079 18173 9088 18207
rect 9036 18164 9088 18173
rect 9128 18207 9180 18216
rect 9128 18173 9137 18207
rect 9137 18173 9171 18207
rect 9171 18173 9180 18207
rect 11704 18207 11756 18216
rect 9128 18164 9180 18173
rect 11704 18173 11713 18207
rect 11713 18173 11747 18207
rect 11747 18173 11756 18207
rect 11704 18164 11756 18173
rect 16948 18275 17000 18284
rect 12072 18207 12124 18216
rect 12072 18173 12081 18207
rect 12081 18173 12115 18207
rect 12115 18173 12124 18207
rect 12072 18164 12124 18173
rect 12716 18207 12768 18216
rect 12716 18173 12725 18207
rect 12725 18173 12759 18207
rect 12759 18173 12768 18207
rect 12716 18164 12768 18173
rect 16948 18241 16957 18275
rect 16957 18241 16991 18275
rect 16991 18241 17000 18275
rect 16948 18232 17000 18241
rect 17224 18275 17276 18284
rect 17224 18241 17233 18275
rect 17233 18241 17267 18275
rect 17267 18241 17276 18275
rect 17224 18232 17276 18241
rect 13452 18164 13504 18216
rect 12808 18139 12860 18148
rect 12808 18105 12817 18139
rect 12817 18105 12851 18139
rect 12851 18105 12860 18139
rect 12808 18096 12860 18105
rect 18236 18096 18288 18148
rect 4344 18028 4396 18080
rect 7748 18028 7800 18080
rect 9312 18028 9364 18080
rect 12256 18071 12308 18080
rect 12256 18037 12265 18071
rect 12265 18037 12299 18071
rect 12299 18037 12308 18071
rect 12256 18028 12308 18037
rect 6962 17926 7014 17978
rect 7026 17926 7078 17978
rect 7090 17926 7142 17978
rect 7154 17926 7206 17978
rect 12942 17926 12994 17978
rect 13006 17926 13058 17978
rect 13070 17926 13122 17978
rect 13134 17926 13186 17978
rect 7288 17824 7340 17876
rect 11796 17824 11848 17876
rect 12808 17824 12860 17876
rect 4436 17799 4488 17808
rect 4436 17765 4445 17799
rect 4445 17765 4479 17799
rect 4479 17765 4488 17799
rect 4436 17756 4488 17765
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 4620 17731 4672 17740
rect 4620 17697 4629 17731
rect 4629 17697 4663 17731
rect 4663 17697 4672 17731
rect 4620 17688 4672 17697
rect 3608 17552 3660 17604
rect 7380 17688 7432 17740
rect 7748 17688 7800 17740
rect 12532 17756 12584 17808
rect 13268 17756 13320 17808
rect 11520 17731 11572 17740
rect 11520 17697 11529 17731
rect 11529 17697 11563 17731
rect 11563 17697 11572 17731
rect 11520 17688 11572 17697
rect 11704 17731 11756 17740
rect 11704 17697 11713 17731
rect 11713 17697 11747 17731
rect 11747 17697 11756 17731
rect 11704 17688 11756 17697
rect 11888 17731 11940 17740
rect 11888 17697 11897 17731
rect 11897 17697 11931 17731
rect 11931 17697 11940 17731
rect 11888 17688 11940 17697
rect 12072 17731 12124 17740
rect 12072 17697 12081 17731
rect 12081 17697 12115 17731
rect 12115 17697 12124 17731
rect 12072 17688 12124 17697
rect 13176 17731 13228 17740
rect 13176 17697 13185 17731
rect 13185 17697 13219 17731
rect 13219 17697 13228 17731
rect 13176 17688 13228 17697
rect 12348 17663 12400 17672
rect 12348 17629 12357 17663
rect 12357 17629 12391 17663
rect 12391 17629 12400 17663
rect 12348 17620 12400 17629
rect 9680 17552 9732 17604
rect 12256 17552 12308 17604
rect 12716 17620 12768 17672
rect 13452 17731 13504 17740
rect 13452 17697 13461 17731
rect 13461 17697 13495 17731
rect 13495 17697 13504 17731
rect 14924 17756 14976 17808
rect 13452 17688 13504 17697
rect 14280 17688 14332 17740
rect 15016 17688 15068 17740
rect 1676 17484 1728 17536
rect 3792 17484 3844 17536
rect 4804 17527 4856 17536
rect 4804 17493 4813 17527
rect 4813 17493 4847 17527
rect 4847 17493 4856 17527
rect 4804 17484 4856 17493
rect 10324 17484 10376 17536
rect 11244 17484 11296 17536
rect 11704 17484 11756 17536
rect 12348 17484 12400 17536
rect 13360 17552 13412 17604
rect 14648 17620 14700 17672
rect 13544 17484 13596 17536
rect 13820 17484 13872 17536
rect 14832 17484 14884 17536
rect 3972 17382 4024 17434
rect 4036 17382 4088 17434
rect 4100 17382 4152 17434
rect 4164 17382 4216 17434
rect 9952 17382 10004 17434
rect 10016 17382 10068 17434
rect 10080 17382 10132 17434
rect 10144 17382 10196 17434
rect 15932 17382 15984 17434
rect 15996 17382 16048 17434
rect 16060 17382 16112 17434
rect 16124 17382 16176 17434
rect 4620 17280 4672 17332
rect 12072 17323 12124 17332
rect 4896 17187 4948 17196
rect 3608 17119 3660 17128
rect 3608 17085 3617 17119
rect 3617 17085 3651 17119
rect 3651 17085 3660 17119
rect 3608 17076 3660 17085
rect 3792 17076 3844 17128
rect 4528 17076 4580 17128
rect 4896 17153 4905 17187
rect 4905 17153 4939 17187
rect 4939 17153 4948 17187
rect 4896 17144 4948 17153
rect 9680 17187 9732 17196
rect 9680 17153 9689 17187
rect 9689 17153 9723 17187
rect 9723 17153 9732 17187
rect 9680 17144 9732 17153
rect 9772 17144 9824 17196
rect 11336 17212 11388 17264
rect 12072 17289 12081 17323
rect 12081 17289 12115 17323
rect 12115 17289 12124 17323
rect 12072 17280 12124 17289
rect 13084 17280 13136 17332
rect 13268 17280 13320 17332
rect 13452 17280 13504 17332
rect 14924 17212 14976 17264
rect 1860 17008 1912 17060
rect 4436 17008 4488 17060
rect 4712 17119 4764 17128
rect 4712 17085 4721 17119
rect 4721 17085 4755 17119
rect 4755 17085 4764 17119
rect 4988 17119 5040 17128
rect 4712 17076 4764 17085
rect 4988 17085 4997 17119
rect 4997 17085 5031 17119
rect 5031 17085 5040 17119
rect 4988 17076 5040 17085
rect 7748 17076 7800 17128
rect 9036 17076 9088 17128
rect 10600 17076 10652 17128
rect 11244 17076 11296 17128
rect 11336 17076 11388 17128
rect 16396 17144 16448 17196
rect 13084 17076 13136 17128
rect 13360 17076 13412 17128
rect 17224 17144 17276 17196
rect 8116 17008 8168 17060
rect 10048 17051 10100 17060
rect 10048 17017 10057 17051
rect 10057 17017 10091 17051
rect 10091 17017 10100 17051
rect 10048 17008 10100 17017
rect 10784 17008 10836 17060
rect 11704 17051 11756 17060
rect 11704 17017 11713 17051
rect 11713 17017 11747 17051
rect 11747 17017 11756 17051
rect 11704 17008 11756 17017
rect 12256 17008 12308 17060
rect 13728 17008 13780 17060
rect 13820 17051 13872 17060
rect 13820 17017 13829 17051
rect 13829 17017 13863 17051
rect 13863 17017 13872 17051
rect 13820 17008 13872 17017
rect 14832 17008 14884 17060
rect 4804 16940 4856 16992
rect 7564 16983 7616 16992
rect 7564 16949 7573 16983
rect 7573 16949 7607 16983
rect 7607 16949 7616 16983
rect 7564 16940 7616 16949
rect 9956 16940 10008 16992
rect 10692 16940 10744 16992
rect 16764 17076 16816 17128
rect 17040 17051 17092 17060
rect 17040 17017 17049 17051
rect 17049 17017 17083 17051
rect 17083 17017 17092 17051
rect 17040 17008 17092 17017
rect 16580 16940 16632 16992
rect 16672 16940 16724 16992
rect 17500 17076 17552 17128
rect 6962 16838 7014 16890
rect 7026 16838 7078 16890
rect 7090 16838 7142 16890
rect 7154 16838 7206 16890
rect 12942 16838 12994 16890
rect 13006 16838 13058 16890
rect 13070 16838 13122 16890
rect 13134 16838 13186 16890
rect 4712 16736 4764 16788
rect 16396 16779 16448 16788
rect 16396 16745 16405 16779
rect 16405 16745 16439 16779
rect 16439 16745 16448 16779
rect 16396 16736 16448 16745
rect 16580 16736 16632 16788
rect 7564 16668 7616 16720
rect 4804 16600 4856 16652
rect 4988 16643 5040 16652
rect 4988 16609 4997 16643
rect 4997 16609 5031 16643
rect 5031 16609 5040 16643
rect 4988 16600 5040 16609
rect 4896 16575 4948 16584
rect 4896 16541 4905 16575
rect 4905 16541 4939 16575
rect 4939 16541 4948 16575
rect 5908 16600 5960 16652
rect 9956 16643 10008 16652
rect 9956 16609 9965 16643
rect 9965 16609 9999 16643
rect 9999 16609 10008 16643
rect 9956 16600 10008 16609
rect 10232 16643 10284 16652
rect 10232 16609 10241 16643
rect 10241 16609 10275 16643
rect 10275 16609 10284 16643
rect 10232 16600 10284 16609
rect 10416 16643 10468 16652
rect 10416 16609 10425 16643
rect 10425 16609 10459 16643
rect 10459 16609 10468 16643
rect 10416 16600 10468 16609
rect 10600 16643 10652 16652
rect 10600 16609 10609 16643
rect 10609 16609 10643 16643
rect 10643 16609 10652 16643
rect 10600 16600 10652 16609
rect 10784 16643 10836 16652
rect 10784 16609 10793 16643
rect 10793 16609 10827 16643
rect 10827 16609 10836 16643
rect 10784 16600 10836 16609
rect 16672 16668 16724 16720
rect 16764 16643 16816 16652
rect 16764 16609 16773 16643
rect 16773 16609 16807 16643
rect 16807 16609 16816 16643
rect 16764 16600 16816 16609
rect 18512 16736 18564 16788
rect 17040 16600 17092 16652
rect 18052 16600 18104 16652
rect 6552 16575 6604 16584
rect 4896 16532 4948 16541
rect 6552 16541 6561 16575
rect 6561 16541 6595 16575
rect 6595 16541 6604 16575
rect 6552 16532 6604 16541
rect 6920 16532 6972 16584
rect 9404 16532 9456 16584
rect 17224 16532 17276 16584
rect 4804 16439 4856 16448
rect 4804 16405 4813 16439
rect 4813 16405 4847 16439
rect 4847 16405 4856 16439
rect 4804 16396 4856 16405
rect 8300 16439 8352 16448
rect 8300 16405 8309 16439
rect 8309 16405 8343 16439
rect 8343 16405 8352 16439
rect 8300 16396 8352 16405
rect 17960 16396 18012 16448
rect 3972 16294 4024 16346
rect 4036 16294 4088 16346
rect 4100 16294 4152 16346
rect 4164 16294 4216 16346
rect 9952 16294 10004 16346
rect 10016 16294 10068 16346
rect 10080 16294 10132 16346
rect 10144 16294 10196 16346
rect 15932 16294 15984 16346
rect 15996 16294 16048 16346
rect 16060 16294 16112 16346
rect 16124 16294 16176 16346
rect 6920 16235 6972 16244
rect 6920 16201 6929 16235
rect 6929 16201 6963 16235
rect 6963 16201 6972 16235
rect 6920 16192 6972 16201
rect 4528 16124 4580 16176
rect 3608 15988 3660 16040
rect 7472 16056 7524 16108
rect 8116 16124 8168 16176
rect 9680 16124 9732 16176
rect 10324 16124 10376 16176
rect 10600 16192 10652 16244
rect 7196 16031 7248 16040
rect 7196 15997 7205 16031
rect 7205 15997 7239 16031
rect 7239 15997 7248 16031
rect 7196 15988 7248 15997
rect 9588 15988 9640 16040
rect 4252 15920 4304 15972
rect 4436 15920 4488 15972
rect 5172 15920 5224 15972
rect 8300 15920 8352 15972
rect 9772 15920 9824 15972
rect 2872 15852 2924 15904
rect 13728 16124 13780 16176
rect 12808 16056 12860 16108
rect 10048 16031 10100 16040
rect 10048 15997 10057 16031
rect 10057 15997 10091 16031
rect 10091 15997 10100 16031
rect 10048 15988 10100 15997
rect 10324 16031 10376 16040
rect 10324 15997 10333 16031
rect 10333 15997 10367 16031
rect 10367 15997 10376 16031
rect 10324 15988 10376 15997
rect 11060 15988 11112 16040
rect 11980 15988 12032 16040
rect 13268 15988 13320 16040
rect 13544 15988 13596 16040
rect 14464 16031 14516 16040
rect 14464 15997 14473 16031
rect 14473 15997 14507 16031
rect 14507 15997 14516 16031
rect 14464 15988 14516 15997
rect 16396 16056 16448 16108
rect 12072 15963 12124 15972
rect 12072 15929 12081 15963
rect 12081 15929 12115 15963
rect 12115 15929 12124 15963
rect 12072 15920 12124 15929
rect 12164 15963 12216 15972
rect 12164 15929 12173 15963
rect 12173 15929 12207 15963
rect 12207 15929 12216 15963
rect 14556 15963 14608 15972
rect 12164 15920 12216 15929
rect 14556 15929 14565 15963
rect 14565 15929 14599 15963
rect 14599 15929 14608 15963
rect 14556 15920 14608 15929
rect 15016 16031 15068 16040
rect 15016 15997 15033 16031
rect 15033 15997 15067 16031
rect 15067 15997 15068 16031
rect 15016 15988 15068 15997
rect 16580 15920 16632 15972
rect 17132 15920 17184 15972
rect 17960 15920 18012 15972
rect 13452 15852 13504 15904
rect 14280 15895 14332 15904
rect 14280 15861 14289 15895
rect 14289 15861 14323 15895
rect 14323 15861 14332 15895
rect 14280 15852 14332 15861
rect 14832 15852 14884 15904
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 6962 15750 7014 15802
rect 7026 15750 7078 15802
rect 7090 15750 7142 15802
rect 7154 15750 7206 15802
rect 12942 15750 12994 15802
rect 13006 15750 13058 15802
rect 13070 15750 13122 15802
rect 13134 15750 13186 15802
rect 7472 15691 7524 15700
rect 7472 15657 7481 15691
rect 7481 15657 7515 15691
rect 7515 15657 7524 15691
rect 7472 15648 7524 15657
rect 10048 15648 10100 15700
rect 12164 15648 12216 15700
rect 13268 15648 13320 15700
rect 14924 15648 14976 15700
rect 16948 15648 17000 15700
rect 17132 15691 17184 15700
rect 17132 15657 17141 15691
rect 17141 15657 17175 15691
rect 17175 15657 17184 15691
rect 17132 15648 17184 15657
rect 17224 15691 17276 15700
rect 17224 15657 17233 15691
rect 17233 15657 17267 15691
rect 17267 15657 17276 15691
rect 17224 15648 17276 15657
rect 2872 15580 2924 15632
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 1860 15555 1912 15564
rect 1860 15521 1869 15555
rect 1869 15521 1903 15555
rect 1903 15521 1912 15555
rect 1860 15512 1912 15521
rect 4804 15623 4856 15632
rect 4804 15589 4813 15623
rect 4813 15589 4847 15623
rect 4847 15589 4856 15623
rect 4804 15580 4856 15589
rect 4252 15555 4304 15564
rect 4252 15521 4261 15555
rect 4261 15521 4295 15555
rect 4295 15521 4304 15555
rect 4252 15512 4304 15521
rect 4436 15512 4488 15564
rect 4528 15555 4580 15564
rect 4528 15521 4537 15555
rect 4537 15521 4571 15555
rect 4571 15521 4580 15555
rect 4988 15555 5040 15564
rect 4528 15512 4580 15521
rect 4988 15521 4997 15555
rect 4997 15521 5031 15555
rect 5031 15521 5040 15555
rect 4988 15512 5040 15521
rect 12716 15580 12768 15632
rect 13452 15623 13504 15632
rect 13452 15589 13461 15623
rect 13461 15589 13495 15623
rect 13495 15589 13504 15623
rect 13452 15580 13504 15589
rect 14280 15580 14332 15632
rect 15200 15580 15252 15632
rect 7472 15555 7524 15564
rect 7472 15521 7481 15555
rect 7481 15521 7515 15555
rect 7515 15521 7524 15555
rect 7472 15512 7524 15521
rect 7656 15555 7708 15564
rect 7656 15521 7665 15555
rect 7665 15521 7699 15555
rect 7699 15521 7708 15555
rect 7656 15512 7708 15521
rect 9588 15512 9640 15564
rect 12072 15512 12124 15564
rect 16580 15555 16632 15564
rect 16580 15521 16589 15555
rect 16589 15521 16623 15555
rect 16623 15521 16632 15555
rect 16580 15512 16632 15521
rect 16948 15555 17000 15564
rect 11888 15444 11940 15496
rect 13728 15487 13780 15496
rect 13728 15453 13737 15487
rect 13737 15453 13771 15487
rect 13771 15453 13780 15487
rect 13728 15444 13780 15453
rect 16948 15521 16957 15555
rect 16957 15521 16991 15555
rect 16991 15521 17000 15555
rect 16948 15512 17000 15521
rect 17224 15512 17276 15564
rect 17408 15555 17460 15564
rect 17408 15521 17417 15555
rect 17417 15521 17451 15555
rect 17451 15521 17460 15555
rect 17408 15512 17460 15521
rect 17592 15555 17644 15564
rect 17592 15521 17601 15555
rect 17601 15521 17635 15555
rect 17635 15521 17644 15555
rect 17592 15512 17644 15521
rect 17868 15512 17920 15564
rect 18696 15555 18748 15564
rect 18696 15521 18705 15555
rect 18705 15521 18739 15555
rect 18739 15521 18748 15555
rect 18696 15512 18748 15521
rect 4804 15376 4856 15428
rect 5356 15376 5408 15428
rect 1768 15308 1820 15360
rect 4436 15308 4488 15360
rect 5448 15308 5500 15360
rect 5724 15308 5776 15360
rect 11704 15308 11756 15360
rect 12440 15308 12492 15360
rect 12716 15308 12768 15360
rect 15016 15308 15068 15360
rect 15752 15308 15804 15360
rect 17868 15351 17920 15360
rect 17868 15317 17877 15351
rect 17877 15317 17911 15351
rect 17911 15317 17920 15351
rect 17868 15308 17920 15317
rect 17960 15308 18012 15360
rect 3972 15206 4024 15258
rect 4036 15206 4088 15258
rect 4100 15206 4152 15258
rect 4164 15206 4216 15258
rect 9952 15206 10004 15258
rect 10016 15206 10068 15258
rect 10080 15206 10132 15258
rect 10144 15206 10196 15258
rect 15932 15206 15984 15258
rect 15996 15206 16048 15258
rect 16060 15206 16112 15258
rect 16124 15206 16176 15258
rect 4988 15104 5040 15156
rect 5356 15147 5408 15156
rect 5356 15113 5365 15147
rect 5365 15113 5399 15147
rect 5399 15113 5408 15147
rect 5356 15104 5408 15113
rect 7656 15104 7708 15156
rect 9680 15147 9732 15156
rect 4712 14968 4764 15020
rect 5632 15036 5684 15088
rect 4436 14900 4488 14952
rect 7288 15036 7340 15088
rect 7564 15036 7616 15088
rect 5080 14900 5132 14952
rect 5448 14900 5500 14952
rect 5724 14943 5776 14952
rect 5724 14909 5733 14943
rect 5733 14909 5767 14943
rect 5767 14909 5776 14943
rect 5724 14900 5776 14909
rect 5908 14900 5960 14952
rect 7380 14900 7432 14952
rect 7932 14900 7984 14952
rect 8208 14900 8260 14952
rect 9680 15113 9689 15147
rect 9689 15113 9723 15147
rect 9723 15113 9732 15147
rect 9680 15104 9732 15113
rect 10416 15147 10468 15156
rect 10416 15113 10425 15147
rect 10425 15113 10459 15147
rect 10459 15113 10468 15147
rect 10416 15104 10468 15113
rect 8116 14875 8168 14884
rect 5264 14764 5316 14816
rect 7288 14764 7340 14816
rect 8116 14841 8125 14875
rect 8125 14841 8159 14875
rect 8159 14841 8168 14875
rect 8116 14832 8168 14841
rect 10968 14900 11020 14952
rect 11888 14943 11940 14952
rect 11888 14909 11897 14943
rect 11897 14909 11931 14943
rect 11931 14909 11940 14943
rect 11888 14900 11940 14909
rect 12164 14943 12216 14952
rect 12164 14909 12173 14943
rect 12173 14909 12207 14943
rect 12207 14909 12216 14943
rect 12164 14900 12216 14909
rect 10324 14832 10376 14884
rect 12072 14875 12124 14884
rect 12072 14841 12081 14875
rect 12081 14841 12115 14875
rect 12115 14841 12124 14875
rect 14832 15036 14884 15088
rect 14556 14900 14608 14952
rect 14832 14900 14884 14952
rect 16396 14900 16448 14952
rect 17592 14968 17644 15020
rect 17868 14900 17920 14952
rect 12072 14832 12124 14841
rect 17408 14832 17460 14884
rect 17592 14832 17644 14884
rect 8300 14764 8352 14816
rect 11520 14764 11572 14816
rect 14648 14807 14700 14816
rect 14648 14773 14657 14807
rect 14657 14773 14691 14807
rect 14691 14773 14700 14807
rect 14648 14764 14700 14773
rect 14740 14764 14792 14816
rect 14924 14764 14976 14816
rect 6962 14662 7014 14714
rect 7026 14662 7078 14714
rect 7090 14662 7142 14714
rect 7154 14662 7206 14714
rect 12942 14662 12994 14714
rect 13006 14662 13058 14714
rect 13070 14662 13122 14714
rect 13134 14662 13186 14714
rect 7472 14560 7524 14612
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 2596 14424 2648 14476
rect 4988 14424 5040 14476
rect 5908 14492 5960 14544
rect 5448 14467 5500 14476
rect 4804 14399 4856 14408
rect 4804 14365 4813 14399
rect 4813 14365 4847 14399
rect 4847 14365 4856 14399
rect 4804 14356 4856 14365
rect 5448 14433 5457 14467
rect 5457 14433 5491 14467
rect 5491 14433 5500 14467
rect 5448 14424 5500 14433
rect 5724 14424 5776 14476
rect 7012 14467 7064 14476
rect 7012 14433 7021 14467
rect 7021 14433 7055 14467
rect 7055 14433 7064 14467
rect 7012 14424 7064 14433
rect 7196 14424 7248 14476
rect 6184 14356 6236 14408
rect 7564 14356 7616 14408
rect 5448 14288 5500 14340
rect 7380 14288 7432 14340
rect 7840 14399 7892 14408
rect 7840 14365 7849 14399
rect 7849 14365 7883 14399
rect 7883 14365 7892 14399
rect 7840 14356 7892 14365
rect 8116 14560 8168 14612
rect 10968 14603 11020 14612
rect 10968 14569 10977 14603
rect 10977 14569 11011 14603
rect 11011 14569 11020 14603
rect 10968 14560 11020 14569
rect 11520 14560 11572 14612
rect 16764 14560 16816 14612
rect 8208 14424 8260 14476
rect 11520 14399 11572 14408
rect 11520 14365 11529 14399
rect 11529 14365 11563 14399
rect 11563 14365 11572 14399
rect 11520 14356 11572 14365
rect 12532 14356 12584 14408
rect 17592 14424 17644 14476
rect 17776 14356 17828 14408
rect 8024 14331 8076 14340
rect 8024 14297 8033 14331
rect 8033 14297 8067 14331
rect 8067 14297 8076 14331
rect 8024 14288 8076 14297
rect 2504 14220 2556 14272
rect 4896 14263 4948 14272
rect 4896 14229 4905 14263
rect 4905 14229 4939 14263
rect 4939 14229 4948 14263
rect 4896 14220 4948 14229
rect 5724 14220 5776 14272
rect 7472 14263 7524 14272
rect 7472 14229 7481 14263
rect 7481 14229 7515 14263
rect 7515 14229 7524 14263
rect 7472 14220 7524 14229
rect 7656 14220 7708 14272
rect 9404 14288 9456 14340
rect 9220 14220 9272 14272
rect 3972 14118 4024 14170
rect 4036 14118 4088 14170
rect 4100 14118 4152 14170
rect 4164 14118 4216 14170
rect 9952 14118 10004 14170
rect 10016 14118 10068 14170
rect 10080 14118 10132 14170
rect 10144 14118 10196 14170
rect 15932 14118 15984 14170
rect 15996 14118 16048 14170
rect 16060 14118 16112 14170
rect 16124 14118 16176 14170
rect 7012 14016 7064 14068
rect 7288 14016 7340 14068
rect 11060 14016 11112 14068
rect 14648 14016 14700 14068
rect 15660 14016 15712 14068
rect 16396 14059 16448 14068
rect 16396 14025 16405 14059
rect 16405 14025 16439 14059
rect 16439 14025 16448 14059
rect 16396 14016 16448 14025
rect 18512 14059 18564 14068
rect 18512 14025 18521 14059
rect 18521 14025 18555 14059
rect 18555 14025 18564 14059
rect 18512 14016 18564 14025
rect 4528 13880 4580 13932
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 1492 13812 1544 13864
rect 2504 13855 2556 13864
rect 2504 13821 2513 13855
rect 2513 13821 2547 13855
rect 2547 13821 2556 13855
rect 2504 13812 2556 13821
rect 4896 13855 4948 13864
rect 4896 13821 4900 13855
rect 4900 13821 4934 13855
rect 4934 13821 4948 13855
rect 4896 13812 4948 13821
rect 5448 13855 5500 13864
rect 5448 13821 5449 13855
rect 5449 13821 5483 13855
rect 5483 13821 5500 13855
rect 5724 13855 5776 13864
rect 1584 13719 1636 13728
rect 1584 13685 1593 13719
rect 1593 13685 1627 13719
rect 1627 13685 1636 13719
rect 1584 13676 1636 13685
rect 3056 13719 3108 13728
rect 3056 13685 3065 13719
rect 3065 13685 3099 13719
rect 3099 13685 3108 13719
rect 3056 13676 3108 13685
rect 4804 13676 4856 13728
rect 5080 13787 5132 13796
rect 5080 13753 5089 13787
rect 5089 13753 5123 13787
rect 5123 13753 5132 13787
rect 5448 13812 5500 13821
rect 5724 13821 5733 13855
rect 5733 13821 5767 13855
rect 5767 13821 5776 13855
rect 5724 13812 5776 13821
rect 7196 13855 7248 13864
rect 7196 13821 7200 13855
rect 7200 13821 7234 13855
rect 7234 13821 7248 13855
rect 7196 13812 7248 13821
rect 7472 13855 7524 13864
rect 7472 13821 7517 13855
rect 7517 13821 7524 13855
rect 7472 13812 7524 13821
rect 5080 13744 5132 13753
rect 6828 13676 6880 13728
rect 7380 13787 7432 13796
rect 7380 13753 7389 13787
rect 7389 13753 7423 13787
rect 7423 13753 7432 13787
rect 8024 13812 8076 13864
rect 9220 13855 9272 13864
rect 9220 13821 9229 13855
rect 9229 13821 9263 13855
rect 9263 13821 9272 13855
rect 9220 13812 9272 13821
rect 9496 13812 9548 13864
rect 9864 13812 9916 13864
rect 13268 13880 13320 13932
rect 15844 13880 15896 13932
rect 15292 13855 15344 13864
rect 7380 13744 7432 13753
rect 9588 13719 9640 13728
rect 9588 13685 9597 13719
rect 9597 13685 9631 13719
rect 9631 13685 9640 13719
rect 9588 13676 9640 13685
rect 13452 13719 13504 13728
rect 13452 13685 13461 13719
rect 13461 13685 13495 13719
rect 13495 13685 13504 13719
rect 13452 13676 13504 13685
rect 15016 13676 15068 13728
rect 15292 13821 15301 13855
rect 15301 13821 15335 13855
rect 15335 13821 15344 13855
rect 15292 13812 15344 13821
rect 15476 13855 15528 13864
rect 15476 13821 15485 13855
rect 15485 13821 15519 13855
rect 15519 13821 15528 13855
rect 15476 13812 15528 13821
rect 15752 13812 15804 13864
rect 17408 13855 17460 13864
rect 17408 13821 17417 13855
rect 17417 13821 17451 13855
rect 17451 13821 17460 13855
rect 17408 13812 17460 13821
rect 17592 13855 17644 13864
rect 17592 13821 17601 13855
rect 17601 13821 17635 13855
rect 17635 13821 17644 13855
rect 17592 13812 17644 13821
rect 17776 13855 17828 13864
rect 17776 13821 17785 13855
rect 17785 13821 17819 13855
rect 17819 13821 17828 13855
rect 17776 13812 17828 13821
rect 18696 13855 18748 13864
rect 18696 13821 18705 13855
rect 18705 13821 18739 13855
rect 18739 13821 18748 13855
rect 18696 13812 18748 13821
rect 17500 13787 17552 13796
rect 17500 13753 17509 13787
rect 17509 13753 17543 13787
rect 17543 13753 17552 13787
rect 17500 13744 17552 13753
rect 6962 13574 7014 13626
rect 7026 13574 7078 13626
rect 7090 13574 7142 13626
rect 7154 13574 7206 13626
rect 12942 13574 12994 13626
rect 13006 13574 13058 13626
rect 13070 13574 13122 13626
rect 13134 13574 13186 13626
rect 1492 13515 1544 13524
rect 1492 13481 1501 13515
rect 1501 13481 1535 13515
rect 1535 13481 1544 13515
rect 1492 13472 1544 13481
rect 1952 13515 2004 13524
rect 1952 13481 1961 13515
rect 1961 13481 1995 13515
rect 1995 13481 2004 13515
rect 1952 13472 2004 13481
rect 3056 13472 3108 13524
rect 5080 13472 5132 13524
rect 5448 13472 5500 13524
rect 9680 13515 9732 13524
rect 9680 13481 9689 13515
rect 9689 13481 9723 13515
rect 9723 13481 9732 13515
rect 9680 13472 9732 13481
rect 12532 13515 12584 13524
rect 12532 13481 12541 13515
rect 12541 13481 12575 13515
rect 12575 13481 12584 13515
rect 12532 13472 12584 13481
rect 12808 13472 12860 13524
rect 2596 13379 2648 13388
rect 2596 13345 2605 13379
rect 2605 13345 2639 13379
rect 2639 13345 2648 13379
rect 2596 13336 2648 13345
rect 2872 13336 2924 13388
rect 11428 13404 11480 13456
rect 9128 13379 9180 13388
rect 2044 13311 2096 13320
rect 2044 13277 2053 13311
rect 2053 13277 2087 13311
rect 2087 13277 2096 13311
rect 2044 13268 2096 13277
rect 9128 13345 9137 13379
rect 9137 13345 9171 13379
rect 9171 13345 9180 13379
rect 9128 13336 9180 13345
rect 9404 13379 9456 13388
rect 9404 13345 9413 13379
rect 9413 13345 9447 13379
rect 9447 13345 9456 13379
rect 9404 13336 9456 13345
rect 9496 13379 9548 13388
rect 9496 13345 9505 13379
rect 9505 13345 9539 13379
rect 9539 13345 9548 13379
rect 9496 13336 9548 13345
rect 13820 13379 13872 13388
rect 3240 13311 3292 13320
rect 3240 13277 3249 13311
rect 3249 13277 3283 13311
rect 3283 13277 3292 13311
rect 3240 13268 3292 13277
rect 7932 13268 7984 13320
rect 9588 13268 9640 13320
rect 10416 13268 10468 13320
rect 12808 13268 12860 13320
rect 13820 13345 13829 13379
rect 13829 13345 13863 13379
rect 13863 13345 13872 13379
rect 13820 13336 13872 13345
rect 15292 13472 15344 13524
rect 15384 13472 15436 13524
rect 17408 13472 17460 13524
rect 18052 13472 18104 13524
rect 14832 13379 14884 13388
rect 14832 13345 14841 13379
rect 14841 13345 14875 13379
rect 14875 13345 14884 13379
rect 14832 13336 14884 13345
rect 15016 13379 15068 13388
rect 15016 13345 15025 13379
rect 15025 13345 15059 13379
rect 15059 13345 15068 13379
rect 15016 13336 15068 13345
rect 4896 13200 4948 13252
rect 5172 13200 5224 13252
rect 7196 13200 7248 13252
rect 13452 13200 13504 13252
rect 14740 13268 14792 13320
rect 15752 13379 15804 13388
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 15844 13379 15896 13388
rect 15844 13345 15853 13379
rect 15853 13345 15887 13379
rect 15887 13345 15896 13379
rect 15844 13336 15896 13345
rect 17132 13336 17184 13388
rect 17500 13336 17552 13388
rect 15384 13268 15436 13320
rect 15660 13268 15712 13320
rect 15476 13200 15528 13252
rect 4528 13132 4580 13184
rect 11888 13175 11940 13184
rect 11888 13141 11897 13175
rect 11897 13141 11931 13175
rect 11931 13141 11940 13175
rect 11888 13132 11940 13141
rect 13268 13175 13320 13184
rect 13268 13141 13277 13175
rect 13277 13141 13311 13175
rect 13311 13141 13320 13175
rect 13268 13132 13320 13141
rect 17776 13200 17828 13252
rect 16396 13132 16448 13184
rect 18052 13175 18104 13184
rect 18052 13141 18061 13175
rect 18061 13141 18095 13175
rect 18095 13141 18104 13175
rect 18052 13132 18104 13141
rect 3972 13030 4024 13082
rect 4036 13030 4088 13082
rect 4100 13030 4152 13082
rect 4164 13030 4216 13082
rect 9952 13030 10004 13082
rect 10016 13030 10068 13082
rect 10080 13030 10132 13082
rect 10144 13030 10196 13082
rect 15932 13030 15984 13082
rect 15996 13030 16048 13082
rect 16060 13030 16112 13082
rect 16124 13030 16176 13082
rect 3240 12928 3292 12980
rect 11428 12928 11480 12980
rect 15476 12928 15528 12980
rect 4896 12860 4948 12912
rect 5080 12860 5132 12912
rect 5632 12903 5684 12912
rect 5632 12869 5641 12903
rect 5641 12869 5675 12903
rect 5675 12869 5684 12903
rect 5632 12860 5684 12869
rect 7196 12903 7248 12912
rect 7196 12869 7205 12903
rect 7205 12869 7239 12903
rect 7239 12869 7248 12903
rect 7196 12860 7248 12869
rect 7380 12860 7432 12912
rect 7656 12860 7708 12912
rect 7932 12903 7984 12912
rect 4804 12835 4856 12844
rect 4804 12801 4813 12835
rect 4813 12801 4847 12835
rect 4847 12801 4856 12835
rect 4804 12792 4856 12801
rect 5356 12767 5408 12776
rect 5356 12733 5365 12767
rect 5365 12733 5399 12767
rect 5399 12733 5408 12767
rect 5356 12724 5408 12733
rect 5908 12792 5960 12844
rect 6920 12792 6972 12844
rect 6276 12724 6328 12776
rect 7564 12724 7616 12776
rect 7932 12869 7941 12903
rect 7941 12869 7975 12903
rect 7975 12869 7984 12903
rect 7932 12860 7984 12869
rect 9772 12792 9824 12844
rect 8208 12724 8260 12776
rect 11060 12724 11112 12776
rect 12624 12792 12676 12844
rect 14740 12792 14792 12844
rect 13820 12724 13872 12776
rect 16580 12724 16632 12776
rect 17132 12767 17184 12776
rect 17132 12733 17141 12767
rect 17141 12733 17175 12767
rect 17175 12733 17184 12767
rect 17132 12724 17184 12733
rect 11244 12656 11296 12708
rect 11980 12656 12032 12708
rect 13268 12656 13320 12708
rect 18052 12656 18104 12708
rect 4160 12588 4212 12640
rect 6828 12588 6880 12640
rect 10508 12588 10560 12640
rect 17500 12631 17552 12640
rect 17500 12597 17509 12631
rect 17509 12597 17543 12631
rect 17543 12597 17552 12631
rect 17500 12588 17552 12597
rect 6962 12486 7014 12538
rect 7026 12486 7078 12538
rect 7090 12486 7142 12538
rect 7154 12486 7206 12538
rect 12942 12486 12994 12538
rect 13006 12486 13058 12538
rect 13070 12486 13122 12538
rect 13134 12486 13186 12538
rect 1492 12087 1544 12096
rect 1492 12053 1501 12087
rect 1501 12053 1535 12087
rect 1535 12053 1544 12087
rect 1492 12044 1544 12053
rect 4160 12384 4212 12436
rect 5356 12384 5408 12436
rect 6276 12427 6328 12436
rect 2872 12359 2924 12368
rect 2872 12325 2881 12359
rect 2881 12325 2915 12359
rect 2915 12325 2924 12359
rect 2872 12316 2924 12325
rect 5080 12316 5132 12368
rect 6276 12393 6285 12427
rect 6285 12393 6319 12427
rect 6319 12393 6328 12427
rect 6276 12384 6328 12393
rect 16304 12384 16356 12436
rect 2964 12248 3016 12300
rect 11060 12316 11112 12368
rect 5540 12180 5592 12232
rect 7012 12248 7064 12300
rect 7748 12248 7800 12300
rect 9128 12248 9180 12300
rect 11152 12248 11204 12300
rect 11888 12248 11940 12300
rect 9312 12180 9364 12232
rect 13820 12316 13872 12368
rect 14188 12316 14240 12368
rect 12624 12248 12676 12300
rect 12808 12291 12860 12300
rect 12808 12257 12817 12291
rect 12817 12257 12851 12291
rect 12851 12257 12860 12291
rect 12808 12248 12860 12257
rect 13268 12248 13320 12300
rect 16856 12248 16908 12300
rect 18052 12384 18104 12436
rect 17500 12316 17552 12368
rect 18236 12316 18288 12368
rect 12716 12112 12768 12164
rect 4896 12044 4948 12096
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 9496 12044 9548 12096
rect 12624 12044 12676 12096
rect 13636 12044 13688 12096
rect 14924 12044 14976 12096
rect 3972 11942 4024 11994
rect 4036 11942 4088 11994
rect 4100 11942 4152 11994
rect 4164 11942 4216 11994
rect 9952 11942 10004 11994
rect 10016 11942 10068 11994
rect 10080 11942 10132 11994
rect 10144 11942 10196 11994
rect 15932 11942 15984 11994
rect 15996 11942 16048 11994
rect 16060 11942 16112 11994
rect 16124 11942 16176 11994
rect 2964 11883 3016 11892
rect 2964 11849 2973 11883
rect 2973 11849 3007 11883
rect 3007 11849 3016 11883
rect 2964 11840 3016 11849
rect 4528 11883 4580 11892
rect 4528 11849 4537 11883
rect 4537 11849 4571 11883
rect 4571 11849 4580 11883
rect 4528 11840 4580 11849
rect 5080 11840 5132 11892
rect 5540 11840 5592 11892
rect 6552 11840 6604 11892
rect 2044 11772 2096 11824
rect 1768 11747 1820 11756
rect 1768 11713 1777 11747
rect 1777 11713 1811 11747
rect 1811 11713 1820 11747
rect 1768 11704 1820 11713
rect 5080 11704 5132 11756
rect 2872 11679 2924 11688
rect 2872 11645 2881 11679
rect 2881 11645 2915 11679
rect 2915 11645 2924 11679
rect 2872 11636 2924 11645
rect 2964 11679 3016 11688
rect 2964 11645 2973 11679
rect 2973 11645 3007 11679
rect 3007 11645 3016 11679
rect 2964 11636 3016 11645
rect 5448 11704 5500 11756
rect 7472 11840 7524 11892
rect 9772 11840 9824 11892
rect 12808 11840 12860 11892
rect 18236 11840 18288 11892
rect 9496 11772 9548 11824
rect 6920 11747 6972 11756
rect 6920 11713 6929 11747
rect 6929 11713 6963 11747
rect 6963 11713 6972 11747
rect 6920 11704 6972 11713
rect 8300 11704 8352 11756
rect 12624 11747 12676 11756
rect 4160 11568 4212 11620
rect 4804 11568 4856 11620
rect 6368 11568 6420 11620
rect 8208 11636 8260 11688
rect 8668 11636 8720 11688
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12624 11704 12676 11713
rect 14188 11747 14240 11756
rect 14188 11713 14197 11747
rect 14197 11713 14231 11747
rect 14231 11713 14240 11747
rect 14188 11704 14240 11713
rect 15292 11704 15344 11756
rect 9404 11636 9456 11688
rect 7012 11568 7064 11620
rect 7656 11568 7708 11620
rect 4712 11500 4764 11552
rect 8484 11500 8536 11552
rect 9312 11568 9364 11620
rect 9772 11636 9824 11688
rect 10416 11568 10468 11620
rect 12532 11568 12584 11620
rect 13636 11568 13688 11620
rect 14924 11568 14976 11620
rect 16028 11568 16080 11620
rect 16304 11636 16356 11688
rect 16856 11636 16908 11688
rect 18696 11679 18748 11688
rect 18696 11645 18705 11679
rect 18705 11645 18739 11679
rect 18739 11645 18748 11679
rect 18696 11636 18748 11645
rect 17132 11500 17184 11552
rect 6962 11398 7014 11450
rect 7026 11398 7078 11450
rect 7090 11398 7142 11450
rect 7154 11398 7206 11450
rect 12942 11398 12994 11450
rect 13006 11398 13058 11450
rect 13070 11398 13122 11450
rect 13134 11398 13186 11450
rect 2964 11296 3016 11348
rect 4160 11339 4212 11348
rect 4160 11305 4169 11339
rect 4169 11305 4203 11339
rect 4203 11305 4212 11339
rect 4160 11296 4212 11305
rect 4988 11296 5040 11348
rect 8208 11339 8260 11348
rect 3700 11228 3752 11280
rect 8208 11305 8217 11339
rect 8217 11305 8251 11339
rect 8251 11305 8260 11339
rect 8208 11296 8260 11305
rect 12532 11296 12584 11348
rect 13728 11296 13780 11348
rect 17316 11296 17368 11348
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 2780 11160 2832 11169
rect 4620 11160 4672 11212
rect 5172 11160 5224 11212
rect 6276 11271 6328 11280
rect 6276 11237 6285 11271
rect 6285 11237 6319 11271
rect 6319 11237 6328 11271
rect 6276 11228 6328 11237
rect 16396 11271 16448 11280
rect 16396 11237 16405 11271
rect 16405 11237 16439 11271
rect 16439 11237 16448 11271
rect 16396 11228 16448 11237
rect 17132 11228 17184 11280
rect 5448 11092 5500 11144
rect 6368 11092 6420 11144
rect 7564 11092 7616 11144
rect 8484 11160 8536 11212
rect 9220 11160 9272 11212
rect 8944 11092 8996 11144
rect 11428 11203 11480 11212
rect 9680 11092 9732 11144
rect 11428 11169 11437 11203
rect 11437 11169 11471 11203
rect 11471 11169 11480 11203
rect 11428 11160 11480 11169
rect 13728 11160 13780 11212
rect 16028 11160 16080 11212
rect 11336 11092 11388 11144
rect 8484 11024 8536 11076
rect 11060 11024 11112 11076
rect 12624 11024 12676 11076
rect 5356 10956 5408 11008
rect 10324 10956 10376 11008
rect 15476 10956 15528 11008
rect 3972 10854 4024 10906
rect 4036 10854 4088 10906
rect 4100 10854 4152 10906
rect 4164 10854 4216 10906
rect 9952 10854 10004 10906
rect 10016 10854 10068 10906
rect 10080 10854 10132 10906
rect 10144 10854 10196 10906
rect 15932 10854 15984 10906
rect 15996 10854 16048 10906
rect 16060 10854 16112 10906
rect 16124 10854 16176 10906
rect 4804 10752 4856 10804
rect 6184 10795 6236 10804
rect 6184 10761 6193 10795
rect 6193 10761 6227 10795
rect 6227 10761 6236 10795
rect 6184 10752 6236 10761
rect 7288 10795 7340 10804
rect 4620 10684 4672 10736
rect 7288 10761 7297 10795
rect 7297 10761 7331 10795
rect 7331 10761 7340 10795
rect 7288 10752 7340 10761
rect 9680 10752 9732 10804
rect 10324 10752 10376 10804
rect 11428 10752 11480 10804
rect 4804 10616 4856 10668
rect 9404 10659 9456 10668
rect 5172 10548 5224 10600
rect 6368 10548 6420 10600
rect 6736 10548 6788 10600
rect 5080 10480 5132 10532
rect 7840 10548 7892 10600
rect 8300 10591 8352 10600
rect 8024 10480 8076 10532
rect 8300 10557 8309 10591
rect 8309 10557 8343 10591
rect 8343 10557 8352 10591
rect 8300 10548 8352 10557
rect 8484 10591 8536 10600
rect 8484 10557 8493 10591
rect 8493 10557 8527 10591
rect 8527 10557 8536 10591
rect 8484 10548 8536 10557
rect 8668 10591 8720 10600
rect 8668 10557 8677 10591
rect 8677 10557 8711 10591
rect 8711 10557 8720 10591
rect 8668 10548 8720 10557
rect 8944 10548 8996 10600
rect 9404 10625 9413 10659
rect 9413 10625 9447 10659
rect 9447 10625 9456 10659
rect 9404 10616 9456 10625
rect 9496 10591 9548 10600
rect 9496 10557 9505 10591
rect 9505 10557 9539 10591
rect 9539 10557 9548 10591
rect 9496 10548 9548 10557
rect 9772 10548 9824 10600
rect 11152 10684 11204 10736
rect 11060 10659 11112 10668
rect 11060 10625 11069 10659
rect 11069 10625 11103 10659
rect 11103 10625 11112 10659
rect 14372 10684 14424 10736
rect 11060 10616 11112 10625
rect 13636 10659 13688 10668
rect 13636 10625 13645 10659
rect 13645 10625 13679 10659
rect 13679 10625 13688 10659
rect 13636 10616 13688 10625
rect 12716 10548 12768 10600
rect 15108 10548 15160 10600
rect 15384 10591 15436 10600
rect 15384 10557 15393 10591
rect 15393 10557 15427 10591
rect 15427 10557 15436 10591
rect 15384 10548 15436 10557
rect 5356 10412 5408 10464
rect 8208 10412 8260 10464
rect 10600 10455 10652 10464
rect 10600 10421 10609 10455
rect 10609 10421 10643 10455
rect 10643 10421 10652 10455
rect 10600 10412 10652 10421
rect 11152 10412 11204 10464
rect 12348 10412 12400 10464
rect 18512 10480 18564 10532
rect 13268 10412 13320 10464
rect 15752 10412 15804 10464
rect 6962 10310 7014 10362
rect 7026 10310 7078 10362
rect 7090 10310 7142 10362
rect 7154 10310 7206 10362
rect 12942 10310 12994 10362
rect 13006 10310 13058 10362
rect 13070 10310 13122 10362
rect 13134 10310 13186 10362
rect 2780 10208 2832 10260
rect 4712 10251 4764 10260
rect 4712 10217 4721 10251
rect 4721 10217 4755 10251
rect 4755 10217 4764 10251
rect 4712 10208 4764 10217
rect 6552 10208 6604 10260
rect 12716 10208 12768 10260
rect 2964 10072 3016 10124
rect 3516 10115 3568 10124
rect 3516 10081 3525 10115
rect 3525 10081 3559 10115
rect 3559 10081 3568 10115
rect 3516 10072 3568 10081
rect 8208 10140 8260 10192
rect 4528 10072 4580 10124
rect 4988 10072 5040 10124
rect 6184 10072 6236 10124
rect 7288 10072 7340 10124
rect 9220 10115 9272 10124
rect 9220 10081 9229 10115
rect 9229 10081 9263 10115
rect 9263 10081 9272 10115
rect 9220 10072 9272 10081
rect 2780 9979 2832 9988
rect 2780 9945 2789 9979
rect 2789 9945 2823 9979
rect 2823 9945 2832 9979
rect 2780 9936 2832 9945
rect 5080 10004 5132 10056
rect 5356 10047 5408 10056
rect 5356 10013 5365 10047
rect 5365 10013 5399 10047
rect 5399 10013 5408 10047
rect 5356 10004 5408 10013
rect 7656 10004 7708 10056
rect 8300 10004 8352 10056
rect 9496 10072 9548 10124
rect 9680 10072 9732 10124
rect 10600 10140 10652 10192
rect 13544 10208 13596 10260
rect 15108 10251 15160 10260
rect 15108 10217 15117 10251
rect 15117 10217 15151 10251
rect 15151 10217 15160 10251
rect 15108 10208 15160 10217
rect 15476 10251 15528 10260
rect 15476 10217 15485 10251
rect 15485 10217 15519 10251
rect 15519 10217 15528 10251
rect 15476 10208 15528 10217
rect 16580 10208 16632 10260
rect 17960 10208 18012 10260
rect 12348 10072 12400 10124
rect 13636 10072 13688 10124
rect 14556 10072 14608 10124
rect 15108 10072 15160 10124
rect 9588 10004 9640 10056
rect 11428 10047 11480 10056
rect 11428 10013 11437 10047
rect 11437 10013 11471 10047
rect 11471 10013 11480 10047
rect 11428 10004 11480 10013
rect 4436 9868 4488 9920
rect 5172 9868 5224 9920
rect 6644 9911 6696 9920
rect 6644 9877 6653 9911
rect 6653 9877 6687 9911
rect 6687 9877 6696 9911
rect 6644 9868 6696 9877
rect 12808 9868 12860 9920
rect 15752 9868 15804 9920
rect 17500 9911 17552 9920
rect 17500 9877 17509 9911
rect 17509 9877 17543 9911
rect 17543 9877 17552 9911
rect 17500 9868 17552 9877
rect 3972 9766 4024 9818
rect 4036 9766 4088 9818
rect 4100 9766 4152 9818
rect 4164 9766 4216 9818
rect 9952 9766 10004 9818
rect 10016 9766 10068 9818
rect 10080 9766 10132 9818
rect 10144 9766 10196 9818
rect 15932 9766 15984 9818
rect 15996 9766 16048 9818
rect 16060 9766 16112 9818
rect 16124 9766 16176 9818
rect 4620 9664 4672 9716
rect 8944 9664 8996 9716
rect 15384 9664 15436 9716
rect 4528 9596 4580 9648
rect 2044 9528 2096 9580
rect 5264 9596 5316 9648
rect 6276 9596 6328 9648
rect 7288 9596 7340 9648
rect 7656 9639 7708 9648
rect 5080 9528 5132 9580
rect 6644 9528 6696 9580
rect 7656 9605 7665 9639
rect 7665 9605 7699 9639
rect 7699 9605 7708 9639
rect 7656 9596 7708 9605
rect 18512 9639 18564 9648
rect 18512 9605 18521 9639
rect 18521 9605 18555 9639
rect 18555 9605 18564 9639
rect 18512 9596 18564 9605
rect 8300 9528 8352 9580
rect 4896 9503 4948 9512
rect 1584 9392 1636 9444
rect 1860 9367 1912 9376
rect 1860 9333 1869 9367
rect 1869 9333 1903 9367
rect 1903 9333 1912 9367
rect 1860 9324 1912 9333
rect 2320 9324 2372 9376
rect 4344 9324 4396 9376
rect 4896 9469 4905 9503
rect 4905 9469 4939 9503
rect 4939 9469 4948 9503
rect 4896 9460 4948 9469
rect 4988 9392 5040 9444
rect 5356 9392 5408 9444
rect 6736 9392 6788 9444
rect 14556 9460 14608 9512
rect 15752 9503 15804 9512
rect 15752 9469 15761 9503
rect 15761 9469 15795 9503
rect 15795 9469 15804 9503
rect 18696 9503 18748 9512
rect 15752 9460 15804 9469
rect 18696 9469 18705 9503
rect 18705 9469 18739 9503
rect 18739 9469 18748 9503
rect 18696 9460 18748 9469
rect 15476 9392 15528 9444
rect 6828 9324 6880 9376
rect 6962 9222 7014 9274
rect 7026 9222 7078 9274
rect 7090 9222 7142 9274
rect 7154 9222 7206 9274
rect 12942 9222 12994 9274
rect 13006 9222 13058 9274
rect 13070 9222 13122 9274
rect 13134 9222 13186 9274
rect 1860 9120 1912 9172
rect 2504 9052 2556 9104
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 4896 9120 4948 9172
rect 5356 9120 5408 9172
rect 9128 9120 9180 9172
rect 4528 9052 4580 9104
rect 4712 9052 4764 9104
rect 11612 9120 11664 9172
rect 14556 9163 14608 9172
rect 5264 9027 5316 9036
rect 5264 8993 5273 9027
rect 5273 8993 5307 9027
rect 5307 8993 5316 9027
rect 5264 8984 5316 8993
rect 6276 8984 6328 9036
rect 4988 8916 5040 8968
rect 7656 8984 7708 9036
rect 8208 8984 8260 9036
rect 8576 8984 8628 9036
rect 9680 9052 9732 9104
rect 14556 9129 14565 9163
rect 14565 9129 14599 9163
rect 14599 9129 14608 9163
rect 14556 9120 14608 9129
rect 12348 8984 12400 9036
rect 13268 8984 13320 9036
rect 8852 8916 8904 8968
rect 11428 8916 11480 8968
rect 12164 8916 12216 8968
rect 12900 8916 12952 8968
rect 1400 8891 1452 8900
rect 1400 8857 1409 8891
rect 1409 8857 1443 8891
rect 1443 8857 1452 8891
rect 1400 8848 1452 8857
rect 2780 8891 2832 8900
rect 2780 8857 2789 8891
rect 2789 8857 2823 8891
rect 2823 8857 2832 8891
rect 2780 8848 2832 8857
rect 4620 8848 4672 8900
rect 5264 8848 5316 8900
rect 6644 8848 6696 8900
rect 7380 8848 7432 8900
rect 9680 8848 9732 8900
rect 4528 8780 4580 8832
rect 8300 8823 8352 8832
rect 8300 8789 8309 8823
rect 8309 8789 8343 8823
rect 8343 8789 8352 8823
rect 8300 8780 8352 8789
rect 8944 8780 8996 8832
rect 9772 8823 9824 8832
rect 9772 8789 9781 8823
rect 9781 8789 9815 8823
rect 9815 8789 9824 8823
rect 9772 8780 9824 8789
rect 10324 8780 10376 8832
rect 14464 8780 14516 8832
rect 3972 8678 4024 8730
rect 4036 8678 4088 8730
rect 4100 8678 4152 8730
rect 4164 8678 4216 8730
rect 9952 8678 10004 8730
rect 10016 8678 10068 8730
rect 10080 8678 10132 8730
rect 10144 8678 10196 8730
rect 15932 8678 15984 8730
rect 15996 8678 16048 8730
rect 16060 8678 16112 8730
rect 16124 8678 16176 8730
rect 8576 8576 8628 8628
rect 9680 8576 9732 8628
rect 12900 8619 12952 8628
rect 12900 8585 12909 8619
rect 12909 8585 12943 8619
rect 12943 8585 12952 8619
rect 12900 8576 12952 8585
rect 2320 8483 2372 8492
rect 2320 8449 2329 8483
rect 2329 8449 2363 8483
rect 2363 8449 2372 8483
rect 2320 8440 2372 8449
rect 4344 8440 4396 8492
rect 4712 8440 4764 8492
rect 7288 8440 7340 8492
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 9312 8440 9364 8492
rect 2780 8372 2832 8424
rect 3148 8372 3200 8424
rect 3424 8372 3476 8424
rect 2504 8304 2556 8356
rect 6000 8372 6052 8424
rect 8208 8304 8260 8356
rect 11060 8372 11112 8424
rect 12348 8415 12400 8424
rect 12348 8381 12357 8415
rect 12357 8381 12391 8415
rect 12391 8381 12400 8415
rect 12348 8372 12400 8381
rect 14464 8415 14516 8424
rect 14464 8381 14473 8415
rect 14473 8381 14507 8415
rect 14507 8381 14516 8415
rect 14464 8372 14516 8381
rect 14556 8372 14608 8424
rect 15476 8415 15528 8424
rect 15476 8381 15485 8415
rect 15485 8381 15519 8415
rect 15519 8381 15528 8415
rect 15476 8372 15528 8381
rect 16672 8415 16724 8424
rect 16672 8381 16681 8415
rect 16681 8381 16715 8415
rect 16715 8381 16724 8415
rect 16672 8372 16724 8381
rect 17500 8372 17552 8424
rect 11244 8304 11296 8356
rect 4712 8236 4764 8288
rect 5356 8279 5408 8288
rect 5356 8245 5365 8279
rect 5365 8245 5399 8279
rect 5399 8245 5408 8279
rect 5356 8236 5408 8245
rect 8484 8279 8536 8288
rect 8484 8245 8493 8279
rect 8493 8245 8527 8279
rect 8527 8245 8536 8279
rect 17132 8347 17184 8356
rect 17132 8313 17141 8347
rect 17141 8313 17175 8347
rect 17175 8313 17184 8347
rect 17132 8304 17184 8313
rect 8484 8236 8536 8245
rect 6962 8134 7014 8186
rect 7026 8134 7078 8186
rect 7090 8134 7142 8186
rect 7154 8134 7206 8186
rect 12942 8134 12994 8186
rect 13006 8134 13058 8186
rect 13070 8134 13122 8186
rect 13134 8134 13186 8186
rect 2504 8075 2556 8084
rect 2504 8041 2513 8075
rect 2513 8041 2547 8075
rect 2547 8041 2556 8075
rect 2504 8032 2556 8041
rect 2688 8032 2740 8084
rect 8484 8075 8536 8084
rect 8484 8041 8493 8075
rect 8493 8041 8527 8075
rect 8527 8041 8536 8075
rect 8484 8032 8536 8041
rect 8668 8032 8720 8084
rect 9128 8032 9180 8084
rect 17132 8032 17184 8084
rect 4528 8007 4580 8016
rect 4528 7973 4537 8007
rect 4537 7973 4571 8007
rect 4571 7973 4580 8007
rect 4528 7964 4580 7973
rect 7472 8007 7524 8016
rect 7472 7973 7481 8007
rect 7481 7973 7515 8007
rect 7515 7973 7524 8007
rect 7472 7964 7524 7973
rect 11060 8007 11112 8016
rect 11060 7973 11069 8007
rect 11069 7973 11103 8007
rect 11103 7973 11112 8007
rect 11060 7964 11112 7973
rect 7840 7939 7892 7948
rect 7840 7905 7849 7939
rect 7849 7905 7883 7939
rect 7883 7905 7892 7939
rect 7840 7896 7892 7905
rect 8668 7939 8720 7948
rect 8668 7905 8677 7939
rect 8677 7905 8711 7939
rect 8711 7905 8720 7939
rect 8668 7896 8720 7905
rect 8852 7939 8904 7948
rect 8852 7905 8861 7939
rect 8861 7905 8895 7939
rect 8895 7905 8904 7939
rect 8852 7896 8904 7905
rect 8944 7939 8996 7948
rect 8944 7905 8953 7939
rect 8953 7905 8987 7939
rect 8987 7905 8996 7939
rect 9128 7939 9180 7948
rect 8944 7896 8996 7905
rect 9128 7905 9137 7939
rect 9137 7905 9171 7939
rect 9171 7905 9180 7939
rect 9128 7896 9180 7905
rect 4712 7828 4764 7880
rect 9772 7760 9824 7812
rect 2504 7692 2556 7744
rect 8852 7692 8904 7744
rect 9588 7692 9640 7744
rect 16764 7692 16816 7744
rect 3972 7590 4024 7642
rect 4036 7590 4088 7642
rect 4100 7590 4152 7642
rect 4164 7590 4216 7642
rect 9952 7590 10004 7642
rect 10016 7590 10068 7642
rect 10080 7590 10132 7642
rect 10144 7590 10196 7642
rect 15932 7590 15984 7642
rect 15996 7590 16048 7642
rect 16060 7590 16112 7642
rect 16124 7590 16176 7642
rect 13360 7531 13412 7540
rect 13360 7497 13369 7531
rect 13369 7497 13403 7531
rect 13403 7497 13412 7531
rect 13360 7488 13412 7497
rect 2504 7463 2556 7472
rect 2504 7429 2513 7463
rect 2513 7429 2547 7463
rect 2547 7429 2556 7463
rect 2504 7420 2556 7429
rect 16764 7463 16816 7472
rect 16764 7429 16773 7463
rect 16773 7429 16807 7463
rect 16807 7429 16816 7463
rect 16764 7420 16816 7429
rect 2504 7284 2556 7336
rect 4620 7284 4672 7336
rect 6644 7327 6696 7336
rect 6644 7293 6653 7327
rect 6653 7293 6687 7327
rect 6687 7293 6696 7327
rect 6644 7284 6696 7293
rect 7288 7327 7340 7336
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 8944 7284 8996 7336
rect 12624 7284 12676 7336
rect 13820 7327 13872 7336
rect 6828 7216 6880 7268
rect 9128 7216 9180 7268
rect 13820 7293 13829 7327
rect 13829 7293 13863 7327
rect 13863 7293 13872 7327
rect 13820 7284 13872 7293
rect 15752 7327 15804 7336
rect 15752 7293 15761 7327
rect 15761 7293 15795 7327
rect 15795 7293 15804 7327
rect 15752 7284 15804 7293
rect 16672 7352 16724 7404
rect 16396 7327 16448 7336
rect 16396 7293 16405 7327
rect 16405 7293 16439 7327
rect 16439 7293 16448 7327
rect 16396 7284 16448 7293
rect 13636 7216 13688 7268
rect 3332 7148 3384 7200
rect 3792 7191 3844 7200
rect 3792 7157 3801 7191
rect 3801 7157 3835 7191
rect 3835 7157 3844 7191
rect 3792 7148 3844 7157
rect 5264 7148 5316 7200
rect 7748 7191 7800 7200
rect 7748 7157 7757 7191
rect 7757 7157 7791 7191
rect 7791 7157 7800 7191
rect 7748 7148 7800 7157
rect 12072 7148 12124 7200
rect 15752 7148 15804 7200
rect 16396 7148 16448 7200
rect 16488 7148 16540 7200
rect 6962 7046 7014 7098
rect 7026 7046 7078 7098
rect 7090 7046 7142 7098
rect 7154 7046 7206 7098
rect 12942 7046 12994 7098
rect 13006 7046 13058 7098
rect 13070 7046 13122 7098
rect 13134 7046 13186 7098
rect 3792 6944 3844 6996
rect 12072 6987 12124 6996
rect 4804 6919 4856 6928
rect 4804 6885 4813 6919
rect 4813 6885 4847 6919
rect 4847 6885 4856 6919
rect 4804 6876 4856 6885
rect 7840 6876 7892 6928
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 2504 6808 2556 6860
rect 3148 6851 3200 6860
rect 3148 6817 3157 6851
rect 3157 6817 3191 6851
rect 3191 6817 3200 6851
rect 3148 6808 3200 6817
rect 4712 6851 4764 6860
rect 4712 6817 4721 6851
rect 4721 6817 4755 6851
rect 4755 6817 4764 6851
rect 4712 6808 4764 6817
rect 4988 6851 5040 6860
rect 4988 6817 4997 6851
rect 4997 6817 5031 6851
rect 5031 6817 5040 6851
rect 4988 6808 5040 6817
rect 5724 6851 5776 6860
rect 5724 6817 5733 6851
rect 5733 6817 5767 6851
rect 5767 6817 5776 6851
rect 5724 6808 5776 6817
rect 5908 6851 5960 6860
rect 5908 6817 5917 6851
rect 5917 6817 5951 6851
rect 5951 6817 5960 6851
rect 5908 6808 5960 6817
rect 6644 6851 6696 6860
rect 6644 6817 6653 6851
rect 6653 6817 6687 6851
rect 6687 6817 6696 6851
rect 6644 6808 6696 6817
rect 8576 6808 8628 6860
rect 12072 6953 12081 6987
rect 12081 6953 12115 6987
rect 12115 6953 12124 6987
rect 12072 6944 12124 6953
rect 13360 6987 13412 6996
rect 13360 6953 13369 6987
rect 13369 6953 13403 6987
rect 13403 6953 13412 6987
rect 13360 6944 13412 6953
rect 13820 6987 13872 6996
rect 13820 6953 13829 6987
rect 13829 6953 13863 6987
rect 13863 6953 13872 6987
rect 13820 6944 13872 6953
rect 16488 6919 16540 6928
rect 9220 6808 9272 6860
rect 9772 6808 9824 6860
rect 10508 6808 10560 6860
rect 10692 6851 10744 6860
rect 10692 6817 10701 6851
rect 10701 6817 10735 6851
rect 10735 6817 10744 6851
rect 10692 6808 10744 6817
rect 10600 6740 10652 6792
rect 12624 6808 12676 6860
rect 13636 6851 13688 6860
rect 13636 6817 13645 6851
rect 13645 6817 13679 6851
rect 13679 6817 13688 6851
rect 14740 6851 14792 6860
rect 13636 6808 13688 6817
rect 14740 6817 14749 6851
rect 14749 6817 14783 6851
rect 14783 6817 14792 6851
rect 14740 6808 14792 6817
rect 16488 6885 16497 6919
rect 16497 6885 16531 6919
rect 16531 6885 16540 6919
rect 16488 6876 16540 6885
rect 18696 6851 18748 6860
rect 18696 6817 18705 6851
rect 18705 6817 18739 6851
rect 18739 6817 18748 6851
rect 18696 6808 18748 6817
rect 8668 6672 8720 6724
rect 9772 6672 9824 6724
rect 12164 6672 12216 6724
rect 13728 6740 13780 6792
rect 15016 6783 15068 6792
rect 15016 6749 15025 6783
rect 15025 6749 15059 6783
rect 15059 6749 15068 6783
rect 15016 6740 15068 6749
rect 3332 6604 3384 6656
rect 12348 6604 12400 6656
rect 12716 6604 12768 6656
rect 14372 6647 14424 6656
rect 14372 6613 14381 6647
rect 14381 6613 14415 6647
rect 14415 6613 14424 6647
rect 14372 6604 14424 6613
rect 3972 6502 4024 6554
rect 4036 6502 4088 6554
rect 4100 6502 4152 6554
rect 4164 6502 4216 6554
rect 9952 6502 10004 6554
rect 10016 6502 10068 6554
rect 10080 6502 10132 6554
rect 10144 6502 10196 6554
rect 15932 6502 15984 6554
rect 15996 6502 16048 6554
rect 16060 6502 16112 6554
rect 16124 6502 16176 6554
rect 1676 6332 1728 6384
rect 5908 6400 5960 6452
rect 9772 6443 9824 6452
rect 9772 6409 9781 6443
rect 9781 6409 9815 6443
rect 9815 6409 9824 6443
rect 9772 6400 9824 6409
rect 14372 6400 14424 6452
rect 12716 6375 12768 6384
rect 1584 6264 1636 6316
rect 12716 6341 12725 6375
rect 12725 6341 12759 6375
rect 12759 6341 12768 6375
rect 12716 6332 12768 6341
rect 6644 6196 6696 6248
rect 7932 6239 7984 6248
rect 7932 6205 7941 6239
rect 7941 6205 7975 6239
rect 7975 6205 7984 6239
rect 7932 6196 7984 6205
rect 8668 6264 8720 6316
rect 15752 6400 15804 6452
rect 15016 6332 15068 6384
rect 8576 6196 8628 6248
rect 6736 6171 6788 6180
rect 6736 6137 6745 6171
rect 6745 6137 6779 6171
rect 6779 6137 6788 6171
rect 6736 6128 6788 6137
rect 7840 6128 7892 6180
rect 9220 6128 9272 6180
rect 10508 6196 10560 6248
rect 10784 6196 10836 6248
rect 12348 6239 12400 6248
rect 12348 6205 12357 6239
rect 12357 6205 12391 6239
rect 12391 6205 12400 6239
rect 12348 6196 12400 6205
rect 14832 6239 14884 6248
rect 14832 6205 14841 6239
rect 14841 6205 14875 6239
rect 14875 6205 14884 6239
rect 14832 6196 14884 6205
rect 15292 6239 15344 6248
rect 10692 6128 10744 6180
rect 15292 6205 15301 6239
rect 15301 6205 15335 6239
rect 15335 6205 15344 6239
rect 15292 6196 15344 6205
rect 15476 6128 15528 6180
rect 12716 6103 12768 6112
rect 12716 6069 12725 6103
rect 12725 6069 12759 6103
rect 12759 6069 12768 6103
rect 12716 6060 12768 6069
rect 14832 6060 14884 6112
rect 16212 6060 16264 6112
rect 6962 5958 7014 6010
rect 7026 5958 7078 6010
rect 7090 5958 7142 6010
rect 7154 5958 7206 6010
rect 12942 5958 12994 6010
rect 13006 5958 13058 6010
rect 13070 5958 13122 6010
rect 13134 5958 13186 6010
rect 3516 5856 3568 5908
rect 4896 5856 4948 5908
rect 6644 5899 6696 5908
rect 3240 5831 3292 5840
rect 3240 5797 3249 5831
rect 3249 5797 3283 5831
rect 3283 5797 3292 5831
rect 3240 5788 3292 5797
rect 6644 5865 6653 5899
rect 6653 5865 6687 5899
rect 6687 5865 6696 5899
rect 6644 5856 6696 5865
rect 6828 5856 6880 5908
rect 7932 5856 7984 5908
rect 9220 5856 9272 5908
rect 10784 5899 10836 5908
rect 10784 5865 10793 5899
rect 10793 5865 10827 5899
rect 10827 5865 10836 5899
rect 10784 5856 10836 5865
rect 14740 5856 14792 5908
rect 12716 5788 12768 5840
rect 4436 5720 4488 5772
rect 4712 5720 4764 5772
rect 5908 5720 5960 5772
rect 10508 5720 10560 5772
rect 12348 5720 12400 5772
rect 12624 5763 12676 5772
rect 12624 5729 12633 5763
rect 12633 5729 12667 5763
rect 12667 5729 12676 5763
rect 12624 5720 12676 5729
rect 7288 5695 7340 5704
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 14740 5763 14792 5772
rect 14740 5729 14749 5763
rect 14749 5729 14783 5763
rect 14783 5729 14792 5763
rect 14740 5720 14792 5729
rect 15292 5763 15344 5772
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 15476 5763 15528 5772
rect 15476 5729 15485 5763
rect 15485 5729 15519 5763
rect 15519 5729 15528 5763
rect 15476 5720 15528 5729
rect 16396 5788 16448 5840
rect 16212 5763 16264 5772
rect 16212 5729 16221 5763
rect 16221 5729 16255 5763
rect 16255 5729 16264 5763
rect 16212 5720 16264 5729
rect 15568 5584 15620 5636
rect 16304 5652 16356 5704
rect 18420 5584 18472 5636
rect 18512 5516 18564 5568
rect 3972 5414 4024 5466
rect 4036 5414 4088 5466
rect 4100 5414 4152 5466
rect 4164 5414 4216 5466
rect 9952 5414 10004 5466
rect 10016 5414 10068 5466
rect 10080 5414 10132 5466
rect 10144 5414 10196 5466
rect 15932 5414 15984 5466
rect 15996 5414 16048 5466
rect 16060 5414 16112 5466
rect 16124 5414 16176 5466
rect 3240 5108 3292 5160
rect 4712 5108 4764 5160
rect 5356 5108 5408 5160
rect 16396 5176 16448 5228
rect 6368 5108 6420 5160
rect 12716 5108 12768 5160
rect 14280 5108 14332 5160
rect 14832 5108 14884 5160
rect 12440 5083 12492 5092
rect 2412 4972 2464 5024
rect 12440 5049 12449 5083
rect 12449 5049 12483 5083
rect 12483 5049 12492 5083
rect 12440 5040 12492 5049
rect 15568 5108 15620 5160
rect 16212 5151 16264 5160
rect 16212 5117 16221 5151
rect 16221 5117 16255 5151
rect 16255 5117 16264 5151
rect 16212 5108 16264 5117
rect 5908 5015 5960 5024
rect 5908 4981 5917 5015
rect 5917 4981 5951 5015
rect 5951 4981 5960 5015
rect 5908 4972 5960 4981
rect 15660 5015 15712 5024
rect 15660 4981 15669 5015
rect 15669 4981 15703 5015
rect 15703 4981 15712 5015
rect 15660 4972 15712 4981
rect 16488 4972 16540 5024
rect 6962 4870 7014 4922
rect 7026 4870 7078 4922
rect 7090 4870 7142 4922
rect 7154 4870 7206 4922
rect 12942 4870 12994 4922
rect 13006 4870 13058 4922
rect 13070 4870 13122 4922
rect 13134 4870 13186 4922
rect 1492 4811 1544 4820
rect 1492 4777 1501 4811
rect 1501 4777 1535 4811
rect 1535 4777 1544 4811
rect 1492 4768 1544 4777
rect 6368 4811 6420 4820
rect 6368 4777 6377 4811
rect 6377 4777 6411 4811
rect 6411 4777 6420 4811
rect 6368 4768 6420 4777
rect 3332 4743 3384 4752
rect 3332 4709 3341 4743
rect 3341 4709 3375 4743
rect 3375 4709 3384 4743
rect 3332 4700 3384 4709
rect 10508 4768 10560 4820
rect 14740 4768 14792 4820
rect 18512 4811 18564 4820
rect 18512 4777 18521 4811
rect 18521 4777 18555 4811
rect 18555 4777 18564 4811
rect 18512 4768 18564 4777
rect 8024 4700 8076 4752
rect 2412 4675 2464 4684
rect 2412 4641 2421 4675
rect 2421 4641 2455 4675
rect 2455 4641 2464 4675
rect 2412 4632 2464 4641
rect 10784 4700 10836 4752
rect 11152 4700 11204 4752
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 10692 4675 10744 4684
rect 10692 4641 10701 4675
rect 10701 4641 10735 4675
rect 10735 4641 10744 4675
rect 16488 4700 16540 4752
rect 10692 4632 10744 4641
rect 12164 4632 12216 4684
rect 16304 4632 16356 4684
rect 18696 4675 18748 4684
rect 4436 4564 4488 4616
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 7288 4564 7340 4573
rect 11612 4607 11664 4616
rect 8116 4496 8168 4548
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 15476 4607 15528 4616
rect 15476 4573 15485 4607
rect 15485 4573 15519 4607
rect 15519 4573 15528 4607
rect 15476 4564 15528 4573
rect 15660 4607 15712 4616
rect 15660 4573 15669 4607
rect 15669 4573 15703 4607
rect 15703 4573 15712 4607
rect 15660 4564 15712 4573
rect 18696 4641 18705 4675
rect 18705 4641 18739 4675
rect 18739 4641 18748 4675
rect 18696 4632 18748 4641
rect 2320 4471 2372 4480
rect 2320 4437 2329 4471
rect 2329 4437 2363 4471
rect 2363 4437 2372 4471
rect 2320 4428 2372 4437
rect 10508 4428 10560 4480
rect 16396 4496 16448 4548
rect 17960 4496 18012 4548
rect 18144 4496 18196 4548
rect 13084 4428 13136 4480
rect 3972 4326 4024 4378
rect 4036 4326 4088 4378
rect 4100 4326 4152 4378
rect 4164 4326 4216 4378
rect 9952 4326 10004 4378
rect 10016 4326 10068 4378
rect 10080 4326 10132 4378
rect 10144 4326 10196 4378
rect 15932 4326 15984 4378
rect 15996 4326 16048 4378
rect 16060 4326 16112 4378
rect 16124 4326 16176 4378
rect 7288 4224 7340 4276
rect 7748 4224 7800 4276
rect 10692 4224 10744 4276
rect 7196 4156 7248 4208
rect 8024 4088 8076 4140
rect 11612 4156 11664 4208
rect 7380 4020 7432 4072
rect 7748 4063 7800 4072
rect 7748 4029 7757 4063
rect 7757 4029 7791 4063
rect 7791 4029 7800 4063
rect 7748 4020 7800 4029
rect 8576 4020 8628 4072
rect 10324 4020 10376 4072
rect 12164 4088 12216 4140
rect 12440 4088 12492 4140
rect 13084 4063 13136 4072
rect 6552 3952 6604 4004
rect 9772 3884 9824 3936
rect 10600 3952 10652 4004
rect 11244 3952 11296 4004
rect 11336 3884 11388 3936
rect 11980 3927 12032 3936
rect 11980 3893 11989 3927
rect 11989 3893 12023 3927
rect 12023 3893 12032 3927
rect 11980 3884 12032 3893
rect 13084 4029 13093 4063
rect 13093 4029 13127 4063
rect 13127 4029 13136 4063
rect 13728 4088 13780 4140
rect 13084 4020 13136 4029
rect 13544 3927 13596 3936
rect 13544 3893 13553 3927
rect 13553 3893 13587 3927
rect 13587 3893 13596 3927
rect 13544 3884 13596 3893
rect 6962 3782 7014 3834
rect 7026 3782 7078 3834
rect 7090 3782 7142 3834
rect 7154 3782 7206 3834
rect 12942 3782 12994 3834
rect 13006 3782 13058 3834
rect 13070 3782 13122 3834
rect 13134 3782 13186 3834
rect 11152 3723 11204 3732
rect 5908 3612 5960 3664
rect 8116 3655 8168 3664
rect 8116 3621 8125 3655
rect 8125 3621 8159 3655
rect 8159 3621 8168 3655
rect 8116 3612 8168 3621
rect 11152 3689 11161 3723
rect 11161 3689 11195 3723
rect 11195 3689 11204 3723
rect 11152 3680 11204 3689
rect 13544 3680 13596 3732
rect 15384 3612 15436 3664
rect 8392 3544 8444 3596
rect 10968 3544 11020 3596
rect 11336 3544 11388 3596
rect 17868 3544 17920 3596
rect 14832 3519 14884 3528
rect 4896 3408 4948 3460
rect 4436 3340 4488 3392
rect 9772 3408 9824 3460
rect 14832 3485 14841 3519
rect 14841 3485 14875 3519
rect 14875 3485 14884 3519
rect 14832 3476 14884 3485
rect 15016 3519 15068 3528
rect 15016 3485 15025 3519
rect 15025 3485 15059 3519
rect 15059 3485 15068 3519
rect 15016 3476 15068 3485
rect 14004 3383 14056 3392
rect 14004 3349 14013 3383
rect 14013 3349 14047 3383
rect 14047 3349 14056 3383
rect 14004 3340 14056 3349
rect 14372 3383 14424 3392
rect 14372 3349 14381 3383
rect 14381 3349 14415 3383
rect 14415 3349 14424 3383
rect 14372 3340 14424 3349
rect 15476 3408 15528 3460
rect 16396 3476 16448 3528
rect 18512 3340 18564 3392
rect 3972 3238 4024 3290
rect 4036 3238 4088 3290
rect 4100 3238 4152 3290
rect 4164 3238 4216 3290
rect 9952 3238 10004 3290
rect 10016 3238 10068 3290
rect 10080 3238 10132 3290
rect 10144 3238 10196 3290
rect 15932 3238 15984 3290
rect 15996 3238 16048 3290
rect 16060 3238 16112 3290
rect 16124 3238 16176 3290
rect 5908 3179 5960 3188
rect 5908 3145 5917 3179
rect 5917 3145 5951 3179
rect 5951 3145 5960 3179
rect 5908 3136 5960 3145
rect 8392 3179 8444 3188
rect 8392 3145 8401 3179
rect 8401 3145 8435 3179
rect 8435 3145 8444 3179
rect 8392 3136 8444 3145
rect 10416 3136 10468 3188
rect 10968 3179 11020 3188
rect 10968 3145 10977 3179
rect 10977 3145 11011 3179
rect 11011 3145 11020 3179
rect 10968 3136 11020 3145
rect 2320 3000 2372 3052
rect 4896 3068 4948 3120
rect 1400 2975 1452 2984
rect 1400 2941 1409 2975
rect 1409 2941 1443 2975
rect 1443 2941 1452 2975
rect 1400 2932 1452 2941
rect 5724 2932 5776 2984
rect 8576 3000 8628 3052
rect 8300 2864 8352 2916
rect 9312 2932 9364 2984
rect 9956 2975 10008 2984
rect 9956 2941 9965 2975
rect 9965 2941 9999 2975
rect 9999 2941 10008 2975
rect 9956 2932 10008 2941
rect 14832 3136 14884 3188
rect 12164 3068 12216 3120
rect 15016 3068 15068 3120
rect 12808 3000 12860 3052
rect 16396 3000 16448 3052
rect 13268 2932 13320 2984
rect 13728 2975 13780 2984
rect 13728 2941 13737 2975
rect 13737 2941 13771 2975
rect 13771 2941 13780 2975
rect 13728 2932 13780 2941
rect 14372 2932 14424 2984
rect 15384 2932 15436 2984
rect 18696 2975 18748 2984
rect 18696 2941 18705 2975
rect 18705 2941 18739 2975
rect 18739 2941 18748 2975
rect 18696 2932 18748 2941
rect 13820 2907 13872 2916
rect 13820 2873 13829 2907
rect 13829 2873 13863 2907
rect 13863 2873 13872 2907
rect 13820 2864 13872 2873
rect 16396 2864 16448 2916
rect 7932 2796 7984 2848
rect 8484 2796 8536 2848
rect 12808 2796 12860 2848
rect 6962 2694 7014 2746
rect 7026 2694 7078 2746
rect 7090 2694 7142 2746
rect 7154 2694 7206 2746
rect 12942 2694 12994 2746
rect 13006 2694 13058 2746
rect 13070 2694 13122 2746
rect 13134 2694 13186 2746
rect 3424 2635 3476 2644
rect 2320 2524 2372 2576
rect 3424 2601 3433 2635
rect 3433 2601 3467 2635
rect 3467 2601 3476 2635
rect 3424 2592 3476 2601
rect 4804 2635 4856 2644
rect 4804 2601 4813 2635
rect 4813 2601 4847 2635
rect 4847 2601 4856 2635
rect 4804 2592 4856 2601
rect 5724 2592 5776 2644
rect 7932 2635 7984 2644
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 8300 2592 8352 2644
rect 9588 2635 9640 2644
rect 9588 2601 9597 2635
rect 9597 2601 9631 2635
rect 9631 2601 9640 2635
rect 9956 2635 10008 2644
rect 9588 2592 9640 2601
rect 9956 2601 9965 2635
rect 9965 2601 9999 2635
rect 9999 2601 10008 2635
rect 9956 2592 10008 2601
rect 10600 2635 10652 2644
rect 10600 2601 10609 2635
rect 10609 2601 10643 2635
rect 10643 2601 10652 2635
rect 10600 2592 10652 2601
rect 11980 2592 12032 2644
rect 13268 2592 13320 2644
rect 13820 2592 13872 2644
rect 15568 2635 15620 2644
rect 15568 2601 15577 2635
rect 15577 2601 15611 2635
rect 15611 2601 15620 2635
rect 15568 2592 15620 2601
rect 16580 2635 16632 2644
rect 16580 2601 16589 2635
rect 16589 2601 16623 2635
rect 16623 2601 16632 2635
rect 18512 2635 18564 2644
rect 16580 2592 16632 2601
rect 18512 2601 18521 2635
rect 18521 2601 18555 2635
rect 18555 2601 18564 2635
rect 18512 2592 18564 2601
rect 9312 2524 9364 2576
rect 14280 2524 14332 2576
rect 15016 2567 15068 2576
rect 15016 2533 15025 2567
rect 15025 2533 15059 2567
rect 15059 2533 15068 2567
rect 15016 2524 15068 2533
rect 15200 2524 15252 2576
rect 16396 2524 16448 2576
rect 480 2456 532 2508
rect 3240 2499 3292 2508
rect 3240 2465 3249 2499
rect 3249 2465 3283 2499
rect 3283 2465 3292 2499
rect 3240 2456 3292 2465
rect 4620 2499 4672 2508
rect 4620 2465 4629 2499
rect 4629 2465 4663 2499
rect 4663 2465 4672 2499
rect 4620 2456 4672 2465
rect 6000 2456 6052 2508
rect 8392 2456 8444 2508
rect 7288 2388 7340 2440
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 7840 2388 7892 2440
rect 9220 2456 9272 2508
rect 10600 2456 10652 2508
rect 11980 2499 12032 2508
rect 11980 2465 11989 2499
rect 11989 2465 12023 2499
rect 12023 2465 12032 2499
rect 11980 2456 12032 2465
rect 12808 2499 12860 2508
rect 12808 2465 12817 2499
rect 12817 2465 12851 2499
rect 12851 2465 12860 2499
rect 12808 2456 12860 2465
rect 14004 2499 14056 2508
rect 14004 2465 14013 2499
rect 14013 2465 14047 2499
rect 14047 2465 14056 2499
rect 14004 2456 14056 2465
rect 14372 2499 14424 2508
rect 14372 2465 14381 2499
rect 14381 2465 14415 2499
rect 14415 2465 14424 2499
rect 14372 2456 14424 2465
rect 13820 2388 13872 2440
rect 16580 2456 16632 2508
rect 17960 2363 18012 2372
rect 17960 2329 17969 2363
rect 17969 2329 18003 2363
rect 18003 2329 18012 2363
rect 17960 2320 18012 2329
rect 3972 2150 4024 2202
rect 4036 2150 4088 2202
rect 4100 2150 4152 2202
rect 4164 2150 4216 2202
rect 9952 2150 10004 2202
rect 10016 2150 10068 2202
rect 10080 2150 10132 2202
rect 10144 2150 10196 2202
rect 15932 2150 15984 2202
rect 15996 2150 16048 2202
rect 16060 2150 16112 2202
rect 16124 2150 16176 2202
rect 19156 1411 19208 1420
rect 19156 1377 19165 1411
rect 19165 1377 19199 1411
rect 19199 1377 19208 1411
rect 19156 1368 19208 1377
<< metal2 >>
rect 938 21540 994 22340
rect 2318 21540 2374 22340
rect 3698 21540 3754 22340
rect 5538 21540 5594 22340
rect 6918 21540 6974 22340
rect 8298 21540 8354 22340
rect 9678 21540 9734 22340
rect 11518 21540 11574 22340
rect 12898 21540 12954 22340
rect 14278 21540 14334 22340
rect 15658 21540 15714 22340
rect 17498 21540 17554 22340
rect 18878 21540 18934 22340
rect 952 19990 980 21540
rect 1490 20496 1546 20505
rect 1490 20431 1546 20440
rect 1504 20058 1532 20431
rect 1492 20052 1544 20058
rect 1492 19994 1544 20000
rect 940 19984 992 19990
rect 940 19926 992 19932
rect 2332 19922 2360 21540
rect 3712 19922 3740 21540
rect 5552 19922 5580 21540
rect 6932 20346 6960 21540
rect 6840 20318 6960 20346
rect 6840 19938 6868 20318
rect 6936 20156 7232 20176
rect 6992 20154 7016 20156
rect 7072 20154 7096 20156
rect 7152 20154 7176 20156
rect 7014 20102 7016 20154
rect 7078 20102 7090 20154
rect 7152 20102 7154 20154
rect 6992 20100 7016 20102
rect 7072 20100 7096 20102
rect 7152 20100 7176 20102
rect 6936 20080 7232 20100
rect 6840 19922 6960 19938
rect 8312 19922 8340 21540
rect 9692 19922 9720 21540
rect 11532 19922 11560 21540
rect 12912 20346 12940 21540
rect 12820 20318 12940 20346
rect 12820 19922 12848 20318
rect 12916 20156 13212 20176
rect 12972 20154 12996 20156
rect 13052 20154 13076 20156
rect 13132 20154 13156 20156
rect 12994 20102 12996 20154
rect 13058 20102 13070 20154
rect 13132 20102 13134 20154
rect 12972 20100 12996 20102
rect 13052 20100 13076 20102
rect 13132 20100 13156 20102
rect 12916 20080 13212 20100
rect 14292 19922 14320 21540
rect 15672 19922 15700 21540
rect 17512 19922 17540 21540
rect 18326 20496 18382 20505
rect 18326 20431 18382 20440
rect 18340 19922 18368 20431
rect 18892 19990 18920 21540
rect 18880 19984 18932 19990
rect 18880 19926 18932 19932
rect 1584 19916 1636 19922
rect 1584 19858 1636 19864
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 3700 19916 3752 19922
rect 3700 19858 3752 19864
rect 5540 19916 5592 19922
rect 6840 19916 6972 19922
rect 6840 19910 6920 19916
rect 5540 19858 5592 19864
rect 6920 19858 6972 19864
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 1596 19514 1624 19858
rect 9588 19780 9640 19786
rect 9588 19722 9640 19728
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 18420 19780 18472 19786
rect 18420 19722 18472 19728
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 2504 19712 2556 19718
rect 2504 19654 2556 19660
rect 3700 19712 3752 19718
rect 3700 19654 3752 19660
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 1398 17776 1454 17785
rect 1398 17711 1400 17720
rect 1452 17711 1454 17720
rect 1400 17682 1452 17688
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1398 15736 1454 15745
rect 1398 15671 1454 15680
rect 1412 15570 1440 15671
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1504 13870 1532 14418
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1412 13705 1440 13806
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 1504 13530 1532 13806
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1492 13524 1544 13530
rect 1492 13466 1544 13472
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1504 11665 1532 12038
rect 1490 11656 1546 11665
rect 1490 11591 1546 11600
rect 1596 9450 1624 13670
rect 1584 9444 1636 9450
rect 1584 9386 1636 9392
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1398 8936 1454 8945
rect 1398 8871 1400 8880
rect 1452 8871 1454 8880
rect 1400 8842 1452 8848
rect 1398 6896 1454 6905
rect 1398 6831 1400 6840
rect 1452 6831 1454 6840
rect 1400 6802 1452 6808
rect 1596 6322 1624 8978
rect 1688 6390 1716 17478
rect 1872 17066 1900 19246
rect 1860 17060 1912 17066
rect 1860 17002 1912 17008
rect 1872 15570 1900 17002
rect 1860 15564 1912 15570
rect 1860 15506 1912 15512
rect 1768 15360 1820 15366
rect 1768 15302 1820 15308
rect 1780 11762 1808 15302
rect 1964 13530 1992 19654
rect 2516 16574 2544 19654
rect 3424 19236 3476 19242
rect 3424 19178 3476 19184
rect 3436 18970 3464 19178
rect 3424 18964 3476 18970
rect 3424 18906 3476 18912
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 3620 17610 3648 18770
rect 3608 17604 3660 17610
rect 3608 17546 3660 17552
rect 3620 17134 3648 17546
rect 3608 17128 3660 17134
rect 3608 17070 3660 17076
rect 2516 16546 2728 16574
rect 2596 14476 2648 14482
rect 2596 14418 2648 14424
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2516 13870 2544 14214
rect 2504 13864 2556 13870
rect 2504 13806 2556 13812
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2056 11830 2084 13262
rect 2044 11824 2096 11830
rect 2044 11766 2096 11772
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 2056 9586 2084 11766
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 1872 9178 1900 9318
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 2332 8498 2360 9318
rect 2516 9110 2544 13806
rect 2608 13394 2636 14418
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2504 8356 2556 8362
rect 2504 8298 2556 8304
rect 2516 8090 2544 8298
rect 2700 8090 2728 16546
rect 3620 16046 3648 17070
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 2872 15904 2924 15910
rect 2872 15846 2924 15852
rect 2884 15638 2912 15846
rect 2872 15632 2924 15638
rect 2872 15574 2924 15580
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 3068 13530 3096 13670
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2884 12374 2912 13330
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3252 12986 3280 13262
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 2976 11898 3004 12242
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2792 10266 2820 11154
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2792 9994 2820 10202
rect 2884 10112 2912 11630
rect 2976 11354 3004 11630
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 3712 11286 3740 19654
rect 3946 19612 4242 19632
rect 4002 19610 4026 19612
rect 4082 19610 4106 19612
rect 4162 19610 4186 19612
rect 4024 19558 4026 19610
rect 4088 19558 4100 19610
rect 4162 19558 4164 19610
rect 4002 19556 4026 19558
rect 4082 19556 4106 19558
rect 4162 19556 4186 19558
rect 3946 19536 4242 19556
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 3896 18970 3924 19314
rect 4804 19236 4856 19242
rect 4804 19178 4856 19184
rect 5816 19236 5868 19242
rect 5816 19178 5868 19184
rect 4436 19168 4488 19174
rect 4436 19110 4488 19116
rect 3884 18964 3936 18970
rect 3884 18906 3936 18912
rect 4448 18834 4476 19110
rect 4436 18828 4488 18834
rect 4436 18770 4488 18776
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 3946 18524 4242 18544
rect 4002 18522 4026 18524
rect 4082 18522 4106 18524
rect 4162 18522 4186 18524
rect 4024 18470 4026 18522
rect 4088 18470 4100 18522
rect 4162 18470 4164 18522
rect 4002 18468 4026 18470
rect 4082 18468 4106 18470
rect 4162 18468 4186 18470
rect 3946 18448 4242 18468
rect 4356 18086 4384 18566
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4356 17660 4384 18022
rect 4448 17814 4476 18770
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4632 18222 4660 18702
rect 4816 18222 4844 19178
rect 5828 18970 5856 19178
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 4620 18216 4672 18222
rect 4540 18176 4620 18204
rect 4436 17808 4488 17814
rect 4436 17750 4488 17756
rect 4356 17632 4476 17660
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3804 17134 3832 17478
rect 3946 17436 4242 17456
rect 4002 17434 4026 17436
rect 4082 17434 4106 17436
rect 4162 17434 4186 17436
rect 4024 17382 4026 17434
rect 4088 17382 4100 17434
rect 4162 17382 4164 17434
rect 4002 17380 4026 17382
rect 4082 17380 4106 17382
rect 4162 17380 4186 17382
rect 3946 17360 4242 17380
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 4448 17066 4476 17632
rect 4540 17134 4568 18176
rect 4620 18158 4672 18164
rect 4804 18216 4856 18222
rect 4804 18158 4856 18164
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4632 17338 4660 17682
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4528 17128 4580 17134
rect 4528 17070 4580 17076
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4436 17060 4488 17066
rect 4436 17002 4488 17008
rect 3946 16348 4242 16368
rect 4002 16346 4026 16348
rect 4082 16346 4106 16348
rect 4162 16346 4186 16348
rect 4024 16294 4026 16346
rect 4088 16294 4100 16346
rect 4162 16294 4164 16346
rect 4002 16292 4026 16294
rect 4082 16292 4106 16294
rect 4162 16292 4186 16294
rect 3946 16272 4242 16292
rect 4448 15978 4476 17002
rect 4540 16182 4568 17070
rect 4724 16794 4752 17070
rect 4816 16998 4844 17478
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4528 16176 4580 16182
rect 4528 16118 4580 16124
rect 4252 15972 4304 15978
rect 4252 15914 4304 15920
rect 4436 15972 4488 15978
rect 4436 15914 4488 15920
rect 4264 15570 4292 15914
rect 4540 15570 4568 16118
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4436 15564 4488 15570
rect 4436 15506 4488 15512
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 4448 15366 4476 15506
rect 4436 15360 4488 15366
rect 4436 15302 4488 15308
rect 3946 15260 4242 15280
rect 4002 15258 4026 15260
rect 4082 15258 4106 15260
rect 4162 15258 4186 15260
rect 4024 15206 4026 15258
rect 4088 15206 4100 15258
rect 4162 15206 4164 15258
rect 4002 15204 4026 15206
rect 4082 15204 4106 15206
rect 4162 15204 4186 15206
rect 3946 15184 4242 15204
rect 4448 14958 4476 15302
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 3946 14172 4242 14192
rect 4002 14170 4026 14172
rect 4082 14170 4106 14172
rect 4162 14170 4186 14172
rect 4024 14118 4026 14170
rect 4088 14118 4100 14170
rect 4162 14118 4164 14170
rect 4002 14116 4026 14118
rect 4082 14116 4106 14118
rect 4162 14116 4186 14118
rect 3946 14096 4242 14116
rect 4540 13938 4568 15506
rect 4724 15026 4752 16730
rect 4816 16658 4844 16934
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4908 16590 4936 17138
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 5000 16658 5028 17070
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 4896 16584 4948 16590
rect 4896 16526 4948 16532
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4816 15638 4844 16390
rect 5172 15972 5224 15978
rect 5172 15914 5224 15920
rect 4804 15632 4856 15638
rect 4804 15574 4856 15580
rect 4988 15564 5040 15570
rect 4988 15506 5040 15512
rect 4804 15428 4856 15434
rect 4804 15370 4856 15376
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4816 14414 4844 15370
rect 5000 15162 5028 15506
rect 4988 15156 5040 15162
rect 4988 15098 5040 15104
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 4988 14476 5040 14482
rect 5092 14464 5120 14894
rect 5040 14436 5120 14464
rect 4988 14418 5040 14424
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4908 13870 4936 14214
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 3946 13084 4242 13104
rect 4002 13082 4026 13084
rect 4082 13082 4106 13084
rect 4162 13082 4186 13084
rect 4024 13030 4026 13082
rect 4088 13030 4100 13082
rect 4162 13030 4164 13082
rect 4002 13028 4026 13030
rect 4082 13028 4106 13030
rect 4162 13028 4186 13030
rect 3946 13008 4242 13028
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4172 12442 4200 12582
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 3946 11996 4242 12016
rect 4002 11994 4026 11996
rect 4082 11994 4106 11996
rect 4162 11994 4186 11996
rect 4024 11942 4026 11994
rect 4088 11942 4100 11994
rect 4162 11942 4164 11994
rect 4002 11940 4026 11942
rect 4082 11940 4106 11942
rect 4162 11940 4186 11942
rect 3946 11920 4242 11940
rect 4540 11898 4568 13126
rect 4816 12850 4844 13670
rect 4896 13252 4948 13258
rect 4896 13194 4948 13200
rect 4908 12918 4936 13194
rect 4896 12912 4948 12918
rect 4896 12854 4948 12860
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4160 11620 4212 11626
rect 4160 11562 4212 11568
rect 4804 11620 4856 11626
rect 4804 11562 4856 11568
rect 4172 11354 4200 11562
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 3700 11280 3752 11286
rect 3700 11222 3752 11228
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 3946 10908 4242 10928
rect 4002 10906 4026 10908
rect 4082 10906 4106 10908
rect 4162 10906 4186 10908
rect 4024 10854 4026 10906
rect 4088 10854 4100 10906
rect 4162 10854 4164 10906
rect 4002 10852 4026 10854
rect 4082 10852 4106 10854
rect 4162 10852 4186 10854
rect 3946 10832 4242 10852
rect 4632 10742 4660 11154
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 2964 10124 3016 10130
rect 2884 10084 2964 10112
rect 2964 10066 3016 10072
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2780 8900 2832 8906
rect 2780 8842 2832 8848
rect 2792 8430 2820 8842
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2516 7478 2544 7686
rect 2504 7472 2556 7478
rect 2504 7414 2556 7420
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2516 6866 2544 7278
rect 3160 6866 3188 8366
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 3344 6662 3372 7142
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 1676 6384 1728 6390
rect 1676 6326 1728 6332
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 3252 5166 3280 5782
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 1490 4856 1546 4865
rect 1490 4791 1492 4800
rect 1544 4791 1546 4800
rect 1492 4762 1544 4768
rect 2424 4690 2452 4966
rect 3344 4758 3372 6598
rect 3332 4752 3384 4758
rect 3332 4694 3384 4700
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2332 3058 2360 4422
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1412 2825 1440 2926
rect 1398 2816 1454 2825
rect 1398 2751 1454 2760
rect 2332 2582 2360 2994
rect 3436 2650 3464 8366
rect 3528 5914 3556 10066
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 3946 9820 4242 9840
rect 4002 9818 4026 9820
rect 4082 9818 4106 9820
rect 4162 9818 4186 9820
rect 4024 9766 4026 9818
rect 4088 9766 4100 9818
rect 4162 9766 4164 9818
rect 4002 9764 4026 9766
rect 4082 9764 4106 9766
rect 4162 9764 4186 9766
rect 3946 9744 4242 9764
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 3946 8732 4242 8752
rect 4002 8730 4026 8732
rect 4082 8730 4106 8732
rect 4162 8730 4186 8732
rect 4024 8678 4026 8730
rect 4088 8678 4100 8730
rect 4162 8678 4164 8730
rect 4002 8676 4026 8678
rect 4082 8676 4106 8678
rect 4162 8676 4186 8678
rect 3946 8656 4242 8676
rect 4356 8498 4384 9318
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 3946 7644 4242 7664
rect 4002 7642 4026 7644
rect 4082 7642 4106 7644
rect 4162 7642 4186 7644
rect 4024 7590 4026 7642
rect 4088 7590 4100 7642
rect 4162 7590 4164 7642
rect 4002 7588 4026 7590
rect 4082 7588 4106 7590
rect 4162 7588 4186 7590
rect 3946 7568 4242 7588
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 3804 7002 3832 7142
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3946 6556 4242 6576
rect 4002 6554 4026 6556
rect 4082 6554 4106 6556
rect 4162 6554 4186 6556
rect 4024 6502 4026 6554
rect 4088 6502 4100 6554
rect 4162 6502 4164 6554
rect 4002 6500 4026 6502
rect 4082 6500 4106 6502
rect 4162 6500 4186 6502
rect 3946 6480 4242 6500
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 4448 5778 4476 9862
rect 4540 9654 4568 10066
rect 4632 9722 4660 10678
rect 4724 10266 4752 11494
rect 4816 10810 4844 11562
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4816 10674 4844 10746
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4540 9110 4568 9590
rect 4528 9104 4580 9110
rect 4528 9046 4580 9052
rect 4632 8906 4660 9658
rect 4908 9602 4936 12038
rect 5000 11354 5028 14418
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 5092 13530 5120 13738
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 5092 12918 5120 13466
rect 5184 13258 5212 15914
rect 5356 15428 5408 15434
rect 5356 15370 5408 15376
rect 5368 15162 5396 15370
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5460 14958 5488 15302
rect 5632 15088 5684 15094
rect 5632 15030 5684 15036
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5172 13252 5224 13258
rect 5172 13194 5224 13200
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 5276 12434 5304 14758
rect 5460 14482 5488 14894
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 5460 13870 5488 14282
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5460 13530 5488 13806
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5644 12918 5672 15030
rect 5736 14958 5764 15302
rect 5920 14958 5948 16594
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5736 14482 5764 14894
rect 5920 14550 5948 14894
rect 5908 14544 5960 14550
rect 5908 14486 5960 14492
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5736 13870 5764 14214
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5920 12850 5948 14486
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5368 12442 5396 12718
rect 5184 12406 5304 12434
rect 5356 12436 5408 12442
rect 5080 12368 5132 12374
rect 5080 12310 5132 12316
rect 5092 11898 5120 12310
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 5092 10538 5120 11698
rect 5184 11218 5212 12406
rect 5356 12378 5408 12384
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5184 10606 5212 11154
rect 5368 11014 5396 12378
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 11898 5580 12174
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5460 11150 5488 11698
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 4816 9574 4936 9602
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4540 8022 4568 8774
rect 4528 8016 4580 8022
rect 4528 7958 4580 7964
rect 4632 7342 4660 8842
rect 4724 8498 4752 9046
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4724 8294 4752 8434
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4724 7886 4752 8230
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4724 6866 4752 7822
rect 4816 7018 4844 9574
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4908 9178 4936 9454
rect 5000 9450 5028 10066
rect 5092 10062 5120 10474
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 5092 9586 5120 9998
rect 5184 9926 5212 10542
rect 5368 10470 5396 10950
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 10062 5396 10406
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5172 9920 5224 9926
rect 5368 9908 5396 9998
rect 5172 9862 5224 9868
rect 5276 9880 5396 9908
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 5000 8974 5028 9386
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 5184 8922 5212 9862
rect 5276 9654 5304 9880
rect 5460 9738 5488 11086
rect 5368 9710 5488 9738
rect 5264 9648 5316 9654
rect 5264 9590 5316 9596
rect 5276 9042 5304 9590
rect 5368 9450 5396 9710
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5368 9178 5396 9386
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 4816 6990 4936 7018
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 3946 5468 4242 5488
rect 4002 5466 4026 5468
rect 4082 5466 4106 5468
rect 4162 5466 4186 5468
rect 4024 5414 4026 5466
rect 4088 5414 4100 5466
rect 4162 5414 4164 5466
rect 4002 5412 4026 5414
rect 4082 5412 4106 5414
rect 4162 5412 4186 5414
rect 3946 5392 4242 5412
rect 4724 5166 4752 5714
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 3946 4380 4242 4400
rect 4002 4378 4026 4380
rect 4082 4378 4106 4380
rect 4162 4378 4186 4380
rect 4024 4326 4026 4378
rect 4088 4326 4100 4378
rect 4162 4326 4164 4378
rect 4002 4324 4026 4326
rect 4082 4324 4106 4326
rect 4162 4324 4186 4326
rect 3946 4304 4242 4324
rect 4448 3398 4476 4558
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 3946 3292 4242 3312
rect 4002 3290 4026 3292
rect 4082 3290 4106 3292
rect 4162 3290 4186 3292
rect 4024 3238 4026 3290
rect 4088 3238 4100 3290
rect 4162 3238 4164 3290
rect 4002 3236 4026 3238
rect 4082 3236 4106 3238
rect 4162 3236 4186 3238
rect 3946 3216 4242 3236
rect 4816 2650 4844 6870
rect 4908 5914 4936 6990
rect 5000 6866 5028 8910
rect 5184 8906 5304 8922
rect 5184 8900 5316 8906
rect 5184 8894 5264 8900
rect 5264 8842 5316 8848
rect 5276 7206 5304 8842
rect 6012 8430 6040 19654
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 6460 19236 6512 19242
rect 6460 19178 6512 19184
rect 7288 19236 7340 19242
rect 7288 19178 7340 19184
rect 6472 18222 6500 19178
rect 6936 19068 7232 19088
rect 6992 19066 7016 19068
rect 7072 19066 7096 19068
rect 7152 19066 7176 19068
rect 7014 19014 7016 19066
rect 7078 19014 7090 19066
rect 7152 19014 7154 19066
rect 6992 19012 7016 19014
rect 7072 19012 7096 19014
rect 7152 19012 7176 19014
rect 6936 18992 7232 19012
rect 7300 18834 7328 19178
rect 8220 19174 8248 19246
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6748 18290 6776 18566
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6460 18216 6512 18222
rect 6460 18158 6512 18164
rect 6472 16572 6500 18158
rect 7288 18148 7340 18154
rect 7288 18090 7340 18096
rect 6936 17980 7232 18000
rect 6992 17978 7016 17980
rect 7072 17978 7096 17980
rect 7152 17978 7176 17980
rect 7014 17926 7016 17978
rect 7078 17926 7090 17978
rect 7152 17926 7154 17978
rect 6992 17924 7016 17926
rect 7072 17924 7096 17926
rect 7152 17924 7176 17926
rect 6936 17904 7232 17924
rect 7300 17882 7328 18090
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7392 17746 7420 18702
rect 7576 18698 7604 19110
rect 7748 18896 7800 18902
rect 7944 18873 7972 19110
rect 7748 18838 7800 18844
rect 7930 18864 7986 18873
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 7760 18426 7788 18838
rect 7930 18799 7932 18808
rect 7984 18799 7986 18808
rect 7932 18770 7984 18776
rect 8208 18692 8260 18698
rect 8208 18634 8260 18640
rect 7748 18420 7800 18426
rect 7748 18362 7800 18368
rect 8220 18154 8248 18634
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8312 18222 8340 18566
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 8208 18148 8260 18154
rect 8208 18090 8260 18096
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7760 17746 7788 18022
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7760 17134 7788 17682
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 6936 16892 7232 16912
rect 6992 16890 7016 16892
rect 7072 16890 7096 16892
rect 7152 16890 7176 16892
rect 7014 16838 7016 16890
rect 7078 16838 7090 16890
rect 7152 16838 7154 16890
rect 6992 16836 7016 16838
rect 7072 16836 7096 16838
rect 7152 16836 7176 16838
rect 6936 16816 7232 16836
rect 7576 16726 7604 16934
rect 7564 16720 7616 16726
rect 7564 16662 7616 16668
rect 6552 16584 6604 16590
rect 6472 16544 6552 16572
rect 6552 16526 6604 16532
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6196 10810 6224 14350
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 6288 12442 6316 12718
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6288 11286 6316 12378
rect 6564 11898 6592 16526
rect 6932 16250 6960 16526
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7196 16040 7248 16046
rect 7248 15988 7328 15994
rect 7196 15982 7328 15988
rect 7208 15966 7328 15982
rect 6936 15804 7232 15824
rect 6992 15802 7016 15804
rect 7072 15802 7096 15804
rect 7152 15802 7176 15804
rect 7014 15750 7016 15802
rect 7078 15750 7090 15802
rect 7152 15750 7154 15802
rect 6992 15748 7016 15750
rect 7072 15748 7096 15750
rect 7152 15748 7176 15750
rect 6936 15728 7232 15748
rect 7300 15094 7328 15966
rect 7484 15706 7512 16050
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7472 15564 7524 15570
rect 7472 15506 7524 15512
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7288 15088 7340 15094
rect 7288 15030 7340 15036
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 6936 14716 7232 14736
rect 6992 14714 7016 14716
rect 7072 14714 7096 14716
rect 7152 14714 7176 14716
rect 7014 14662 7016 14714
rect 7078 14662 7090 14714
rect 7152 14662 7154 14714
rect 6992 14660 7016 14662
rect 7072 14660 7096 14662
rect 7152 14660 7176 14662
rect 6936 14640 7232 14660
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7024 14074 7052 14418
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7208 13870 7236 14418
rect 7300 14074 7328 14758
rect 7392 14346 7420 14894
rect 7484 14618 7512 15506
rect 7668 15162 7696 15506
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7564 15088 7616 15094
rect 7564 15030 7616 15036
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7576 14414 7604 15030
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 12832 6868 13670
rect 6936 13628 7232 13648
rect 6992 13626 7016 13628
rect 7072 13626 7096 13628
rect 7152 13626 7176 13628
rect 7014 13574 7016 13626
rect 7078 13574 7090 13626
rect 7152 13574 7154 13626
rect 6992 13572 7016 13574
rect 7072 13572 7096 13574
rect 7152 13572 7176 13574
rect 6936 13552 7232 13572
rect 7196 13252 7248 13258
rect 7196 13194 7248 13200
rect 7208 12918 7236 13194
rect 7196 12912 7248 12918
rect 7196 12854 7248 12860
rect 6920 12844 6972 12850
rect 6840 12804 6920 12832
rect 6920 12786 6972 12792
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6840 12434 6868 12582
rect 6936 12540 7232 12560
rect 6992 12538 7016 12540
rect 7072 12538 7096 12540
rect 7152 12538 7176 12540
rect 7014 12486 7016 12538
rect 7078 12486 7090 12538
rect 7152 12486 7154 12538
rect 6992 12484 7016 12486
rect 7072 12484 7096 12486
rect 7152 12484 7176 12486
rect 6936 12464 7232 12484
rect 6840 12406 6960 12434
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6932 11762 6960 12406
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 7024 11626 7052 12242
rect 6368 11620 6420 11626
rect 6368 11562 6420 11568
rect 7012 11620 7064 11626
rect 7012 11562 7064 11568
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6196 10130 6224 10746
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6288 9654 6316 11222
rect 6380 11150 6408 11562
rect 6936 11452 7232 11472
rect 6992 11450 7016 11452
rect 7072 11450 7096 11452
rect 7152 11450 7176 11452
rect 7014 11398 7016 11450
rect 7078 11398 7090 11450
rect 7152 11398 7154 11450
rect 6992 11396 7016 11398
rect 7072 11396 7096 11398
rect 7152 11396 7176 11398
rect 6936 11376 7232 11396
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6380 10606 6408 11086
rect 7300 10810 7328 14010
rect 7484 13870 7512 14214
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7392 12918 7420 13738
rect 7668 12918 7696 14214
rect 7380 12912 7432 12918
rect 7380 12854 7432 12860
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6288 9042 6316 9590
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4908 3466 4936 5850
rect 5368 5166 5396 8230
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 4908 3126 4936 3402
rect 4896 3120 4948 3126
rect 4896 3062 4948 3068
rect 5736 2990 5764 6802
rect 5920 6458 5948 6802
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 5920 5030 5948 5714
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 6380 4826 6408 5102
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6564 4010 6592 10202
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6656 9586 6684 9862
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6656 8906 6684 9522
rect 6748 9450 6776 10542
rect 6936 10364 7232 10384
rect 6992 10362 7016 10364
rect 7072 10362 7096 10364
rect 7152 10362 7176 10364
rect 7014 10310 7016 10362
rect 7078 10310 7090 10362
rect 7152 10310 7154 10362
rect 6992 10308 7016 10310
rect 7072 10308 7096 10310
rect 7152 10308 7176 10310
rect 6936 10288 7232 10308
rect 7300 10130 7328 10746
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7300 9654 7328 10066
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6644 8900 6696 8906
rect 6644 8842 6696 8848
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6656 6866 6684 7278
rect 6840 7274 6868 9318
rect 6936 9276 7232 9296
rect 6992 9274 7016 9276
rect 7072 9274 7096 9276
rect 7152 9274 7176 9276
rect 7014 9222 7016 9274
rect 7078 9222 7090 9274
rect 7152 9222 7154 9274
rect 6992 9220 7016 9222
rect 7072 9220 7096 9222
rect 7152 9220 7176 9222
rect 6936 9200 7232 9220
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 6936 8188 7232 8208
rect 6992 8186 7016 8188
rect 7072 8186 7096 8188
rect 7152 8186 7176 8188
rect 7014 8134 7016 8186
rect 7078 8134 7090 8186
rect 7152 8134 7154 8186
rect 6992 8132 7016 8134
rect 7072 8132 7096 8134
rect 7152 8132 7176 8134
rect 6936 8112 7232 8132
rect 7300 7342 7328 8434
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 6828 7268 6880 7274
rect 6828 7210 6880 7216
rect 6644 6860 6696 6866
rect 6696 6820 6776 6848
rect 6644 6802 6696 6808
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6656 5914 6684 6190
rect 6748 6186 6776 6820
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6840 5914 6868 7210
rect 6936 7100 7232 7120
rect 6992 7098 7016 7100
rect 7072 7098 7096 7100
rect 7152 7098 7176 7100
rect 7014 7046 7016 7098
rect 7078 7046 7090 7098
rect 7152 7046 7154 7098
rect 6992 7044 7016 7046
rect 7072 7044 7096 7046
rect 7152 7044 7176 7046
rect 6936 7024 7232 7044
rect 6936 6012 7232 6032
rect 6992 6010 7016 6012
rect 7072 6010 7096 6012
rect 7152 6010 7176 6012
rect 7014 5958 7016 6010
rect 7078 5958 7090 6010
rect 7152 5958 7154 6010
rect 6992 5956 7016 5958
rect 7072 5956 7096 5958
rect 7152 5956 7176 5958
rect 6936 5936 7232 5956
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 7300 5710 7328 7278
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 6936 4924 7232 4944
rect 6992 4922 7016 4924
rect 7072 4922 7096 4924
rect 7152 4922 7176 4924
rect 7014 4870 7016 4922
rect 7078 4870 7090 4922
rect 7152 4870 7154 4922
rect 6992 4868 7016 4870
rect 7072 4868 7096 4870
rect 7152 4868 7176 4870
rect 6936 4848 7232 4868
rect 7300 4706 7328 5646
rect 7208 4678 7328 4706
rect 7208 4214 7236 4678
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7300 4282 7328 4558
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7196 4208 7248 4214
rect 7248 4156 7328 4162
rect 7196 4150 7328 4156
rect 7208 4134 7328 4150
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6936 3836 7232 3856
rect 6992 3834 7016 3836
rect 7072 3834 7096 3836
rect 7152 3834 7176 3836
rect 7014 3782 7016 3834
rect 7078 3782 7090 3834
rect 7152 3782 7154 3834
rect 6992 3780 7016 3782
rect 7072 3780 7096 3782
rect 7152 3780 7176 3782
rect 6936 3760 7232 3780
rect 5908 3664 5960 3670
rect 5908 3606 5960 3612
rect 5920 3194 5948 3606
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5736 2650 5764 2926
rect 6936 2748 7232 2768
rect 6992 2746 7016 2748
rect 7072 2746 7096 2748
rect 7152 2746 7176 2748
rect 7014 2694 7016 2746
rect 7078 2694 7090 2746
rect 7152 2694 7154 2746
rect 6992 2692 7016 2694
rect 7072 2692 7096 2694
rect 7152 2692 7176 2694
rect 6936 2672 7232 2692
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 2320 2576 2372 2582
rect 2320 2518 2372 2524
rect 480 2508 532 2514
rect 480 2450 532 2456
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 492 800 520 2450
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 1872 800 1900 2314
rect 3252 800 3280 2450
rect 3946 2204 4242 2224
rect 4002 2202 4026 2204
rect 4082 2202 4106 2204
rect 4162 2202 4186 2204
rect 4024 2150 4026 2202
rect 4088 2150 4100 2202
rect 4162 2150 4164 2202
rect 4002 2148 4026 2150
rect 4082 2148 4106 2150
rect 4162 2148 4186 2150
rect 3946 2128 4242 2148
rect 4632 800 4660 2450
rect 6012 800 6040 2450
rect 7300 2446 7328 4134
rect 7392 4078 7420 8842
rect 7484 8022 7512 11834
rect 7576 11150 7604 12718
rect 7760 12306 7788 17070
rect 8116 17060 8168 17066
rect 8116 17002 8168 17008
rect 8128 16182 8156 17002
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8116 16176 8168 16182
rect 8116 16118 8168 16124
rect 8312 15978 8340 16390
rect 8300 15972 8352 15978
rect 8300 15914 8352 15920
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 7840 14408 7892 14414
rect 7840 14350 7892 14356
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7668 11626 7696 12038
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7668 9654 7696 9998
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7668 9042 7696 9590
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7760 7206 7788 12242
rect 7852 10606 7880 14350
rect 7944 13326 7972 14894
rect 8116 14884 8168 14890
rect 8116 14826 8168 14832
rect 8128 14618 8156 14826
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8220 14482 8248 14894
rect 8312 14822 8340 15914
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8024 14340 8076 14346
rect 8024 14282 8076 14288
rect 8036 13870 8064 14282
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7944 12918 7972 13262
rect 7932 12912 7984 12918
rect 7932 12854 7984 12860
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8220 11694 8248 12718
rect 8312 11762 8340 14758
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8220 11354 8248 11630
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8312 10690 8340 11698
rect 8036 10662 8340 10690
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 8036 10538 8064 10662
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8220 10198 8248 10406
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8220 9042 8248 10134
rect 8312 10062 8340 10542
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8312 9586 8340 9998
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8220 8362 8248 8978
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7852 6934 7880 7890
rect 7840 6928 7892 6934
rect 7840 6870 7892 6876
rect 7852 6186 7880 6870
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 7840 6180 7892 6186
rect 7840 6122 7892 6128
rect 7944 5914 7972 6190
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7760 4078 7788 4218
rect 8036 4146 8064 4694
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 8128 3670 8156 4490
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8312 3074 8340 8774
rect 8404 8498 8432 19654
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8576 18896 8628 18902
rect 8574 18864 8576 18873
rect 8628 18864 8630 18873
rect 8574 18799 8630 18808
rect 8588 18698 8616 18799
rect 8576 18692 8628 18698
rect 8576 18634 8628 18640
rect 8864 18630 8892 19314
rect 9128 19236 9180 19242
rect 9128 19178 9180 19184
rect 9140 18970 9168 19178
rect 9128 18964 9180 18970
rect 9128 18906 9180 18912
rect 9312 18828 9364 18834
rect 9312 18770 9364 18776
rect 9128 18692 9180 18698
rect 9128 18634 9180 18640
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 9140 18222 9168 18634
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 9048 17134 9076 18158
rect 9324 18086 9352 18770
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 9404 16584 9456 16590
rect 9404 16526 9456 16532
rect 9416 14346 9444 16526
rect 9600 16046 9628 19722
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 9926 19612 10222 19632
rect 9982 19610 10006 19612
rect 10062 19610 10086 19612
rect 10142 19610 10166 19612
rect 10004 19558 10006 19610
rect 10068 19558 10080 19610
rect 10142 19558 10144 19610
rect 9982 19556 10006 19558
rect 10062 19556 10086 19558
rect 10142 19556 10166 19558
rect 9926 19536 10222 19556
rect 9926 18524 10222 18544
rect 9982 18522 10006 18524
rect 10062 18522 10086 18524
rect 10142 18522 10166 18524
rect 10004 18470 10006 18522
rect 10068 18470 10080 18522
rect 10142 18470 10144 18522
rect 9982 18468 10006 18470
rect 10062 18468 10086 18470
rect 10142 18468 10166 18470
rect 9926 18448 10222 18468
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 9692 17202 9720 17546
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 9926 17436 10222 17456
rect 9982 17434 10006 17436
rect 10062 17434 10086 17436
rect 10142 17434 10166 17436
rect 10004 17382 10006 17434
rect 10068 17382 10080 17434
rect 10142 17382 10144 17434
rect 9982 17380 10006 17382
rect 10062 17380 10086 17382
rect 10142 17380 10166 17382
rect 9926 17360 10222 17380
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9600 15570 9628 15982
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9692 15162 9720 16118
rect 9784 15978 9812 17138
rect 10336 17082 10364 17478
rect 10060 17066 10364 17082
rect 10048 17060 10364 17066
rect 10100 17054 10364 17060
rect 10048 17002 10100 17008
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9968 16658 9996 16934
rect 10244 16658 10272 17054
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 9926 16348 10222 16368
rect 9982 16346 10006 16348
rect 10062 16346 10086 16348
rect 10142 16346 10166 16348
rect 10004 16294 10006 16346
rect 10068 16294 10080 16346
rect 10142 16294 10144 16346
rect 9982 16292 10006 16294
rect 10062 16292 10086 16294
rect 10142 16292 10166 16294
rect 9926 16272 10222 16292
rect 10324 16176 10376 16182
rect 10324 16118 10376 16124
rect 10336 16046 10364 16118
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 10060 15706 10088 15982
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 9926 15260 10222 15280
rect 9982 15258 10006 15260
rect 10062 15258 10086 15260
rect 10142 15258 10166 15260
rect 10004 15206 10006 15258
rect 10068 15206 10080 15258
rect 10142 15206 10144 15258
rect 9982 15204 10006 15206
rect 10062 15204 10086 15206
rect 10142 15204 10166 15206
rect 9926 15184 10222 15204
rect 10428 15162 10456 16594
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10324 14884 10376 14890
rect 10324 14826 10376 14832
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9232 13870 9260 14214
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9416 13394 9444 14282
rect 9926 14172 10222 14192
rect 9982 14170 10006 14172
rect 10062 14170 10086 14172
rect 10142 14170 10166 14172
rect 10004 14118 10006 14170
rect 10068 14118 10080 14170
rect 10142 14118 10144 14170
rect 9982 14116 10006 14118
rect 10062 14116 10086 14118
rect 10142 14116 10166 14118
rect 9926 14096 10222 14116
rect 9496 13864 9548 13870
rect 9864 13864 9916 13870
rect 9548 13824 9864 13852
rect 9496 13806 9548 13812
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9140 12306 9168 13330
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8496 11218 8524 11494
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8496 10606 8524 11018
rect 8680 10606 8708 11630
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8956 10606 8984 11086
rect 8484 10600 8536 10606
rect 8668 10600 8720 10606
rect 8536 10560 8616 10588
rect 8484 10542 8536 10548
rect 8588 9042 8616 10560
rect 8668 10542 8720 10548
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8956 9722 8984 10542
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8496 8090 8524 8230
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8588 6866 8616 8570
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8680 7954 8708 8026
rect 8864 7954 8892 8910
rect 8956 8838 8984 9658
rect 9140 9178 9168 12242
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9324 11626 9352 12174
rect 9508 12102 9536 13330
rect 9600 13326 9628 13670
rect 9692 13530 9720 13824
rect 9864 13806 9916 13812
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9926 13084 10222 13104
rect 9982 13082 10006 13084
rect 10062 13082 10086 13084
rect 10142 13082 10166 13084
rect 10004 13030 10006 13082
rect 10068 13030 10080 13082
rect 10142 13030 10144 13082
rect 9982 13028 10006 13030
rect 10062 13028 10086 13030
rect 10142 13028 10166 13030
rect 9926 13008 10222 13028
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9508 11830 9536 12038
rect 9784 11898 9812 12786
rect 9926 11996 10222 12016
rect 9982 11994 10006 11996
rect 10062 11994 10086 11996
rect 10142 11994 10166 11996
rect 10004 11942 10006 11994
rect 10068 11942 10080 11994
rect 10142 11942 10144 11994
rect 9982 11940 10006 11942
rect 10062 11940 10086 11942
rect 10142 11940 10166 11942
rect 9926 11920 10222 11940
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9232 10130 9260 11154
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 8956 7954 8984 8774
rect 9140 8090 9168 9114
rect 9324 8498 9352 11562
rect 9416 10674 9444 11630
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9508 10606 9536 11766
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9692 10810 9720 11086
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9508 10130 9536 10542
rect 9692 10248 9720 10746
rect 9784 10606 9812 11630
rect 10336 11098 10364 14826
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10428 11626 10456 13262
rect 10520 12646 10548 19654
rect 11244 19372 11296 19378
rect 11244 19314 11296 19320
rect 10600 19236 10652 19242
rect 10600 19178 10652 19184
rect 10612 18970 10640 19178
rect 11256 18970 11284 19314
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11532 18902 11560 19110
rect 11520 18896 11572 18902
rect 11520 18838 11572 18844
rect 11520 18284 11572 18290
rect 11520 18226 11572 18232
rect 11532 17746 11560 18226
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 11256 17134 11284 17478
rect 11336 17264 11388 17270
rect 11336 17206 11388 17212
rect 11348 17134 11376 17206
rect 10600 17128 10652 17134
rect 11244 17128 11296 17134
rect 10652 17088 10732 17116
rect 10600 17070 10652 17076
rect 10704 16998 10732 17088
rect 11244 17070 11296 17076
rect 11336 17128 11388 17134
rect 11336 17070 11388 17076
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10796 16658 10824 17002
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10612 16250 10640 16594
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 10980 14618 11008 14894
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 11072 14074 11100 15982
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11532 14618 11560 14758
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11532 14414 11560 14554
rect 11520 14408 11572 14414
rect 11520 14350 11572 14356
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11428 13456 11480 13462
rect 11428 13398 11480 13404
rect 11440 12986 11468 13398
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 11072 12374 11100 12718
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11256 12434 11284 12650
rect 11256 12406 11376 12434
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10336 11070 10456 11098
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 9926 10908 10222 10928
rect 9982 10906 10006 10908
rect 10062 10906 10086 10908
rect 10142 10906 10166 10908
rect 10004 10854 10006 10906
rect 10068 10854 10080 10906
rect 10142 10854 10144 10906
rect 9982 10852 10006 10854
rect 10062 10852 10086 10854
rect 10142 10852 10166 10854
rect 9926 10832 10222 10852
rect 10336 10810 10364 10950
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9600 10220 9720 10248
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9600 10062 9628 10220
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9692 9110 9720 10066
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9692 8906 9720 9046
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9692 8634 9720 8842
rect 9784 8838 9812 10542
rect 9926 9820 10222 9840
rect 9982 9818 10006 9820
rect 10062 9818 10086 9820
rect 10142 9818 10166 9820
rect 10004 9766 10006 9818
rect 10068 9766 10080 9818
rect 10142 9766 10144 9818
rect 9982 9764 10006 9766
rect 10062 9764 10086 9766
rect 10142 9764 10166 9766
rect 9926 9744 10222 9764
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 9926 8732 10222 8752
rect 9982 8730 10006 8732
rect 10062 8730 10086 8732
rect 10142 8730 10166 8732
rect 10004 8678 10006 8730
rect 10068 8678 10080 8730
rect 10142 8678 10144 8730
rect 9982 8676 10006 8678
rect 10062 8676 10086 8678
rect 10142 8676 10166 8678
rect 9926 8656 10222 8676
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9140 7954 9168 8026
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 8864 7750 8892 7890
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8956 7342 8984 7890
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 9140 7274 9168 7890
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9128 7268 9180 7274
rect 9128 7210 9180 7216
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 8588 6254 8616 6802
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8680 6322 8708 6666
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 9232 6186 9260 6802
rect 9220 6180 9272 6186
rect 9220 6122 9272 6128
rect 9232 5914 9260 6122
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8404 3210 8432 3538
rect 8404 3194 8524 3210
rect 8392 3188 8524 3194
rect 8444 3182 8524 3188
rect 8392 3130 8444 3136
rect 8312 3046 8432 3074
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 7944 2650 7972 2790
rect 8312 2650 8340 2858
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8404 2514 8432 3046
rect 8496 2854 8524 3182
rect 8588 3058 8616 4014
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 9324 2582 9352 2926
rect 9600 2650 9628 7686
rect 9784 6866 9812 7754
rect 9926 7644 10222 7664
rect 9982 7642 10006 7644
rect 10062 7642 10086 7644
rect 10142 7642 10166 7644
rect 10004 7590 10006 7642
rect 10068 7590 10080 7642
rect 10142 7590 10144 7642
rect 9982 7588 10006 7590
rect 10062 7588 10086 7590
rect 10142 7588 10166 7590
rect 9926 7568 10222 7588
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9784 6458 9812 6666
rect 9926 6556 10222 6576
rect 9982 6554 10006 6556
rect 10062 6554 10086 6556
rect 10142 6554 10166 6556
rect 10004 6502 10006 6554
rect 10068 6502 10080 6554
rect 10142 6502 10144 6554
rect 9982 6500 10006 6502
rect 10062 6500 10086 6502
rect 10142 6500 10166 6502
rect 9926 6480 10222 6500
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9926 5468 10222 5488
rect 9982 5466 10006 5468
rect 10062 5466 10086 5468
rect 10142 5466 10166 5468
rect 10004 5414 10006 5466
rect 10068 5414 10080 5466
rect 10142 5414 10144 5466
rect 9982 5412 10006 5414
rect 10062 5412 10086 5414
rect 10142 5412 10166 5414
rect 9926 5392 10222 5412
rect 9926 4380 10222 4400
rect 9982 4378 10006 4380
rect 10062 4378 10086 4380
rect 10142 4378 10166 4380
rect 10004 4326 10006 4378
rect 10068 4326 10080 4378
rect 10142 4326 10144 4378
rect 9982 4324 10006 4326
rect 10062 4324 10086 4326
rect 10142 4324 10166 4326
rect 9926 4304 10222 4324
rect 10336 4078 10364 8774
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9784 3466 9812 3878
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9926 3292 10222 3312
rect 9982 3290 10006 3292
rect 10062 3290 10086 3292
rect 10142 3290 10166 3292
rect 10004 3238 10006 3290
rect 10068 3238 10080 3290
rect 10142 3238 10144 3290
rect 9982 3236 10006 3238
rect 10062 3236 10086 3238
rect 10142 3236 10166 3238
rect 9926 3216 10222 3236
rect 10428 3194 10456 11070
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11072 10674 11100 11018
rect 11164 10742 11192 12242
rect 11348 11150 11376 12406
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11152 10736 11204 10742
rect 11152 10678 11204 10684
rect 11348 10690 11376 11086
rect 11440 10810 11468 11154
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11164 10470 11192 10678
rect 11348 10662 11468 10690
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 10612 10198 10640 10406
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 11440 10062 11468 10662
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11440 8974 11468 9998
rect 11624 9178 11652 19654
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11716 18222 11744 18566
rect 11808 18358 11836 18770
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11716 17746 11744 18158
rect 11808 17882 11836 18294
rect 11796 17876 11848 17882
rect 11796 17818 11848 17824
rect 11900 17746 11928 19654
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12084 18222 12112 18770
rect 12360 18698 12388 18906
rect 12636 18698 12664 19246
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12348 18692 12400 18698
rect 12348 18634 12400 18640
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 12624 18692 12676 18698
rect 12624 18634 12676 18640
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 12256 18080 12308 18086
rect 12256 18022 12308 18028
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11716 17066 11744 17478
rect 12084 17338 12112 17682
rect 12268 17610 12296 18022
rect 12544 17814 12572 18634
rect 12728 18222 12756 18702
rect 12820 18426 12848 19110
rect 12916 19068 13212 19088
rect 12972 19066 12996 19068
rect 13052 19066 13076 19068
rect 13132 19066 13156 19068
rect 12994 19014 12996 19066
rect 13058 19014 13070 19066
rect 13132 19014 13134 19066
rect 12972 19012 12996 19014
rect 13052 19012 13076 19014
rect 13132 19012 13156 19014
rect 12916 18992 13212 19012
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 12728 17678 12756 18158
rect 12808 18148 12860 18154
rect 12808 18090 12860 18096
rect 12820 17882 12848 18090
rect 12916 17980 13212 18000
rect 12972 17978 12996 17980
rect 13052 17978 13076 17980
rect 13132 17978 13156 17980
rect 12994 17926 12996 17978
rect 13058 17926 13070 17978
rect 13132 17926 13134 17978
rect 12972 17924 12996 17926
rect 13052 17924 13076 17926
rect 13132 17924 13156 17926
rect 12916 17904 13212 17924
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12256 17604 12308 17610
rect 12256 17546 12308 17552
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 12268 17066 12296 17546
rect 12360 17542 12388 17614
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 11704 17060 11756 17066
rect 11704 17002 11756 17008
rect 12256 17060 12308 17066
rect 12256 17002 12308 17008
rect 11716 15366 11744 17002
rect 12820 16114 12848 17818
rect 13268 17808 13320 17814
rect 13268 17750 13320 17756
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 13096 17134 13124 17274
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 13188 17048 13216 17682
rect 13280 17338 13308 17750
rect 13464 17746 13492 18158
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 13360 17604 13412 17610
rect 13360 17546 13412 17552
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13372 17134 13400 17546
rect 13464 17338 13492 17682
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13188 17020 13308 17048
rect 12916 16892 13212 16912
rect 12972 16890 12996 16892
rect 13052 16890 13076 16892
rect 13132 16890 13156 16892
rect 12994 16838 12996 16890
rect 13058 16838 13070 16890
rect 13132 16838 13134 16890
rect 12972 16836 12996 16838
rect 13052 16836 13076 16838
rect 13132 16836 13156 16838
rect 12916 16816 13212 16836
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 13280 16046 13308 17020
rect 13556 16046 13584 17478
rect 11980 16040 12032 16046
rect 11980 15982 12032 15988
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11900 14958 11928 15438
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11900 12306 11928 13126
rect 11992 12714 12020 15982
rect 12072 15972 12124 15978
rect 12072 15914 12124 15920
rect 12164 15972 12216 15978
rect 12164 15914 12216 15920
rect 12084 15570 12112 15914
rect 12176 15706 12204 15914
rect 12916 15804 13212 15824
rect 12972 15802 12996 15804
rect 13052 15802 13076 15804
rect 13132 15802 13156 15804
rect 12994 15750 12996 15802
rect 13058 15750 13070 15802
rect 13132 15750 13134 15802
rect 12972 15748 12996 15750
rect 13052 15748 13076 15750
rect 13132 15748 13156 15750
rect 12916 15728 13212 15748
rect 13280 15706 13308 15982
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 12164 15700 12216 15706
rect 12164 15642 12216 15648
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12084 14890 12112 15506
rect 12176 14958 12204 15642
rect 13464 15638 13492 15846
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 13452 15632 13504 15638
rect 13452 15574 13504 15580
rect 12728 15366 12756 15574
rect 12440 15360 12492 15366
rect 12716 15360 12768 15366
rect 12492 15308 12572 15314
rect 12440 15302 12572 15308
rect 12716 15302 12768 15308
rect 12452 15286 12572 15302
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 12544 14414 12572 15286
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12544 13530 12572 14350
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 11980 12708 12032 12714
rect 11980 12650 12032 12656
rect 12636 12306 12664 12786
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 12728 12170 12756 15302
rect 12916 14716 13212 14736
rect 12972 14714 12996 14716
rect 13052 14714 13076 14716
rect 13132 14714 13156 14716
rect 12994 14662 12996 14714
rect 13058 14662 13070 14714
rect 13132 14662 13134 14714
rect 12972 14660 12996 14662
rect 13052 14660 13076 14662
rect 13132 14660 13156 14662
rect 12916 14640 13212 14660
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 12916 13628 13212 13648
rect 12972 13626 12996 13628
rect 13052 13626 13076 13628
rect 13132 13626 13156 13628
rect 12994 13574 12996 13626
rect 13058 13574 13070 13626
rect 13132 13574 13134 13626
rect 12972 13572 12996 13574
rect 13052 13572 13076 13574
rect 13132 13572 13156 13574
rect 12916 13552 13212 13572
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12820 13326 12848 13466
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12820 12306 12848 13262
rect 13280 13190 13308 13874
rect 13452 13728 13504 13734
rect 13452 13670 13504 13676
rect 13464 13258 13492 13670
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 12916 12540 13212 12560
rect 12972 12538 12996 12540
rect 13052 12538 13076 12540
rect 13132 12538 13156 12540
rect 12994 12486 12996 12538
rect 13058 12486 13070 12538
rect 13132 12486 13134 12538
rect 12972 12484 12996 12486
rect 13052 12484 13076 12486
rect 13132 12484 13156 12486
rect 12916 12464 13212 12484
rect 13280 12306 13308 12650
rect 13648 12434 13676 19722
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 13820 19236 13872 19242
rect 13820 19178 13872 19184
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13740 18766 13768 19110
rect 13832 18970 13860 19178
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13740 17066 13768 18566
rect 14292 17746 14320 18770
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13832 17066 13860 17478
rect 13728 17060 13780 17066
rect 13728 17002 13780 17008
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13740 16182 13768 17002
rect 13728 16176 13780 16182
rect 13728 16118 13780 16124
rect 13740 15502 13768 16118
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14292 15638 14320 15846
rect 14280 15632 14332 15638
rect 14280 15574 14332 15580
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13556 12406 13676 12434
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12636 11762 12664 12038
rect 12820 11898 12848 12242
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12544 11354 12572 11562
rect 12916 11452 13212 11472
rect 12972 11450 12996 11452
rect 13052 11450 13076 11452
rect 13132 11450 13156 11452
rect 12994 11398 12996 11450
rect 13058 11398 13070 11450
rect 13132 11398 13134 11450
rect 12972 11396 12996 11398
rect 13052 11396 13076 11398
rect 13132 11396 13156 11398
rect 12916 11376 13212 11396
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 12360 10130 12388 10406
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 11072 8022 11100 8366
rect 11244 8356 11296 8362
rect 11244 8298 11296 8304
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10520 6254 10548 6802
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 10520 4826 10548 5714
rect 10612 4842 10640 6734
rect 10704 6186 10732 6802
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10796 5914 10824 6190
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10612 4814 10824 4842
rect 10520 4486 10548 4762
rect 10612 4690 10640 4814
rect 10796 4758 10824 4814
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 11152 4752 11204 4758
rect 11152 4694 11204 4700
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 10704 4282 10732 4626
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 9968 2650 9996 2926
rect 10612 2650 10640 3946
rect 11164 3738 11192 4694
rect 11256 4010 11284 8298
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12084 7002 12112 7142
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12176 6730 12204 8910
rect 12360 8430 12388 8978
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12636 7342 12664 11018
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12728 10266 12756 10542
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 12916 10364 13212 10384
rect 12972 10362 12996 10364
rect 13052 10362 13076 10364
rect 13132 10362 13156 10364
rect 12994 10310 12996 10362
rect 13058 10310 13070 10362
rect 13132 10310 13134 10362
rect 12972 10308 12996 10310
rect 13052 10308 13076 10310
rect 13132 10308 13156 10310
rect 12916 10288 13212 10308
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 12176 4690 12204 6666
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12360 6254 12388 6598
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12360 5778 12388 6190
rect 12636 5778 12664 6802
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12728 6390 12756 6598
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12728 5846 12756 6054
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12728 5166 12756 5782
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11624 4214 11652 4558
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 12176 4146 12204 4626
rect 12452 4146 12480 5034
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11348 3602 11376 3878
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 10980 3194 11008 3538
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 11992 2650 12020 3878
rect 12176 3126 12204 4082
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 12820 3058 12848 9862
rect 12916 9276 13212 9296
rect 12972 9274 12996 9276
rect 13052 9274 13076 9276
rect 13132 9274 13156 9276
rect 12994 9222 12996 9274
rect 13058 9222 13070 9274
rect 13132 9222 13134 9274
rect 12972 9220 12996 9222
rect 13052 9220 13076 9222
rect 13132 9220 13156 9222
rect 12916 9200 13212 9220
rect 13280 9042 13308 10406
rect 13556 10266 13584 12406
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13648 11626 13676 12038
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13740 11354 13768 15438
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13832 12782 13860 13330
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13832 12374 13860 12718
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14200 11762 14228 12310
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13740 11218 13768 11290
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13648 10130 13676 10610
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12912 8634 12940 8910
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12916 8188 13212 8208
rect 12972 8186 12996 8188
rect 13052 8186 13076 8188
rect 13132 8186 13156 8188
rect 12994 8134 12996 8186
rect 13058 8134 13070 8186
rect 13132 8134 13134 8186
rect 12972 8132 12996 8134
rect 13052 8132 13076 8134
rect 13132 8132 13156 8134
rect 12916 8112 13212 8132
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 12916 7100 13212 7120
rect 12972 7098 12996 7100
rect 13052 7098 13076 7100
rect 13132 7098 13156 7100
rect 12994 7046 12996 7098
rect 13058 7046 13070 7098
rect 13132 7046 13134 7098
rect 12972 7044 12996 7046
rect 13052 7044 13076 7046
rect 13132 7044 13156 7046
rect 12916 7024 13212 7044
rect 13372 7002 13400 7482
rect 13636 7268 13688 7274
rect 13636 7210 13688 7216
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13648 6866 13676 7210
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13740 6798 13768 11154
rect 14384 10742 14412 19654
rect 15016 19304 15068 19310
rect 15016 19246 15068 19252
rect 14924 17808 14976 17814
rect 14924 17750 14976 17756
rect 14648 17672 14700 17678
rect 14648 17614 14700 17620
rect 14464 16040 14516 16046
rect 14464 15982 14516 15988
rect 14476 14940 14504 15982
rect 14556 15972 14608 15978
rect 14660 15960 14688 17614
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14844 17066 14872 17478
rect 14936 17270 14964 17750
rect 15028 17746 15056 19246
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15488 18902 15516 19110
rect 15672 18970 15700 19654
rect 15906 19612 16202 19632
rect 15962 19610 15986 19612
rect 16042 19610 16066 19612
rect 16122 19610 16146 19612
rect 15984 19558 15986 19610
rect 16048 19558 16060 19610
rect 16122 19558 16124 19610
rect 15962 19556 15986 19558
rect 16042 19556 16066 19558
rect 16122 19556 16146 19558
rect 15906 19536 16202 19556
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 15660 18964 15712 18970
rect 15660 18906 15712 18912
rect 17052 18902 17080 19110
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 17040 18896 17092 18902
rect 17040 18838 17092 18844
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 15906 18524 16202 18544
rect 15962 18522 15986 18524
rect 16042 18522 16066 18524
rect 16122 18522 16146 18524
rect 15984 18470 15986 18522
rect 16048 18470 16060 18522
rect 16122 18470 16124 18522
rect 15962 18468 15986 18470
rect 16042 18468 16066 18470
rect 16122 18468 16146 18470
rect 15906 18448 16202 18468
rect 16960 18290 16988 18702
rect 17236 18630 17264 19246
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17236 18290 17264 18566
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 15016 17740 15068 17746
rect 15016 17682 15068 17688
rect 14924 17264 14976 17270
rect 14924 17206 14976 17212
rect 14832 17060 14884 17066
rect 14832 17002 14884 17008
rect 14936 16402 14964 17206
rect 14608 15932 14688 15960
rect 14556 15914 14608 15920
rect 14556 14952 14608 14958
rect 14476 14912 14556 14940
rect 14556 14894 14608 14900
rect 14660 14822 14688 15932
rect 14844 16374 14964 16402
rect 14844 15910 14872 16374
rect 15028 16046 15056 17682
rect 15906 17436 16202 17456
rect 15962 17434 15986 17436
rect 16042 17434 16066 17436
rect 16122 17434 16146 17436
rect 15984 17382 15986 17434
rect 16048 17382 16060 17434
rect 16122 17382 16124 17434
rect 15962 17380 15986 17382
rect 16042 17380 16066 17382
rect 16122 17380 16146 17382
rect 15906 17360 16202 17380
rect 16396 17196 16448 17202
rect 16396 17138 16448 17144
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 16408 16794 16436 17138
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16592 16794 16620 16934
rect 16396 16788 16448 16794
rect 16396 16730 16448 16736
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16684 16726 16712 16934
rect 16672 16720 16724 16726
rect 16672 16662 16724 16668
rect 16776 16658 16804 17070
rect 17040 17060 17092 17066
rect 17040 17002 17092 17008
rect 17052 16658 17080 17002
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 15906 16348 16202 16368
rect 15962 16346 15986 16348
rect 16042 16346 16066 16348
rect 16122 16346 16146 16348
rect 15984 16294 15986 16346
rect 16048 16294 16060 16346
rect 16122 16294 16124 16346
rect 15962 16292 15986 16294
rect 16042 16292 16066 16294
rect 16122 16292 16146 16294
rect 15906 16272 16202 16292
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 14844 15094 14872 15846
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 14832 15088 14884 15094
rect 14832 15030 14884 15036
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14660 14074 14688 14758
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14752 13326 14780 14758
rect 14844 13394 14872 14894
rect 14936 14822 14964 15642
rect 15028 15366 15056 15982
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15212 15638 15240 15846
rect 15200 15632 15252 15638
rect 15200 15574 15252 15580
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 15660 14068 15712 14074
rect 15764 14056 15792 15302
rect 15906 15260 16202 15280
rect 15962 15258 15986 15260
rect 16042 15258 16066 15260
rect 16122 15258 16146 15260
rect 15984 15206 15986 15258
rect 16048 15206 16060 15258
rect 16122 15206 16124 15258
rect 15962 15204 15986 15206
rect 16042 15204 16066 15206
rect 16122 15204 16146 15206
rect 15906 15184 16202 15204
rect 16408 14958 16436 16050
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 16592 15570 16620 15914
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 15906 14172 16202 14192
rect 15962 14170 15986 14172
rect 16042 14170 16066 14172
rect 16122 14170 16146 14172
rect 15984 14118 15986 14170
rect 16048 14118 16060 14170
rect 16122 14118 16124 14170
rect 15962 14116 15986 14118
rect 16042 14116 16066 14118
rect 16122 14116 16146 14118
rect 15906 14096 16202 14116
rect 16408 14074 16436 14894
rect 16396 14068 16448 14074
rect 15764 14028 15884 14056
rect 15660 14010 15712 14016
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15028 13394 15056 13670
rect 15304 13530 15332 13806
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15396 13410 15424 13466
rect 14832 13388 14884 13394
rect 14832 13330 14884 13336
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 15120 13382 15424 13410
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14844 13274 14872 13330
rect 15120 13274 15148 13382
rect 14752 12850 14780 13262
rect 14844 13246 15148 13274
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 15396 12434 15424 13262
rect 15488 13258 15516 13806
rect 15672 13326 15700 14010
rect 15856 13938 15884 14028
rect 16396 14010 16448 14016
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15764 13394 15792 13806
rect 15856 13394 15884 13874
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15476 13252 15528 13258
rect 15476 13194 15528 13200
rect 15488 12986 15516 13194
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 15906 13084 16202 13104
rect 15962 13082 15986 13084
rect 16042 13082 16066 13084
rect 16122 13082 16146 13084
rect 15984 13030 15986 13082
rect 16048 13030 16060 13082
rect 16122 13030 16124 13082
rect 15962 13028 15986 13030
rect 16042 13028 16066 13030
rect 16122 13028 16146 13030
rect 15906 13008 16202 13028
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15304 12406 15424 12434
rect 16304 12436 16356 12442
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14936 11626 14964 12038
rect 15304 11762 15332 12406
rect 16304 12378 16356 12384
rect 15906 11996 16202 12016
rect 15962 11994 15986 11996
rect 16042 11994 16066 11996
rect 16122 11994 16146 11996
rect 15984 11942 15986 11994
rect 16048 11942 16060 11994
rect 16122 11942 16124 11994
rect 15962 11940 15986 11942
rect 16042 11940 16066 11942
rect 16122 11940 16146 11942
rect 15906 11920 16202 11940
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 16316 11694 16344 12378
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 14924 11620 14976 11626
rect 14924 11562 14976 11568
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 16040 11218 16068 11562
rect 16408 11286 16436 13126
rect 16592 12782 16620 15506
rect 16776 14618 16804 16594
rect 17236 16590 17264 17138
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17132 15972 17184 15978
rect 17132 15914 17184 15920
rect 17144 15706 17172 15914
rect 17236 15706 17264 16526
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 16960 15570 16988 15642
rect 17328 15586 17356 19314
rect 17512 17134 17540 19654
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 18064 18834 18092 19110
rect 18144 18896 18196 18902
rect 18144 18838 18196 18844
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 18064 16658 18092 18770
rect 18052 16652 18104 16658
rect 18052 16594 18104 16600
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 17972 15978 18000 16390
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 17236 15570 17356 15586
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 17224 15564 17356 15570
rect 17276 15558 17356 15564
rect 17408 15564 17460 15570
rect 17224 15506 17276 15512
rect 17408 15506 17460 15512
rect 17592 15564 17644 15570
rect 17592 15506 17644 15512
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17420 14890 17448 15506
rect 17604 15026 17632 15506
rect 17880 15366 17908 15506
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 17880 14958 17908 15302
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17408 14884 17460 14890
rect 17408 14826 17460 14832
rect 17592 14884 17644 14890
rect 17592 14826 17644 14832
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 17604 14482 17632 14826
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17604 13870 17632 14418
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 17788 13870 17816 14350
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17420 13530 17448 13806
rect 17500 13796 17552 13802
rect 17500 13738 17552 13744
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17512 13394 17540 13738
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17144 12782 17172 13330
rect 17788 13258 17816 13806
rect 17776 13252 17828 13258
rect 17776 13194 17828 13200
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17144 12434 17172 12718
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17144 12406 17356 12434
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16868 11694 16896 12242
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17144 11286 17172 11494
rect 17328 11354 17356 12406
rect 17512 12374 17540 12582
rect 17500 12368 17552 12374
rect 17500 12310 17552 12316
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 16396 11280 16448 11286
rect 16396 11222 16448 11228
rect 17132 11280 17184 11286
rect 17132 11222 17184 11228
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15120 10266 15148 10542
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15120 10130 15148 10202
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 14568 9518 14596 10066
rect 15396 9722 15424 10542
rect 15488 10266 15516 10950
rect 15906 10908 16202 10928
rect 15962 10906 15986 10908
rect 16042 10906 16066 10908
rect 16122 10906 16146 10908
rect 15984 10854 15986 10906
rect 16048 10854 16060 10906
rect 16122 10854 16124 10906
rect 15962 10852 15986 10854
rect 16042 10852 16066 10854
rect 16122 10852 16146 10854
rect 15906 10832 16202 10852
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 15764 9926 15792 10406
rect 17972 10266 18000 15302
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 18064 13190 18092 13466
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 18064 12714 18092 13126
rect 18052 12708 18104 12714
rect 18052 12650 18104 12656
rect 18064 12442 18092 12650
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15764 9518 15792 9862
rect 15906 9820 16202 9840
rect 15962 9818 15986 9820
rect 16042 9818 16066 9820
rect 16122 9818 16146 9820
rect 15984 9766 15986 9818
rect 16048 9766 16060 9818
rect 16122 9766 16124 9818
rect 15962 9764 15986 9766
rect 16042 9764 16066 9766
rect 16122 9764 16146 9766
rect 15906 9744 16202 9764
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 14568 9178 14596 9454
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14476 8430 14504 8774
rect 14568 8430 14596 9114
rect 15488 8430 15516 9386
rect 15906 8732 16202 8752
rect 15962 8730 15986 8732
rect 16042 8730 16066 8732
rect 16122 8730 16146 8732
rect 15984 8678 15986 8730
rect 16048 8678 16060 8730
rect 16122 8678 16124 8730
rect 15962 8676 15986 8678
rect 16042 8676 16066 8678
rect 16122 8676 16146 8678
rect 15906 8656 16202 8676
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15906 7644 16202 7664
rect 15962 7642 15986 7644
rect 16042 7642 16066 7644
rect 16122 7642 16146 7644
rect 15984 7590 15986 7642
rect 16048 7590 16060 7642
rect 16122 7590 16124 7642
rect 15962 7588 15986 7590
rect 16042 7588 16066 7590
rect 16122 7588 16146 7590
rect 15906 7568 16202 7588
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 13832 7002 13860 7278
rect 15764 7206 15792 7278
rect 16408 7206 16436 7278
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14384 6458 14412 6598
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 12916 6012 13212 6032
rect 12972 6010 12996 6012
rect 13052 6010 13076 6012
rect 13132 6010 13156 6012
rect 12994 5958 12996 6010
rect 13058 5958 13070 6010
rect 13132 5958 13134 6010
rect 12972 5956 12996 5958
rect 13052 5956 13076 5958
rect 13132 5956 13156 5958
rect 12916 5936 13212 5956
rect 14752 5914 14780 6802
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15028 6390 15056 6734
rect 15764 6458 15792 7142
rect 16500 6934 16528 7142
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 15906 6556 16202 6576
rect 15962 6554 15986 6556
rect 16042 6554 16066 6556
rect 16122 6554 16146 6556
rect 15984 6502 15986 6554
rect 16048 6502 16060 6554
rect 16122 6502 16124 6554
rect 15962 6500 15986 6502
rect 16042 6500 16066 6502
rect 16122 6500 16146 6502
rect 15906 6480 16202 6500
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15016 6384 15068 6390
rect 15016 6326 15068 6332
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 14844 6118 14872 6190
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 12916 4924 13212 4944
rect 12972 4922 12996 4924
rect 13052 4922 13076 4924
rect 13132 4922 13156 4924
rect 12994 4870 12996 4922
rect 13058 4870 13070 4922
rect 13132 4870 13134 4922
rect 12972 4868 12996 4870
rect 13052 4868 13076 4870
rect 13132 4868 13156 4870
rect 12916 4848 13212 4868
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13096 4078 13124 4422
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 12916 3836 13212 3856
rect 12972 3834 12996 3836
rect 13052 3834 13076 3836
rect 13132 3834 13156 3836
rect 12994 3782 12996 3834
rect 13058 3782 13070 3834
rect 13132 3782 13134 3834
rect 12972 3780 12996 3782
rect 13052 3780 13076 3782
rect 13132 3780 13156 3782
rect 12916 3760 13212 3780
rect 13556 3738 13584 3878
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 13740 2990 13768 4082
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 10600 2644 10652 2650
rect 10600 2586 10652 2592
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 9312 2576 9364 2582
rect 9312 2518 9364 2524
rect 12820 2514 12848 2790
rect 12916 2748 13212 2768
rect 12972 2746 12996 2748
rect 13052 2746 13076 2748
rect 13132 2746 13156 2748
rect 12994 2694 12996 2746
rect 13058 2694 13070 2746
rect 13132 2694 13134 2746
rect 12972 2692 12996 2694
rect 13052 2692 13076 2694
rect 13132 2692 13156 2694
rect 12916 2672 13212 2692
rect 13280 2650 13308 2926
rect 13820 2916 13872 2922
rect 13820 2858 13872 2864
rect 13832 2650 13860 2858
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 14016 2514 14044 3334
rect 14292 2582 14320 5102
rect 14752 4826 14780 5714
rect 14844 5166 14872 6054
rect 15304 5778 15332 6190
rect 15476 6180 15528 6186
rect 15476 6122 15528 6128
rect 15488 5778 15516 6122
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16224 5778 16252 6054
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 15568 5636 15620 5642
rect 15568 5578 15620 5584
rect 15580 5166 15608 5578
rect 15906 5468 16202 5488
rect 15962 5466 15986 5468
rect 16042 5466 16066 5468
rect 16122 5466 16146 5468
rect 15984 5414 15986 5466
rect 16048 5414 16060 5466
rect 16122 5414 16124 5466
rect 15962 5412 15986 5414
rect 16042 5412 16066 5414
rect 16122 5412 16146 5414
rect 15906 5392 16202 5412
rect 16316 5250 16344 5646
rect 16224 5222 16344 5250
rect 16408 5234 16436 5782
rect 16396 5228 16448 5234
rect 16224 5166 16252 5222
rect 16396 5170 16448 5176
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 15476 4616 15528 4622
rect 15476 4558 15528 4564
rect 15384 3664 15436 3670
rect 15384 3606 15436 3612
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14384 2990 14412 3334
rect 14844 3194 14872 3470
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 15028 3126 15056 3470
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14280 2576 14332 2582
rect 14280 2518 14332 2524
rect 14384 2514 14412 2926
rect 15028 2582 15056 3062
rect 15396 2990 15424 3606
rect 15488 3466 15516 4558
rect 15476 3460 15528 3466
rect 15476 3402 15528 3408
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 15580 2650 15608 5102
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 15672 4622 15700 4966
rect 16500 4758 16528 4966
rect 16488 4752 16540 4758
rect 16488 4694 16540 4700
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 15906 4380 16202 4400
rect 15962 4378 15986 4380
rect 16042 4378 16066 4380
rect 16122 4378 16146 4380
rect 15984 4326 15986 4378
rect 16048 4326 16060 4378
rect 16122 4326 16124 4378
rect 15962 4324 15986 4326
rect 16042 4324 16066 4326
rect 16122 4324 16146 4326
rect 15906 4304 16202 4324
rect 15906 3292 16202 3312
rect 15962 3290 15986 3292
rect 16042 3290 16066 3292
rect 16122 3290 16146 3292
rect 15984 3238 15986 3290
rect 16048 3238 16060 3290
rect 16122 3238 16124 3290
rect 15962 3236 15986 3238
rect 16042 3236 16066 3238
rect 16122 3236 16146 3238
rect 15906 3216 16202 3236
rect 16316 2938 16344 4626
rect 16396 4548 16448 4554
rect 16396 4490 16448 4496
rect 16408 3534 16436 4490
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16408 3058 16436 3470
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16316 2922 16436 2938
rect 16316 2916 16448 2922
rect 16316 2910 16396 2916
rect 16396 2858 16448 2864
rect 15568 2644 15620 2650
rect 15568 2586 15620 2592
rect 16408 2582 16436 2858
rect 16592 2650 16620 10202
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17512 8430 17540 9862
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 17500 8424 17552 8430
rect 17500 8366 17552 8372
rect 16684 7410 16712 8366
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 17144 8090 17172 8298
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16776 7478 16804 7686
rect 16764 7472 16816 7478
rect 16764 7414 16816 7420
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 18156 4554 18184 18838
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 18248 18154 18276 18566
rect 18236 18148 18288 18154
rect 18236 18090 18288 18096
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 18248 11898 18276 12310
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18432 5642 18460 19722
rect 18696 18692 18748 18698
rect 18696 18634 18748 18640
rect 18708 18465 18736 18634
rect 18694 18456 18750 18465
rect 18694 18391 18750 18400
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18524 14074 18552 16730
rect 18694 15736 18750 15745
rect 18694 15671 18750 15680
rect 18708 15570 18736 15671
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18512 14068 18564 14074
rect 18512 14010 18564 14016
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18708 13705 18736 13806
rect 18694 13696 18750 13705
rect 18694 13631 18750 13640
rect 18696 11688 18748 11694
rect 18694 11656 18696 11665
rect 18748 11656 18750 11665
rect 18694 11591 18750 11600
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18524 9654 18552 10474
rect 18512 9648 18564 9654
rect 18512 9590 18564 9596
rect 18694 9616 18750 9625
rect 18694 9551 18750 9560
rect 18708 9518 18736 9551
rect 18696 9512 18748 9518
rect 18696 9454 18748 9460
rect 18694 6896 18750 6905
rect 18694 6831 18696 6840
rect 18748 6831 18750 6840
rect 18696 6802 18748 6808
rect 18420 5636 18472 5642
rect 18420 5578 18472 5584
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18524 4826 18552 5510
rect 18694 4856 18750 4865
rect 18512 4820 18564 4826
rect 18694 4791 18750 4800
rect 18512 4762 18564 4768
rect 18708 4690 18736 4791
rect 18696 4684 18748 4690
rect 18696 4626 18748 4632
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 18144 4548 18196 4554
rect 18144 4490 18196 4496
rect 17972 4162 18000 4490
rect 17880 4134 18000 4162
rect 17880 3602 17908 4134
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18524 2650 18552 3334
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18708 2825 18736 2926
rect 18694 2816 18750 2825
rect 18694 2751 18750 2760
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 15016 2576 15068 2582
rect 15016 2518 15068 2524
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 16396 2576 16448 2582
rect 16396 2518 16448 2524
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 14004 2508 14056 2514
rect 14004 2450 14056 2456
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 7852 800 7880 2382
rect 9232 800 9260 2450
rect 9926 2204 10222 2224
rect 9982 2202 10006 2204
rect 10062 2202 10086 2204
rect 10142 2202 10166 2204
rect 10004 2150 10006 2202
rect 10068 2150 10080 2202
rect 10142 2150 10144 2202
rect 9982 2148 10006 2150
rect 10062 2148 10086 2150
rect 10142 2148 10166 2150
rect 9926 2128 10222 2148
rect 10612 800 10640 2450
rect 11992 800 12020 2450
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 13832 800 13860 2382
rect 15212 800 15240 2518
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 15906 2204 16202 2224
rect 15962 2202 15986 2204
rect 16042 2202 16066 2204
rect 16122 2202 16146 2204
rect 15984 2150 15986 2202
rect 16048 2150 16060 2202
rect 16122 2150 16124 2202
rect 15962 2148 15986 2150
rect 16042 2148 16066 2150
rect 16122 2148 16146 2150
rect 15906 2128 16202 2148
rect 16592 800 16620 2450
rect 17960 2372 18012 2378
rect 17960 2314 18012 2320
rect 17972 800 18000 2314
rect 19156 1420 19208 1426
rect 19156 1362 19208 1368
rect 478 0 534 800
rect 1858 0 1914 800
rect 3238 0 3294 800
rect 4618 0 4674 800
rect 5998 0 6054 800
rect 7838 0 7894 800
rect 9218 0 9274 800
rect 10598 0 10654 800
rect 11978 0 12034 800
rect 13818 0 13874 800
rect 15198 0 15254 800
rect 16578 0 16634 800
rect 17958 0 18014 800
rect 19168 785 19196 1362
rect 19154 776 19210 785
rect 19154 711 19210 720
<< via2 >>
rect 1490 20440 1546 20496
rect 6936 20154 6992 20156
rect 7016 20154 7072 20156
rect 7096 20154 7152 20156
rect 7176 20154 7232 20156
rect 6936 20102 6962 20154
rect 6962 20102 6992 20154
rect 7016 20102 7026 20154
rect 7026 20102 7072 20154
rect 7096 20102 7142 20154
rect 7142 20102 7152 20154
rect 7176 20102 7206 20154
rect 7206 20102 7232 20154
rect 6936 20100 6992 20102
rect 7016 20100 7072 20102
rect 7096 20100 7152 20102
rect 7176 20100 7232 20102
rect 12916 20154 12972 20156
rect 12996 20154 13052 20156
rect 13076 20154 13132 20156
rect 13156 20154 13212 20156
rect 12916 20102 12942 20154
rect 12942 20102 12972 20154
rect 12996 20102 13006 20154
rect 13006 20102 13052 20154
rect 13076 20102 13122 20154
rect 13122 20102 13132 20154
rect 13156 20102 13186 20154
rect 13186 20102 13212 20154
rect 12916 20100 12972 20102
rect 12996 20100 13052 20102
rect 13076 20100 13132 20102
rect 13156 20100 13212 20102
rect 18326 20440 18382 20496
rect 1398 17740 1454 17776
rect 1398 17720 1400 17740
rect 1400 17720 1452 17740
rect 1452 17720 1454 17740
rect 1398 15680 1454 15736
rect 1398 13640 1454 13696
rect 1490 11600 1546 11656
rect 1398 8900 1454 8936
rect 1398 8880 1400 8900
rect 1400 8880 1452 8900
rect 1452 8880 1454 8900
rect 1398 6860 1454 6896
rect 1398 6840 1400 6860
rect 1400 6840 1452 6860
rect 1452 6840 1454 6860
rect 3946 19610 4002 19612
rect 4026 19610 4082 19612
rect 4106 19610 4162 19612
rect 4186 19610 4242 19612
rect 3946 19558 3972 19610
rect 3972 19558 4002 19610
rect 4026 19558 4036 19610
rect 4036 19558 4082 19610
rect 4106 19558 4152 19610
rect 4152 19558 4162 19610
rect 4186 19558 4216 19610
rect 4216 19558 4242 19610
rect 3946 19556 4002 19558
rect 4026 19556 4082 19558
rect 4106 19556 4162 19558
rect 4186 19556 4242 19558
rect 3946 18522 4002 18524
rect 4026 18522 4082 18524
rect 4106 18522 4162 18524
rect 4186 18522 4242 18524
rect 3946 18470 3972 18522
rect 3972 18470 4002 18522
rect 4026 18470 4036 18522
rect 4036 18470 4082 18522
rect 4106 18470 4152 18522
rect 4152 18470 4162 18522
rect 4186 18470 4216 18522
rect 4216 18470 4242 18522
rect 3946 18468 4002 18470
rect 4026 18468 4082 18470
rect 4106 18468 4162 18470
rect 4186 18468 4242 18470
rect 3946 17434 4002 17436
rect 4026 17434 4082 17436
rect 4106 17434 4162 17436
rect 4186 17434 4242 17436
rect 3946 17382 3972 17434
rect 3972 17382 4002 17434
rect 4026 17382 4036 17434
rect 4036 17382 4082 17434
rect 4106 17382 4152 17434
rect 4152 17382 4162 17434
rect 4186 17382 4216 17434
rect 4216 17382 4242 17434
rect 3946 17380 4002 17382
rect 4026 17380 4082 17382
rect 4106 17380 4162 17382
rect 4186 17380 4242 17382
rect 3946 16346 4002 16348
rect 4026 16346 4082 16348
rect 4106 16346 4162 16348
rect 4186 16346 4242 16348
rect 3946 16294 3972 16346
rect 3972 16294 4002 16346
rect 4026 16294 4036 16346
rect 4036 16294 4082 16346
rect 4106 16294 4152 16346
rect 4152 16294 4162 16346
rect 4186 16294 4216 16346
rect 4216 16294 4242 16346
rect 3946 16292 4002 16294
rect 4026 16292 4082 16294
rect 4106 16292 4162 16294
rect 4186 16292 4242 16294
rect 3946 15258 4002 15260
rect 4026 15258 4082 15260
rect 4106 15258 4162 15260
rect 4186 15258 4242 15260
rect 3946 15206 3972 15258
rect 3972 15206 4002 15258
rect 4026 15206 4036 15258
rect 4036 15206 4082 15258
rect 4106 15206 4152 15258
rect 4152 15206 4162 15258
rect 4186 15206 4216 15258
rect 4216 15206 4242 15258
rect 3946 15204 4002 15206
rect 4026 15204 4082 15206
rect 4106 15204 4162 15206
rect 4186 15204 4242 15206
rect 3946 14170 4002 14172
rect 4026 14170 4082 14172
rect 4106 14170 4162 14172
rect 4186 14170 4242 14172
rect 3946 14118 3972 14170
rect 3972 14118 4002 14170
rect 4026 14118 4036 14170
rect 4036 14118 4082 14170
rect 4106 14118 4152 14170
rect 4152 14118 4162 14170
rect 4186 14118 4216 14170
rect 4216 14118 4242 14170
rect 3946 14116 4002 14118
rect 4026 14116 4082 14118
rect 4106 14116 4162 14118
rect 4186 14116 4242 14118
rect 3946 13082 4002 13084
rect 4026 13082 4082 13084
rect 4106 13082 4162 13084
rect 4186 13082 4242 13084
rect 3946 13030 3972 13082
rect 3972 13030 4002 13082
rect 4026 13030 4036 13082
rect 4036 13030 4082 13082
rect 4106 13030 4152 13082
rect 4152 13030 4162 13082
rect 4186 13030 4216 13082
rect 4216 13030 4242 13082
rect 3946 13028 4002 13030
rect 4026 13028 4082 13030
rect 4106 13028 4162 13030
rect 4186 13028 4242 13030
rect 3946 11994 4002 11996
rect 4026 11994 4082 11996
rect 4106 11994 4162 11996
rect 4186 11994 4242 11996
rect 3946 11942 3972 11994
rect 3972 11942 4002 11994
rect 4026 11942 4036 11994
rect 4036 11942 4082 11994
rect 4106 11942 4152 11994
rect 4152 11942 4162 11994
rect 4186 11942 4216 11994
rect 4216 11942 4242 11994
rect 3946 11940 4002 11942
rect 4026 11940 4082 11942
rect 4106 11940 4162 11942
rect 4186 11940 4242 11942
rect 3946 10906 4002 10908
rect 4026 10906 4082 10908
rect 4106 10906 4162 10908
rect 4186 10906 4242 10908
rect 3946 10854 3972 10906
rect 3972 10854 4002 10906
rect 4026 10854 4036 10906
rect 4036 10854 4082 10906
rect 4106 10854 4152 10906
rect 4152 10854 4162 10906
rect 4186 10854 4216 10906
rect 4216 10854 4242 10906
rect 3946 10852 4002 10854
rect 4026 10852 4082 10854
rect 4106 10852 4162 10854
rect 4186 10852 4242 10854
rect 1490 4820 1546 4856
rect 1490 4800 1492 4820
rect 1492 4800 1544 4820
rect 1544 4800 1546 4820
rect 1398 2760 1454 2816
rect 3946 9818 4002 9820
rect 4026 9818 4082 9820
rect 4106 9818 4162 9820
rect 4186 9818 4242 9820
rect 3946 9766 3972 9818
rect 3972 9766 4002 9818
rect 4026 9766 4036 9818
rect 4036 9766 4082 9818
rect 4106 9766 4152 9818
rect 4152 9766 4162 9818
rect 4186 9766 4216 9818
rect 4216 9766 4242 9818
rect 3946 9764 4002 9766
rect 4026 9764 4082 9766
rect 4106 9764 4162 9766
rect 4186 9764 4242 9766
rect 3946 8730 4002 8732
rect 4026 8730 4082 8732
rect 4106 8730 4162 8732
rect 4186 8730 4242 8732
rect 3946 8678 3972 8730
rect 3972 8678 4002 8730
rect 4026 8678 4036 8730
rect 4036 8678 4082 8730
rect 4106 8678 4152 8730
rect 4152 8678 4162 8730
rect 4186 8678 4216 8730
rect 4216 8678 4242 8730
rect 3946 8676 4002 8678
rect 4026 8676 4082 8678
rect 4106 8676 4162 8678
rect 4186 8676 4242 8678
rect 3946 7642 4002 7644
rect 4026 7642 4082 7644
rect 4106 7642 4162 7644
rect 4186 7642 4242 7644
rect 3946 7590 3972 7642
rect 3972 7590 4002 7642
rect 4026 7590 4036 7642
rect 4036 7590 4082 7642
rect 4106 7590 4152 7642
rect 4152 7590 4162 7642
rect 4186 7590 4216 7642
rect 4216 7590 4242 7642
rect 3946 7588 4002 7590
rect 4026 7588 4082 7590
rect 4106 7588 4162 7590
rect 4186 7588 4242 7590
rect 3946 6554 4002 6556
rect 4026 6554 4082 6556
rect 4106 6554 4162 6556
rect 4186 6554 4242 6556
rect 3946 6502 3972 6554
rect 3972 6502 4002 6554
rect 4026 6502 4036 6554
rect 4036 6502 4082 6554
rect 4106 6502 4152 6554
rect 4152 6502 4162 6554
rect 4186 6502 4216 6554
rect 4216 6502 4242 6554
rect 3946 6500 4002 6502
rect 4026 6500 4082 6502
rect 4106 6500 4162 6502
rect 4186 6500 4242 6502
rect 3946 5466 4002 5468
rect 4026 5466 4082 5468
rect 4106 5466 4162 5468
rect 4186 5466 4242 5468
rect 3946 5414 3972 5466
rect 3972 5414 4002 5466
rect 4026 5414 4036 5466
rect 4036 5414 4082 5466
rect 4106 5414 4152 5466
rect 4152 5414 4162 5466
rect 4186 5414 4216 5466
rect 4216 5414 4242 5466
rect 3946 5412 4002 5414
rect 4026 5412 4082 5414
rect 4106 5412 4162 5414
rect 4186 5412 4242 5414
rect 3946 4378 4002 4380
rect 4026 4378 4082 4380
rect 4106 4378 4162 4380
rect 4186 4378 4242 4380
rect 3946 4326 3972 4378
rect 3972 4326 4002 4378
rect 4026 4326 4036 4378
rect 4036 4326 4082 4378
rect 4106 4326 4152 4378
rect 4152 4326 4162 4378
rect 4186 4326 4216 4378
rect 4216 4326 4242 4378
rect 3946 4324 4002 4326
rect 4026 4324 4082 4326
rect 4106 4324 4162 4326
rect 4186 4324 4242 4326
rect 3946 3290 4002 3292
rect 4026 3290 4082 3292
rect 4106 3290 4162 3292
rect 4186 3290 4242 3292
rect 3946 3238 3972 3290
rect 3972 3238 4002 3290
rect 4026 3238 4036 3290
rect 4036 3238 4082 3290
rect 4106 3238 4152 3290
rect 4152 3238 4162 3290
rect 4186 3238 4216 3290
rect 4216 3238 4242 3290
rect 3946 3236 4002 3238
rect 4026 3236 4082 3238
rect 4106 3236 4162 3238
rect 4186 3236 4242 3238
rect 6936 19066 6992 19068
rect 7016 19066 7072 19068
rect 7096 19066 7152 19068
rect 7176 19066 7232 19068
rect 6936 19014 6962 19066
rect 6962 19014 6992 19066
rect 7016 19014 7026 19066
rect 7026 19014 7072 19066
rect 7096 19014 7142 19066
rect 7142 19014 7152 19066
rect 7176 19014 7206 19066
rect 7206 19014 7232 19066
rect 6936 19012 6992 19014
rect 7016 19012 7072 19014
rect 7096 19012 7152 19014
rect 7176 19012 7232 19014
rect 6936 17978 6992 17980
rect 7016 17978 7072 17980
rect 7096 17978 7152 17980
rect 7176 17978 7232 17980
rect 6936 17926 6962 17978
rect 6962 17926 6992 17978
rect 7016 17926 7026 17978
rect 7026 17926 7072 17978
rect 7096 17926 7142 17978
rect 7142 17926 7152 17978
rect 7176 17926 7206 17978
rect 7206 17926 7232 17978
rect 6936 17924 6992 17926
rect 7016 17924 7072 17926
rect 7096 17924 7152 17926
rect 7176 17924 7232 17926
rect 7930 18828 7986 18864
rect 7930 18808 7932 18828
rect 7932 18808 7984 18828
rect 7984 18808 7986 18828
rect 6936 16890 6992 16892
rect 7016 16890 7072 16892
rect 7096 16890 7152 16892
rect 7176 16890 7232 16892
rect 6936 16838 6962 16890
rect 6962 16838 6992 16890
rect 7016 16838 7026 16890
rect 7026 16838 7072 16890
rect 7096 16838 7142 16890
rect 7142 16838 7152 16890
rect 7176 16838 7206 16890
rect 7206 16838 7232 16890
rect 6936 16836 6992 16838
rect 7016 16836 7072 16838
rect 7096 16836 7152 16838
rect 7176 16836 7232 16838
rect 6936 15802 6992 15804
rect 7016 15802 7072 15804
rect 7096 15802 7152 15804
rect 7176 15802 7232 15804
rect 6936 15750 6962 15802
rect 6962 15750 6992 15802
rect 7016 15750 7026 15802
rect 7026 15750 7072 15802
rect 7096 15750 7142 15802
rect 7142 15750 7152 15802
rect 7176 15750 7206 15802
rect 7206 15750 7232 15802
rect 6936 15748 6992 15750
rect 7016 15748 7072 15750
rect 7096 15748 7152 15750
rect 7176 15748 7232 15750
rect 6936 14714 6992 14716
rect 7016 14714 7072 14716
rect 7096 14714 7152 14716
rect 7176 14714 7232 14716
rect 6936 14662 6962 14714
rect 6962 14662 6992 14714
rect 7016 14662 7026 14714
rect 7026 14662 7072 14714
rect 7096 14662 7142 14714
rect 7142 14662 7152 14714
rect 7176 14662 7206 14714
rect 7206 14662 7232 14714
rect 6936 14660 6992 14662
rect 7016 14660 7072 14662
rect 7096 14660 7152 14662
rect 7176 14660 7232 14662
rect 6936 13626 6992 13628
rect 7016 13626 7072 13628
rect 7096 13626 7152 13628
rect 7176 13626 7232 13628
rect 6936 13574 6962 13626
rect 6962 13574 6992 13626
rect 7016 13574 7026 13626
rect 7026 13574 7072 13626
rect 7096 13574 7142 13626
rect 7142 13574 7152 13626
rect 7176 13574 7206 13626
rect 7206 13574 7232 13626
rect 6936 13572 6992 13574
rect 7016 13572 7072 13574
rect 7096 13572 7152 13574
rect 7176 13572 7232 13574
rect 6936 12538 6992 12540
rect 7016 12538 7072 12540
rect 7096 12538 7152 12540
rect 7176 12538 7232 12540
rect 6936 12486 6962 12538
rect 6962 12486 6992 12538
rect 7016 12486 7026 12538
rect 7026 12486 7072 12538
rect 7096 12486 7142 12538
rect 7142 12486 7152 12538
rect 7176 12486 7206 12538
rect 7206 12486 7232 12538
rect 6936 12484 6992 12486
rect 7016 12484 7072 12486
rect 7096 12484 7152 12486
rect 7176 12484 7232 12486
rect 6936 11450 6992 11452
rect 7016 11450 7072 11452
rect 7096 11450 7152 11452
rect 7176 11450 7232 11452
rect 6936 11398 6962 11450
rect 6962 11398 6992 11450
rect 7016 11398 7026 11450
rect 7026 11398 7072 11450
rect 7096 11398 7142 11450
rect 7142 11398 7152 11450
rect 7176 11398 7206 11450
rect 7206 11398 7232 11450
rect 6936 11396 6992 11398
rect 7016 11396 7072 11398
rect 7096 11396 7152 11398
rect 7176 11396 7232 11398
rect 6936 10362 6992 10364
rect 7016 10362 7072 10364
rect 7096 10362 7152 10364
rect 7176 10362 7232 10364
rect 6936 10310 6962 10362
rect 6962 10310 6992 10362
rect 7016 10310 7026 10362
rect 7026 10310 7072 10362
rect 7096 10310 7142 10362
rect 7142 10310 7152 10362
rect 7176 10310 7206 10362
rect 7206 10310 7232 10362
rect 6936 10308 6992 10310
rect 7016 10308 7072 10310
rect 7096 10308 7152 10310
rect 7176 10308 7232 10310
rect 6936 9274 6992 9276
rect 7016 9274 7072 9276
rect 7096 9274 7152 9276
rect 7176 9274 7232 9276
rect 6936 9222 6962 9274
rect 6962 9222 6992 9274
rect 7016 9222 7026 9274
rect 7026 9222 7072 9274
rect 7096 9222 7142 9274
rect 7142 9222 7152 9274
rect 7176 9222 7206 9274
rect 7206 9222 7232 9274
rect 6936 9220 6992 9222
rect 7016 9220 7072 9222
rect 7096 9220 7152 9222
rect 7176 9220 7232 9222
rect 6936 8186 6992 8188
rect 7016 8186 7072 8188
rect 7096 8186 7152 8188
rect 7176 8186 7232 8188
rect 6936 8134 6962 8186
rect 6962 8134 6992 8186
rect 7016 8134 7026 8186
rect 7026 8134 7072 8186
rect 7096 8134 7142 8186
rect 7142 8134 7152 8186
rect 7176 8134 7206 8186
rect 7206 8134 7232 8186
rect 6936 8132 6992 8134
rect 7016 8132 7072 8134
rect 7096 8132 7152 8134
rect 7176 8132 7232 8134
rect 6936 7098 6992 7100
rect 7016 7098 7072 7100
rect 7096 7098 7152 7100
rect 7176 7098 7232 7100
rect 6936 7046 6962 7098
rect 6962 7046 6992 7098
rect 7016 7046 7026 7098
rect 7026 7046 7072 7098
rect 7096 7046 7142 7098
rect 7142 7046 7152 7098
rect 7176 7046 7206 7098
rect 7206 7046 7232 7098
rect 6936 7044 6992 7046
rect 7016 7044 7072 7046
rect 7096 7044 7152 7046
rect 7176 7044 7232 7046
rect 6936 6010 6992 6012
rect 7016 6010 7072 6012
rect 7096 6010 7152 6012
rect 7176 6010 7232 6012
rect 6936 5958 6962 6010
rect 6962 5958 6992 6010
rect 7016 5958 7026 6010
rect 7026 5958 7072 6010
rect 7096 5958 7142 6010
rect 7142 5958 7152 6010
rect 7176 5958 7206 6010
rect 7206 5958 7232 6010
rect 6936 5956 6992 5958
rect 7016 5956 7072 5958
rect 7096 5956 7152 5958
rect 7176 5956 7232 5958
rect 6936 4922 6992 4924
rect 7016 4922 7072 4924
rect 7096 4922 7152 4924
rect 7176 4922 7232 4924
rect 6936 4870 6962 4922
rect 6962 4870 6992 4922
rect 7016 4870 7026 4922
rect 7026 4870 7072 4922
rect 7096 4870 7142 4922
rect 7142 4870 7152 4922
rect 7176 4870 7206 4922
rect 7206 4870 7232 4922
rect 6936 4868 6992 4870
rect 7016 4868 7072 4870
rect 7096 4868 7152 4870
rect 7176 4868 7232 4870
rect 6936 3834 6992 3836
rect 7016 3834 7072 3836
rect 7096 3834 7152 3836
rect 7176 3834 7232 3836
rect 6936 3782 6962 3834
rect 6962 3782 6992 3834
rect 7016 3782 7026 3834
rect 7026 3782 7072 3834
rect 7096 3782 7142 3834
rect 7142 3782 7152 3834
rect 7176 3782 7206 3834
rect 7206 3782 7232 3834
rect 6936 3780 6992 3782
rect 7016 3780 7072 3782
rect 7096 3780 7152 3782
rect 7176 3780 7232 3782
rect 6936 2746 6992 2748
rect 7016 2746 7072 2748
rect 7096 2746 7152 2748
rect 7176 2746 7232 2748
rect 6936 2694 6962 2746
rect 6962 2694 6992 2746
rect 7016 2694 7026 2746
rect 7026 2694 7072 2746
rect 7096 2694 7142 2746
rect 7142 2694 7152 2746
rect 7176 2694 7206 2746
rect 7206 2694 7232 2746
rect 6936 2692 6992 2694
rect 7016 2692 7072 2694
rect 7096 2692 7152 2694
rect 7176 2692 7232 2694
rect 3946 2202 4002 2204
rect 4026 2202 4082 2204
rect 4106 2202 4162 2204
rect 4186 2202 4242 2204
rect 3946 2150 3972 2202
rect 3972 2150 4002 2202
rect 4026 2150 4036 2202
rect 4036 2150 4082 2202
rect 4106 2150 4152 2202
rect 4152 2150 4162 2202
rect 4186 2150 4216 2202
rect 4216 2150 4242 2202
rect 3946 2148 4002 2150
rect 4026 2148 4082 2150
rect 4106 2148 4162 2150
rect 4186 2148 4242 2150
rect 8574 18844 8576 18864
rect 8576 18844 8628 18864
rect 8628 18844 8630 18864
rect 8574 18808 8630 18844
rect 9926 19610 9982 19612
rect 10006 19610 10062 19612
rect 10086 19610 10142 19612
rect 10166 19610 10222 19612
rect 9926 19558 9952 19610
rect 9952 19558 9982 19610
rect 10006 19558 10016 19610
rect 10016 19558 10062 19610
rect 10086 19558 10132 19610
rect 10132 19558 10142 19610
rect 10166 19558 10196 19610
rect 10196 19558 10222 19610
rect 9926 19556 9982 19558
rect 10006 19556 10062 19558
rect 10086 19556 10142 19558
rect 10166 19556 10222 19558
rect 9926 18522 9982 18524
rect 10006 18522 10062 18524
rect 10086 18522 10142 18524
rect 10166 18522 10222 18524
rect 9926 18470 9952 18522
rect 9952 18470 9982 18522
rect 10006 18470 10016 18522
rect 10016 18470 10062 18522
rect 10086 18470 10132 18522
rect 10132 18470 10142 18522
rect 10166 18470 10196 18522
rect 10196 18470 10222 18522
rect 9926 18468 9982 18470
rect 10006 18468 10062 18470
rect 10086 18468 10142 18470
rect 10166 18468 10222 18470
rect 9926 17434 9982 17436
rect 10006 17434 10062 17436
rect 10086 17434 10142 17436
rect 10166 17434 10222 17436
rect 9926 17382 9952 17434
rect 9952 17382 9982 17434
rect 10006 17382 10016 17434
rect 10016 17382 10062 17434
rect 10086 17382 10132 17434
rect 10132 17382 10142 17434
rect 10166 17382 10196 17434
rect 10196 17382 10222 17434
rect 9926 17380 9982 17382
rect 10006 17380 10062 17382
rect 10086 17380 10142 17382
rect 10166 17380 10222 17382
rect 9926 16346 9982 16348
rect 10006 16346 10062 16348
rect 10086 16346 10142 16348
rect 10166 16346 10222 16348
rect 9926 16294 9952 16346
rect 9952 16294 9982 16346
rect 10006 16294 10016 16346
rect 10016 16294 10062 16346
rect 10086 16294 10132 16346
rect 10132 16294 10142 16346
rect 10166 16294 10196 16346
rect 10196 16294 10222 16346
rect 9926 16292 9982 16294
rect 10006 16292 10062 16294
rect 10086 16292 10142 16294
rect 10166 16292 10222 16294
rect 9926 15258 9982 15260
rect 10006 15258 10062 15260
rect 10086 15258 10142 15260
rect 10166 15258 10222 15260
rect 9926 15206 9952 15258
rect 9952 15206 9982 15258
rect 10006 15206 10016 15258
rect 10016 15206 10062 15258
rect 10086 15206 10132 15258
rect 10132 15206 10142 15258
rect 10166 15206 10196 15258
rect 10196 15206 10222 15258
rect 9926 15204 9982 15206
rect 10006 15204 10062 15206
rect 10086 15204 10142 15206
rect 10166 15204 10222 15206
rect 9926 14170 9982 14172
rect 10006 14170 10062 14172
rect 10086 14170 10142 14172
rect 10166 14170 10222 14172
rect 9926 14118 9952 14170
rect 9952 14118 9982 14170
rect 10006 14118 10016 14170
rect 10016 14118 10062 14170
rect 10086 14118 10132 14170
rect 10132 14118 10142 14170
rect 10166 14118 10196 14170
rect 10196 14118 10222 14170
rect 9926 14116 9982 14118
rect 10006 14116 10062 14118
rect 10086 14116 10142 14118
rect 10166 14116 10222 14118
rect 9926 13082 9982 13084
rect 10006 13082 10062 13084
rect 10086 13082 10142 13084
rect 10166 13082 10222 13084
rect 9926 13030 9952 13082
rect 9952 13030 9982 13082
rect 10006 13030 10016 13082
rect 10016 13030 10062 13082
rect 10086 13030 10132 13082
rect 10132 13030 10142 13082
rect 10166 13030 10196 13082
rect 10196 13030 10222 13082
rect 9926 13028 9982 13030
rect 10006 13028 10062 13030
rect 10086 13028 10142 13030
rect 10166 13028 10222 13030
rect 9926 11994 9982 11996
rect 10006 11994 10062 11996
rect 10086 11994 10142 11996
rect 10166 11994 10222 11996
rect 9926 11942 9952 11994
rect 9952 11942 9982 11994
rect 10006 11942 10016 11994
rect 10016 11942 10062 11994
rect 10086 11942 10132 11994
rect 10132 11942 10142 11994
rect 10166 11942 10196 11994
rect 10196 11942 10222 11994
rect 9926 11940 9982 11942
rect 10006 11940 10062 11942
rect 10086 11940 10142 11942
rect 10166 11940 10222 11942
rect 9926 10906 9982 10908
rect 10006 10906 10062 10908
rect 10086 10906 10142 10908
rect 10166 10906 10222 10908
rect 9926 10854 9952 10906
rect 9952 10854 9982 10906
rect 10006 10854 10016 10906
rect 10016 10854 10062 10906
rect 10086 10854 10132 10906
rect 10132 10854 10142 10906
rect 10166 10854 10196 10906
rect 10196 10854 10222 10906
rect 9926 10852 9982 10854
rect 10006 10852 10062 10854
rect 10086 10852 10142 10854
rect 10166 10852 10222 10854
rect 9926 9818 9982 9820
rect 10006 9818 10062 9820
rect 10086 9818 10142 9820
rect 10166 9818 10222 9820
rect 9926 9766 9952 9818
rect 9952 9766 9982 9818
rect 10006 9766 10016 9818
rect 10016 9766 10062 9818
rect 10086 9766 10132 9818
rect 10132 9766 10142 9818
rect 10166 9766 10196 9818
rect 10196 9766 10222 9818
rect 9926 9764 9982 9766
rect 10006 9764 10062 9766
rect 10086 9764 10142 9766
rect 10166 9764 10222 9766
rect 9926 8730 9982 8732
rect 10006 8730 10062 8732
rect 10086 8730 10142 8732
rect 10166 8730 10222 8732
rect 9926 8678 9952 8730
rect 9952 8678 9982 8730
rect 10006 8678 10016 8730
rect 10016 8678 10062 8730
rect 10086 8678 10132 8730
rect 10132 8678 10142 8730
rect 10166 8678 10196 8730
rect 10196 8678 10222 8730
rect 9926 8676 9982 8678
rect 10006 8676 10062 8678
rect 10086 8676 10142 8678
rect 10166 8676 10222 8678
rect 9926 7642 9982 7644
rect 10006 7642 10062 7644
rect 10086 7642 10142 7644
rect 10166 7642 10222 7644
rect 9926 7590 9952 7642
rect 9952 7590 9982 7642
rect 10006 7590 10016 7642
rect 10016 7590 10062 7642
rect 10086 7590 10132 7642
rect 10132 7590 10142 7642
rect 10166 7590 10196 7642
rect 10196 7590 10222 7642
rect 9926 7588 9982 7590
rect 10006 7588 10062 7590
rect 10086 7588 10142 7590
rect 10166 7588 10222 7590
rect 9926 6554 9982 6556
rect 10006 6554 10062 6556
rect 10086 6554 10142 6556
rect 10166 6554 10222 6556
rect 9926 6502 9952 6554
rect 9952 6502 9982 6554
rect 10006 6502 10016 6554
rect 10016 6502 10062 6554
rect 10086 6502 10132 6554
rect 10132 6502 10142 6554
rect 10166 6502 10196 6554
rect 10196 6502 10222 6554
rect 9926 6500 9982 6502
rect 10006 6500 10062 6502
rect 10086 6500 10142 6502
rect 10166 6500 10222 6502
rect 9926 5466 9982 5468
rect 10006 5466 10062 5468
rect 10086 5466 10142 5468
rect 10166 5466 10222 5468
rect 9926 5414 9952 5466
rect 9952 5414 9982 5466
rect 10006 5414 10016 5466
rect 10016 5414 10062 5466
rect 10086 5414 10132 5466
rect 10132 5414 10142 5466
rect 10166 5414 10196 5466
rect 10196 5414 10222 5466
rect 9926 5412 9982 5414
rect 10006 5412 10062 5414
rect 10086 5412 10142 5414
rect 10166 5412 10222 5414
rect 9926 4378 9982 4380
rect 10006 4378 10062 4380
rect 10086 4378 10142 4380
rect 10166 4378 10222 4380
rect 9926 4326 9952 4378
rect 9952 4326 9982 4378
rect 10006 4326 10016 4378
rect 10016 4326 10062 4378
rect 10086 4326 10132 4378
rect 10132 4326 10142 4378
rect 10166 4326 10196 4378
rect 10196 4326 10222 4378
rect 9926 4324 9982 4326
rect 10006 4324 10062 4326
rect 10086 4324 10142 4326
rect 10166 4324 10222 4326
rect 9926 3290 9982 3292
rect 10006 3290 10062 3292
rect 10086 3290 10142 3292
rect 10166 3290 10222 3292
rect 9926 3238 9952 3290
rect 9952 3238 9982 3290
rect 10006 3238 10016 3290
rect 10016 3238 10062 3290
rect 10086 3238 10132 3290
rect 10132 3238 10142 3290
rect 10166 3238 10196 3290
rect 10196 3238 10222 3290
rect 9926 3236 9982 3238
rect 10006 3236 10062 3238
rect 10086 3236 10142 3238
rect 10166 3236 10222 3238
rect 12916 19066 12972 19068
rect 12996 19066 13052 19068
rect 13076 19066 13132 19068
rect 13156 19066 13212 19068
rect 12916 19014 12942 19066
rect 12942 19014 12972 19066
rect 12996 19014 13006 19066
rect 13006 19014 13052 19066
rect 13076 19014 13122 19066
rect 13122 19014 13132 19066
rect 13156 19014 13186 19066
rect 13186 19014 13212 19066
rect 12916 19012 12972 19014
rect 12996 19012 13052 19014
rect 13076 19012 13132 19014
rect 13156 19012 13212 19014
rect 12916 17978 12972 17980
rect 12996 17978 13052 17980
rect 13076 17978 13132 17980
rect 13156 17978 13212 17980
rect 12916 17926 12942 17978
rect 12942 17926 12972 17978
rect 12996 17926 13006 17978
rect 13006 17926 13052 17978
rect 13076 17926 13122 17978
rect 13122 17926 13132 17978
rect 13156 17926 13186 17978
rect 13186 17926 13212 17978
rect 12916 17924 12972 17926
rect 12996 17924 13052 17926
rect 13076 17924 13132 17926
rect 13156 17924 13212 17926
rect 12916 16890 12972 16892
rect 12996 16890 13052 16892
rect 13076 16890 13132 16892
rect 13156 16890 13212 16892
rect 12916 16838 12942 16890
rect 12942 16838 12972 16890
rect 12996 16838 13006 16890
rect 13006 16838 13052 16890
rect 13076 16838 13122 16890
rect 13122 16838 13132 16890
rect 13156 16838 13186 16890
rect 13186 16838 13212 16890
rect 12916 16836 12972 16838
rect 12996 16836 13052 16838
rect 13076 16836 13132 16838
rect 13156 16836 13212 16838
rect 12916 15802 12972 15804
rect 12996 15802 13052 15804
rect 13076 15802 13132 15804
rect 13156 15802 13212 15804
rect 12916 15750 12942 15802
rect 12942 15750 12972 15802
rect 12996 15750 13006 15802
rect 13006 15750 13052 15802
rect 13076 15750 13122 15802
rect 13122 15750 13132 15802
rect 13156 15750 13186 15802
rect 13186 15750 13212 15802
rect 12916 15748 12972 15750
rect 12996 15748 13052 15750
rect 13076 15748 13132 15750
rect 13156 15748 13212 15750
rect 12916 14714 12972 14716
rect 12996 14714 13052 14716
rect 13076 14714 13132 14716
rect 13156 14714 13212 14716
rect 12916 14662 12942 14714
rect 12942 14662 12972 14714
rect 12996 14662 13006 14714
rect 13006 14662 13052 14714
rect 13076 14662 13122 14714
rect 13122 14662 13132 14714
rect 13156 14662 13186 14714
rect 13186 14662 13212 14714
rect 12916 14660 12972 14662
rect 12996 14660 13052 14662
rect 13076 14660 13132 14662
rect 13156 14660 13212 14662
rect 12916 13626 12972 13628
rect 12996 13626 13052 13628
rect 13076 13626 13132 13628
rect 13156 13626 13212 13628
rect 12916 13574 12942 13626
rect 12942 13574 12972 13626
rect 12996 13574 13006 13626
rect 13006 13574 13052 13626
rect 13076 13574 13122 13626
rect 13122 13574 13132 13626
rect 13156 13574 13186 13626
rect 13186 13574 13212 13626
rect 12916 13572 12972 13574
rect 12996 13572 13052 13574
rect 13076 13572 13132 13574
rect 13156 13572 13212 13574
rect 12916 12538 12972 12540
rect 12996 12538 13052 12540
rect 13076 12538 13132 12540
rect 13156 12538 13212 12540
rect 12916 12486 12942 12538
rect 12942 12486 12972 12538
rect 12996 12486 13006 12538
rect 13006 12486 13052 12538
rect 13076 12486 13122 12538
rect 13122 12486 13132 12538
rect 13156 12486 13186 12538
rect 13186 12486 13212 12538
rect 12916 12484 12972 12486
rect 12996 12484 13052 12486
rect 13076 12484 13132 12486
rect 13156 12484 13212 12486
rect 12916 11450 12972 11452
rect 12996 11450 13052 11452
rect 13076 11450 13132 11452
rect 13156 11450 13212 11452
rect 12916 11398 12942 11450
rect 12942 11398 12972 11450
rect 12996 11398 13006 11450
rect 13006 11398 13052 11450
rect 13076 11398 13122 11450
rect 13122 11398 13132 11450
rect 13156 11398 13186 11450
rect 13186 11398 13212 11450
rect 12916 11396 12972 11398
rect 12996 11396 13052 11398
rect 13076 11396 13132 11398
rect 13156 11396 13212 11398
rect 12916 10362 12972 10364
rect 12996 10362 13052 10364
rect 13076 10362 13132 10364
rect 13156 10362 13212 10364
rect 12916 10310 12942 10362
rect 12942 10310 12972 10362
rect 12996 10310 13006 10362
rect 13006 10310 13052 10362
rect 13076 10310 13122 10362
rect 13122 10310 13132 10362
rect 13156 10310 13186 10362
rect 13186 10310 13212 10362
rect 12916 10308 12972 10310
rect 12996 10308 13052 10310
rect 13076 10308 13132 10310
rect 13156 10308 13212 10310
rect 12916 9274 12972 9276
rect 12996 9274 13052 9276
rect 13076 9274 13132 9276
rect 13156 9274 13212 9276
rect 12916 9222 12942 9274
rect 12942 9222 12972 9274
rect 12996 9222 13006 9274
rect 13006 9222 13052 9274
rect 13076 9222 13122 9274
rect 13122 9222 13132 9274
rect 13156 9222 13186 9274
rect 13186 9222 13212 9274
rect 12916 9220 12972 9222
rect 12996 9220 13052 9222
rect 13076 9220 13132 9222
rect 13156 9220 13212 9222
rect 12916 8186 12972 8188
rect 12996 8186 13052 8188
rect 13076 8186 13132 8188
rect 13156 8186 13212 8188
rect 12916 8134 12942 8186
rect 12942 8134 12972 8186
rect 12996 8134 13006 8186
rect 13006 8134 13052 8186
rect 13076 8134 13122 8186
rect 13122 8134 13132 8186
rect 13156 8134 13186 8186
rect 13186 8134 13212 8186
rect 12916 8132 12972 8134
rect 12996 8132 13052 8134
rect 13076 8132 13132 8134
rect 13156 8132 13212 8134
rect 12916 7098 12972 7100
rect 12996 7098 13052 7100
rect 13076 7098 13132 7100
rect 13156 7098 13212 7100
rect 12916 7046 12942 7098
rect 12942 7046 12972 7098
rect 12996 7046 13006 7098
rect 13006 7046 13052 7098
rect 13076 7046 13122 7098
rect 13122 7046 13132 7098
rect 13156 7046 13186 7098
rect 13186 7046 13212 7098
rect 12916 7044 12972 7046
rect 12996 7044 13052 7046
rect 13076 7044 13132 7046
rect 13156 7044 13212 7046
rect 15906 19610 15962 19612
rect 15986 19610 16042 19612
rect 16066 19610 16122 19612
rect 16146 19610 16202 19612
rect 15906 19558 15932 19610
rect 15932 19558 15962 19610
rect 15986 19558 15996 19610
rect 15996 19558 16042 19610
rect 16066 19558 16112 19610
rect 16112 19558 16122 19610
rect 16146 19558 16176 19610
rect 16176 19558 16202 19610
rect 15906 19556 15962 19558
rect 15986 19556 16042 19558
rect 16066 19556 16122 19558
rect 16146 19556 16202 19558
rect 15906 18522 15962 18524
rect 15986 18522 16042 18524
rect 16066 18522 16122 18524
rect 16146 18522 16202 18524
rect 15906 18470 15932 18522
rect 15932 18470 15962 18522
rect 15986 18470 15996 18522
rect 15996 18470 16042 18522
rect 16066 18470 16112 18522
rect 16112 18470 16122 18522
rect 16146 18470 16176 18522
rect 16176 18470 16202 18522
rect 15906 18468 15962 18470
rect 15986 18468 16042 18470
rect 16066 18468 16122 18470
rect 16146 18468 16202 18470
rect 15906 17434 15962 17436
rect 15986 17434 16042 17436
rect 16066 17434 16122 17436
rect 16146 17434 16202 17436
rect 15906 17382 15932 17434
rect 15932 17382 15962 17434
rect 15986 17382 15996 17434
rect 15996 17382 16042 17434
rect 16066 17382 16112 17434
rect 16112 17382 16122 17434
rect 16146 17382 16176 17434
rect 16176 17382 16202 17434
rect 15906 17380 15962 17382
rect 15986 17380 16042 17382
rect 16066 17380 16122 17382
rect 16146 17380 16202 17382
rect 15906 16346 15962 16348
rect 15986 16346 16042 16348
rect 16066 16346 16122 16348
rect 16146 16346 16202 16348
rect 15906 16294 15932 16346
rect 15932 16294 15962 16346
rect 15986 16294 15996 16346
rect 15996 16294 16042 16346
rect 16066 16294 16112 16346
rect 16112 16294 16122 16346
rect 16146 16294 16176 16346
rect 16176 16294 16202 16346
rect 15906 16292 15962 16294
rect 15986 16292 16042 16294
rect 16066 16292 16122 16294
rect 16146 16292 16202 16294
rect 15906 15258 15962 15260
rect 15986 15258 16042 15260
rect 16066 15258 16122 15260
rect 16146 15258 16202 15260
rect 15906 15206 15932 15258
rect 15932 15206 15962 15258
rect 15986 15206 15996 15258
rect 15996 15206 16042 15258
rect 16066 15206 16112 15258
rect 16112 15206 16122 15258
rect 16146 15206 16176 15258
rect 16176 15206 16202 15258
rect 15906 15204 15962 15206
rect 15986 15204 16042 15206
rect 16066 15204 16122 15206
rect 16146 15204 16202 15206
rect 15906 14170 15962 14172
rect 15986 14170 16042 14172
rect 16066 14170 16122 14172
rect 16146 14170 16202 14172
rect 15906 14118 15932 14170
rect 15932 14118 15962 14170
rect 15986 14118 15996 14170
rect 15996 14118 16042 14170
rect 16066 14118 16112 14170
rect 16112 14118 16122 14170
rect 16146 14118 16176 14170
rect 16176 14118 16202 14170
rect 15906 14116 15962 14118
rect 15986 14116 16042 14118
rect 16066 14116 16122 14118
rect 16146 14116 16202 14118
rect 15906 13082 15962 13084
rect 15986 13082 16042 13084
rect 16066 13082 16122 13084
rect 16146 13082 16202 13084
rect 15906 13030 15932 13082
rect 15932 13030 15962 13082
rect 15986 13030 15996 13082
rect 15996 13030 16042 13082
rect 16066 13030 16112 13082
rect 16112 13030 16122 13082
rect 16146 13030 16176 13082
rect 16176 13030 16202 13082
rect 15906 13028 15962 13030
rect 15986 13028 16042 13030
rect 16066 13028 16122 13030
rect 16146 13028 16202 13030
rect 15906 11994 15962 11996
rect 15986 11994 16042 11996
rect 16066 11994 16122 11996
rect 16146 11994 16202 11996
rect 15906 11942 15932 11994
rect 15932 11942 15962 11994
rect 15986 11942 15996 11994
rect 15996 11942 16042 11994
rect 16066 11942 16112 11994
rect 16112 11942 16122 11994
rect 16146 11942 16176 11994
rect 16176 11942 16202 11994
rect 15906 11940 15962 11942
rect 15986 11940 16042 11942
rect 16066 11940 16122 11942
rect 16146 11940 16202 11942
rect 15906 10906 15962 10908
rect 15986 10906 16042 10908
rect 16066 10906 16122 10908
rect 16146 10906 16202 10908
rect 15906 10854 15932 10906
rect 15932 10854 15962 10906
rect 15986 10854 15996 10906
rect 15996 10854 16042 10906
rect 16066 10854 16112 10906
rect 16112 10854 16122 10906
rect 16146 10854 16176 10906
rect 16176 10854 16202 10906
rect 15906 10852 15962 10854
rect 15986 10852 16042 10854
rect 16066 10852 16122 10854
rect 16146 10852 16202 10854
rect 15906 9818 15962 9820
rect 15986 9818 16042 9820
rect 16066 9818 16122 9820
rect 16146 9818 16202 9820
rect 15906 9766 15932 9818
rect 15932 9766 15962 9818
rect 15986 9766 15996 9818
rect 15996 9766 16042 9818
rect 16066 9766 16112 9818
rect 16112 9766 16122 9818
rect 16146 9766 16176 9818
rect 16176 9766 16202 9818
rect 15906 9764 15962 9766
rect 15986 9764 16042 9766
rect 16066 9764 16122 9766
rect 16146 9764 16202 9766
rect 15906 8730 15962 8732
rect 15986 8730 16042 8732
rect 16066 8730 16122 8732
rect 16146 8730 16202 8732
rect 15906 8678 15932 8730
rect 15932 8678 15962 8730
rect 15986 8678 15996 8730
rect 15996 8678 16042 8730
rect 16066 8678 16112 8730
rect 16112 8678 16122 8730
rect 16146 8678 16176 8730
rect 16176 8678 16202 8730
rect 15906 8676 15962 8678
rect 15986 8676 16042 8678
rect 16066 8676 16122 8678
rect 16146 8676 16202 8678
rect 15906 7642 15962 7644
rect 15986 7642 16042 7644
rect 16066 7642 16122 7644
rect 16146 7642 16202 7644
rect 15906 7590 15932 7642
rect 15932 7590 15962 7642
rect 15986 7590 15996 7642
rect 15996 7590 16042 7642
rect 16066 7590 16112 7642
rect 16112 7590 16122 7642
rect 16146 7590 16176 7642
rect 16176 7590 16202 7642
rect 15906 7588 15962 7590
rect 15986 7588 16042 7590
rect 16066 7588 16122 7590
rect 16146 7588 16202 7590
rect 12916 6010 12972 6012
rect 12996 6010 13052 6012
rect 13076 6010 13132 6012
rect 13156 6010 13212 6012
rect 12916 5958 12942 6010
rect 12942 5958 12972 6010
rect 12996 5958 13006 6010
rect 13006 5958 13052 6010
rect 13076 5958 13122 6010
rect 13122 5958 13132 6010
rect 13156 5958 13186 6010
rect 13186 5958 13212 6010
rect 12916 5956 12972 5958
rect 12996 5956 13052 5958
rect 13076 5956 13132 5958
rect 13156 5956 13212 5958
rect 15906 6554 15962 6556
rect 15986 6554 16042 6556
rect 16066 6554 16122 6556
rect 16146 6554 16202 6556
rect 15906 6502 15932 6554
rect 15932 6502 15962 6554
rect 15986 6502 15996 6554
rect 15996 6502 16042 6554
rect 16066 6502 16112 6554
rect 16112 6502 16122 6554
rect 16146 6502 16176 6554
rect 16176 6502 16202 6554
rect 15906 6500 15962 6502
rect 15986 6500 16042 6502
rect 16066 6500 16122 6502
rect 16146 6500 16202 6502
rect 12916 4922 12972 4924
rect 12996 4922 13052 4924
rect 13076 4922 13132 4924
rect 13156 4922 13212 4924
rect 12916 4870 12942 4922
rect 12942 4870 12972 4922
rect 12996 4870 13006 4922
rect 13006 4870 13052 4922
rect 13076 4870 13122 4922
rect 13122 4870 13132 4922
rect 13156 4870 13186 4922
rect 13186 4870 13212 4922
rect 12916 4868 12972 4870
rect 12996 4868 13052 4870
rect 13076 4868 13132 4870
rect 13156 4868 13212 4870
rect 12916 3834 12972 3836
rect 12996 3834 13052 3836
rect 13076 3834 13132 3836
rect 13156 3834 13212 3836
rect 12916 3782 12942 3834
rect 12942 3782 12972 3834
rect 12996 3782 13006 3834
rect 13006 3782 13052 3834
rect 13076 3782 13122 3834
rect 13122 3782 13132 3834
rect 13156 3782 13186 3834
rect 13186 3782 13212 3834
rect 12916 3780 12972 3782
rect 12996 3780 13052 3782
rect 13076 3780 13132 3782
rect 13156 3780 13212 3782
rect 12916 2746 12972 2748
rect 12996 2746 13052 2748
rect 13076 2746 13132 2748
rect 13156 2746 13212 2748
rect 12916 2694 12942 2746
rect 12942 2694 12972 2746
rect 12996 2694 13006 2746
rect 13006 2694 13052 2746
rect 13076 2694 13122 2746
rect 13122 2694 13132 2746
rect 13156 2694 13186 2746
rect 13186 2694 13212 2746
rect 12916 2692 12972 2694
rect 12996 2692 13052 2694
rect 13076 2692 13132 2694
rect 13156 2692 13212 2694
rect 15906 5466 15962 5468
rect 15986 5466 16042 5468
rect 16066 5466 16122 5468
rect 16146 5466 16202 5468
rect 15906 5414 15932 5466
rect 15932 5414 15962 5466
rect 15986 5414 15996 5466
rect 15996 5414 16042 5466
rect 16066 5414 16112 5466
rect 16112 5414 16122 5466
rect 16146 5414 16176 5466
rect 16176 5414 16202 5466
rect 15906 5412 15962 5414
rect 15986 5412 16042 5414
rect 16066 5412 16122 5414
rect 16146 5412 16202 5414
rect 15906 4378 15962 4380
rect 15986 4378 16042 4380
rect 16066 4378 16122 4380
rect 16146 4378 16202 4380
rect 15906 4326 15932 4378
rect 15932 4326 15962 4378
rect 15986 4326 15996 4378
rect 15996 4326 16042 4378
rect 16066 4326 16112 4378
rect 16112 4326 16122 4378
rect 16146 4326 16176 4378
rect 16176 4326 16202 4378
rect 15906 4324 15962 4326
rect 15986 4324 16042 4326
rect 16066 4324 16122 4326
rect 16146 4324 16202 4326
rect 15906 3290 15962 3292
rect 15986 3290 16042 3292
rect 16066 3290 16122 3292
rect 16146 3290 16202 3292
rect 15906 3238 15932 3290
rect 15932 3238 15962 3290
rect 15986 3238 15996 3290
rect 15996 3238 16042 3290
rect 16066 3238 16112 3290
rect 16112 3238 16122 3290
rect 16146 3238 16176 3290
rect 16176 3238 16202 3290
rect 15906 3236 15962 3238
rect 15986 3236 16042 3238
rect 16066 3236 16122 3238
rect 16146 3236 16202 3238
rect 18694 18400 18750 18456
rect 18694 15680 18750 15736
rect 18694 13640 18750 13696
rect 18694 11636 18696 11656
rect 18696 11636 18748 11656
rect 18748 11636 18750 11656
rect 18694 11600 18750 11636
rect 18694 9560 18750 9616
rect 18694 6860 18750 6896
rect 18694 6840 18696 6860
rect 18696 6840 18748 6860
rect 18748 6840 18750 6860
rect 18694 4800 18750 4856
rect 18694 2760 18750 2816
rect 9926 2202 9982 2204
rect 10006 2202 10062 2204
rect 10086 2202 10142 2204
rect 10166 2202 10222 2204
rect 9926 2150 9952 2202
rect 9952 2150 9982 2202
rect 10006 2150 10016 2202
rect 10016 2150 10062 2202
rect 10086 2150 10132 2202
rect 10132 2150 10142 2202
rect 10166 2150 10196 2202
rect 10196 2150 10222 2202
rect 9926 2148 9982 2150
rect 10006 2148 10062 2150
rect 10086 2148 10142 2150
rect 10166 2148 10222 2150
rect 15906 2202 15962 2204
rect 15986 2202 16042 2204
rect 16066 2202 16122 2204
rect 16146 2202 16202 2204
rect 15906 2150 15932 2202
rect 15932 2150 15962 2202
rect 15986 2150 15996 2202
rect 15996 2150 16042 2202
rect 16066 2150 16112 2202
rect 16112 2150 16122 2202
rect 16146 2150 16176 2202
rect 16176 2150 16202 2202
rect 15906 2148 15962 2150
rect 15986 2148 16042 2150
rect 16066 2148 16122 2150
rect 16146 2148 16202 2150
rect 19154 720 19210 776
<< metal3 >>
rect 0 20498 800 20528
rect 1485 20498 1551 20501
rect 0 20496 1551 20498
rect 0 20440 1490 20496
rect 1546 20440 1551 20496
rect 0 20438 1551 20440
rect 0 20408 800 20438
rect 1485 20435 1551 20438
rect 18321 20498 18387 20501
rect 19396 20498 20196 20528
rect 18321 20496 20196 20498
rect 18321 20440 18326 20496
rect 18382 20440 20196 20496
rect 18321 20438 20196 20440
rect 18321 20435 18387 20438
rect 19396 20408 20196 20438
rect 6924 20160 7244 20161
rect 6924 20096 6932 20160
rect 6996 20096 7012 20160
rect 7076 20096 7092 20160
rect 7156 20096 7172 20160
rect 7236 20096 7244 20160
rect 6924 20095 7244 20096
rect 12904 20160 13224 20161
rect 12904 20096 12912 20160
rect 12976 20096 12992 20160
rect 13056 20096 13072 20160
rect 13136 20096 13152 20160
rect 13216 20096 13224 20160
rect 12904 20095 13224 20096
rect 3934 19616 4254 19617
rect 3934 19552 3942 19616
rect 4006 19552 4022 19616
rect 4086 19552 4102 19616
rect 4166 19552 4182 19616
rect 4246 19552 4254 19616
rect 3934 19551 4254 19552
rect 9914 19616 10234 19617
rect 9914 19552 9922 19616
rect 9986 19552 10002 19616
rect 10066 19552 10082 19616
rect 10146 19552 10162 19616
rect 10226 19552 10234 19616
rect 9914 19551 10234 19552
rect 15894 19616 16214 19617
rect 15894 19552 15902 19616
rect 15966 19552 15982 19616
rect 16046 19552 16062 19616
rect 16126 19552 16142 19616
rect 16206 19552 16214 19616
rect 15894 19551 16214 19552
rect 6924 19072 7244 19073
rect 6924 19008 6932 19072
rect 6996 19008 7012 19072
rect 7076 19008 7092 19072
rect 7156 19008 7172 19072
rect 7236 19008 7244 19072
rect 6924 19007 7244 19008
rect 12904 19072 13224 19073
rect 12904 19008 12912 19072
rect 12976 19008 12992 19072
rect 13056 19008 13072 19072
rect 13136 19008 13152 19072
rect 13216 19008 13224 19072
rect 12904 19007 13224 19008
rect 7925 18866 7991 18869
rect 8569 18866 8635 18869
rect 7925 18864 8635 18866
rect 7925 18808 7930 18864
rect 7986 18808 8574 18864
rect 8630 18808 8635 18864
rect 7925 18806 8635 18808
rect 7925 18803 7991 18806
rect 8569 18803 8635 18806
rect 3934 18528 4254 18529
rect 3934 18464 3942 18528
rect 4006 18464 4022 18528
rect 4086 18464 4102 18528
rect 4166 18464 4182 18528
rect 4246 18464 4254 18528
rect 3934 18463 4254 18464
rect 9914 18528 10234 18529
rect 9914 18464 9922 18528
rect 9986 18464 10002 18528
rect 10066 18464 10082 18528
rect 10146 18464 10162 18528
rect 10226 18464 10234 18528
rect 9914 18463 10234 18464
rect 15894 18528 16214 18529
rect 15894 18464 15902 18528
rect 15966 18464 15982 18528
rect 16046 18464 16062 18528
rect 16126 18464 16142 18528
rect 16206 18464 16214 18528
rect 15894 18463 16214 18464
rect 18689 18458 18755 18461
rect 19396 18458 20196 18488
rect 18689 18456 20196 18458
rect 18689 18400 18694 18456
rect 18750 18400 20196 18456
rect 18689 18398 20196 18400
rect 18689 18395 18755 18398
rect 19396 18368 20196 18398
rect 6924 17984 7244 17985
rect 6924 17920 6932 17984
rect 6996 17920 7012 17984
rect 7076 17920 7092 17984
rect 7156 17920 7172 17984
rect 7236 17920 7244 17984
rect 6924 17919 7244 17920
rect 12904 17984 13224 17985
rect 12904 17920 12912 17984
rect 12976 17920 12992 17984
rect 13056 17920 13072 17984
rect 13136 17920 13152 17984
rect 13216 17920 13224 17984
rect 12904 17919 13224 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 3934 17440 4254 17441
rect 3934 17376 3942 17440
rect 4006 17376 4022 17440
rect 4086 17376 4102 17440
rect 4166 17376 4182 17440
rect 4246 17376 4254 17440
rect 3934 17375 4254 17376
rect 9914 17440 10234 17441
rect 9914 17376 9922 17440
rect 9986 17376 10002 17440
rect 10066 17376 10082 17440
rect 10146 17376 10162 17440
rect 10226 17376 10234 17440
rect 9914 17375 10234 17376
rect 15894 17440 16214 17441
rect 15894 17376 15902 17440
rect 15966 17376 15982 17440
rect 16046 17376 16062 17440
rect 16126 17376 16142 17440
rect 16206 17376 16214 17440
rect 15894 17375 16214 17376
rect 6924 16896 7244 16897
rect 6924 16832 6932 16896
rect 6996 16832 7012 16896
rect 7076 16832 7092 16896
rect 7156 16832 7172 16896
rect 7236 16832 7244 16896
rect 6924 16831 7244 16832
rect 12904 16896 13224 16897
rect 12904 16832 12912 16896
rect 12976 16832 12992 16896
rect 13056 16832 13072 16896
rect 13136 16832 13152 16896
rect 13216 16832 13224 16896
rect 12904 16831 13224 16832
rect 3934 16352 4254 16353
rect 3934 16288 3942 16352
rect 4006 16288 4022 16352
rect 4086 16288 4102 16352
rect 4166 16288 4182 16352
rect 4246 16288 4254 16352
rect 3934 16287 4254 16288
rect 9914 16352 10234 16353
rect 9914 16288 9922 16352
rect 9986 16288 10002 16352
rect 10066 16288 10082 16352
rect 10146 16288 10162 16352
rect 10226 16288 10234 16352
rect 9914 16287 10234 16288
rect 15894 16352 16214 16353
rect 15894 16288 15902 16352
rect 15966 16288 15982 16352
rect 16046 16288 16062 16352
rect 16126 16288 16142 16352
rect 16206 16288 16214 16352
rect 15894 16287 16214 16288
rect 6924 15808 7244 15809
rect 0 15738 800 15768
rect 6924 15744 6932 15808
rect 6996 15744 7012 15808
rect 7076 15744 7092 15808
rect 7156 15744 7172 15808
rect 7236 15744 7244 15808
rect 6924 15743 7244 15744
rect 12904 15808 13224 15809
rect 12904 15744 12912 15808
rect 12976 15744 12992 15808
rect 13056 15744 13072 15808
rect 13136 15744 13152 15808
rect 13216 15744 13224 15808
rect 12904 15743 13224 15744
rect 1393 15738 1459 15741
rect 0 15736 1459 15738
rect 0 15680 1398 15736
rect 1454 15680 1459 15736
rect 0 15678 1459 15680
rect 0 15648 800 15678
rect 1393 15675 1459 15678
rect 18689 15738 18755 15741
rect 19396 15738 20196 15768
rect 18689 15736 20196 15738
rect 18689 15680 18694 15736
rect 18750 15680 20196 15736
rect 18689 15678 20196 15680
rect 18689 15675 18755 15678
rect 19396 15648 20196 15678
rect 3934 15264 4254 15265
rect 3934 15200 3942 15264
rect 4006 15200 4022 15264
rect 4086 15200 4102 15264
rect 4166 15200 4182 15264
rect 4246 15200 4254 15264
rect 3934 15199 4254 15200
rect 9914 15264 10234 15265
rect 9914 15200 9922 15264
rect 9986 15200 10002 15264
rect 10066 15200 10082 15264
rect 10146 15200 10162 15264
rect 10226 15200 10234 15264
rect 9914 15199 10234 15200
rect 15894 15264 16214 15265
rect 15894 15200 15902 15264
rect 15966 15200 15982 15264
rect 16046 15200 16062 15264
rect 16126 15200 16142 15264
rect 16206 15200 16214 15264
rect 15894 15199 16214 15200
rect 6924 14720 7244 14721
rect 6924 14656 6932 14720
rect 6996 14656 7012 14720
rect 7076 14656 7092 14720
rect 7156 14656 7172 14720
rect 7236 14656 7244 14720
rect 6924 14655 7244 14656
rect 12904 14720 13224 14721
rect 12904 14656 12912 14720
rect 12976 14656 12992 14720
rect 13056 14656 13072 14720
rect 13136 14656 13152 14720
rect 13216 14656 13224 14720
rect 12904 14655 13224 14656
rect 3934 14176 4254 14177
rect 3934 14112 3942 14176
rect 4006 14112 4022 14176
rect 4086 14112 4102 14176
rect 4166 14112 4182 14176
rect 4246 14112 4254 14176
rect 3934 14111 4254 14112
rect 9914 14176 10234 14177
rect 9914 14112 9922 14176
rect 9986 14112 10002 14176
rect 10066 14112 10082 14176
rect 10146 14112 10162 14176
rect 10226 14112 10234 14176
rect 9914 14111 10234 14112
rect 15894 14176 16214 14177
rect 15894 14112 15902 14176
rect 15966 14112 15982 14176
rect 16046 14112 16062 14176
rect 16126 14112 16142 14176
rect 16206 14112 16214 14176
rect 15894 14111 16214 14112
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 18689 13698 18755 13701
rect 19396 13698 20196 13728
rect 18689 13696 20196 13698
rect 18689 13640 18694 13696
rect 18750 13640 20196 13696
rect 18689 13638 20196 13640
rect 18689 13635 18755 13638
rect 6924 13632 7244 13633
rect 6924 13568 6932 13632
rect 6996 13568 7012 13632
rect 7076 13568 7092 13632
rect 7156 13568 7172 13632
rect 7236 13568 7244 13632
rect 6924 13567 7244 13568
rect 12904 13632 13224 13633
rect 12904 13568 12912 13632
rect 12976 13568 12992 13632
rect 13056 13568 13072 13632
rect 13136 13568 13152 13632
rect 13216 13568 13224 13632
rect 19396 13608 20196 13638
rect 12904 13567 13224 13568
rect 3934 13088 4254 13089
rect 3934 13024 3942 13088
rect 4006 13024 4022 13088
rect 4086 13024 4102 13088
rect 4166 13024 4182 13088
rect 4246 13024 4254 13088
rect 3934 13023 4254 13024
rect 9914 13088 10234 13089
rect 9914 13024 9922 13088
rect 9986 13024 10002 13088
rect 10066 13024 10082 13088
rect 10146 13024 10162 13088
rect 10226 13024 10234 13088
rect 9914 13023 10234 13024
rect 15894 13088 16214 13089
rect 15894 13024 15902 13088
rect 15966 13024 15982 13088
rect 16046 13024 16062 13088
rect 16126 13024 16142 13088
rect 16206 13024 16214 13088
rect 15894 13023 16214 13024
rect 6924 12544 7244 12545
rect 6924 12480 6932 12544
rect 6996 12480 7012 12544
rect 7076 12480 7092 12544
rect 7156 12480 7172 12544
rect 7236 12480 7244 12544
rect 6924 12479 7244 12480
rect 12904 12544 13224 12545
rect 12904 12480 12912 12544
rect 12976 12480 12992 12544
rect 13056 12480 13072 12544
rect 13136 12480 13152 12544
rect 13216 12480 13224 12544
rect 12904 12479 13224 12480
rect 3934 12000 4254 12001
rect 3934 11936 3942 12000
rect 4006 11936 4022 12000
rect 4086 11936 4102 12000
rect 4166 11936 4182 12000
rect 4246 11936 4254 12000
rect 3934 11935 4254 11936
rect 9914 12000 10234 12001
rect 9914 11936 9922 12000
rect 9986 11936 10002 12000
rect 10066 11936 10082 12000
rect 10146 11936 10162 12000
rect 10226 11936 10234 12000
rect 9914 11935 10234 11936
rect 15894 12000 16214 12001
rect 15894 11936 15902 12000
rect 15966 11936 15982 12000
rect 16046 11936 16062 12000
rect 16126 11936 16142 12000
rect 16206 11936 16214 12000
rect 15894 11935 16214 11936
rect 0 11658 800 11688
rect 1485 11658 1551 11661
rect 0 11656 1551 11658
rect 0 11600 1490 11656
rect 1546 11600 1551 11656
rect 0 11598 1551 11600
rect 0 11568 800 11598
rect 1485 11595 1551 11598
rect 18689 11658 18755 11661
rect 19396 11658 20196 11688
rect 18689 11656 20196 11658
rect 18689 11600 18694 11656
rect 18750 11600 20196 11656
rect 18689 11598 20196 11600
rect 18689 11595 18755 11598
rect 19396 11568 20196 11598
rect 6924 11456 7244 11457
rect 6924 11392 6932 11456
rect 6996 11392 7012 11456
rect 7076 11392 7092 11456
rect 7156 11392 7172 11456
rect 7236 11392 7244 11456
rect 6924 11391 7244 11392
rect 12904 11456 13224 11457
rect 12904 11392 12912 11456
rect 12976 11392 12992 11456
rect 13056 11392 13072 11456
rect 13136 11392 13152 11456
rect 13216 11392 13224 11456
rect 12904 11391 13224 11392
rect 3934 10912 4254 10913
rect 3934 10848 3942 10912
rect 4006 10848 4022 10912
rect 4086 10848 4102 10912
rect 4166 10848 4182 10912
rect 4246 10848 4254 10912
rect 3934 10847 4254 10848
rect 9914 10912 10234 10913
rect 9914 10848 9922 10912
rect 9986 10848 10002 10912
rect 10066 10848 10082 10912
rect 10146 10848 10162 10912
rect 10226 10848 10234 10912
rect 9914 10847 10234 10848
rect 15894 10912 16214 10913
rect 15894 10848 15902 10912
rect 15966 10848 15982 10912
rect 16046 10848 16062 10912
rect 16126 10848 16142 10912
rect 16206 10848 16214 10912
rect 15894 10847 16214 10848
rect 6924 10368 7244 10369
rect 6924 10304 6932 10368
rect 6996 10304 7012 10368
rect 7076 10304 7092 10368
rect 7156 10304 7172 10368
rect 7236 10304 7244 10368
rect 6924 10303 7244 10304
rect 12904 10368 13224 10369
rect 12904 10304 12912 10368
rect 12976 10304 12992 10368
rect 13056 10304 13072 10368
rect 13136 10304 13152 10368
rect 13216 10304 13224 10368
rect 12904 10303 13224 10304
rect 3934 9824 4254 9825
rect 3934 9760 3942 9824
rect 4006 9760 4022 9824
rect 4086 9760 4102 9824
rect 4166 9760 4182 9824
rect 4246 9760 4254 9824
rect 3934 9759 4254 9760
rect 9914 9824 10234 9825
rect 9914 9760 9922 9824
rect 9986 9760 10002 9824
rect 10066 9760 10082 9824
rect 10146 9760 10162 9824
rect 10226 9760 10234 9824
rect 9914 9759 10234 9760
rect 15894 9824 16214 9825
rect 15894 9760 15902 9824
rect 15966 9760 15982 9824
rect 16046 9760 16062 9824
rect 16126 9760 16142 9824
rect 16206 9760 16214 9824
rect 15894 9759 16214 9760
rect 18689 9618 18755 9621
rect 19396 9618 20196 9648
rect 18689 9616 20196 9618
rect 18689 9560 18694 9616
rect 18750 9560 20196 9616
rect 18689 9558 20196 9560
rect 18689 9555 18755 9558
rect 19396 9528 20196 9558
rect 6924 9280 7244 9281
rect 6924 9216 6932 9280
rect 6996 9216 7012 9280
rect 7076 9216 7092 9280
rect 7156 9216 7172 9280
rect 7236 9216 7244 9280
rect 6924 9215 7244 9216
rect 12904 9280 13224 9281
rect 12904 9216 12912 9280
rect 12976 9216 12992 9280
rect 13056 9216 13072 9280
rect 13136 9216 13152 9280
rect 13216 9216 13224 9280
rect 12904 9215 13224 9216
rect 0 8938 800 8968
rect 1393 8938 1459 8941
rect 0 8936 1459 8938
rect 0 8880 1398 8936
rect 1454 8880 1459 8936
rect 0 8878 1459 8880
rect 0 8848 800 8878
rect 1393 8875 1459 8878
rect 3934 8736 4254 8737
rect 3934 8672 3942 8736
rect 4006 8672 4022 8736
rect 4086 8672 4102 8736
rect 4166 8672 4182 8736
rect 4246 8672 4254 8736
rect 3934 8671 4254 8672
rect 9914 8736 10234 8737
rect 9914 8672 9922 8736
rect 9986 8672 10002 8736
rect 10066 8672 10082 8736
rect 10146 8672 10162 8736
rect 10226 8672 10234 8736
rect 9914 8671 10234 8672
rect 15894 8736 16214 8737
rect 15894 8672 15902 8736
rect 15966 8672 15982 8736
rect 16046 8672 16062 8736
rect 16126 8672 16142 8736
rect 16206 8672 16214 8736
rect 15894 8671 16214 8672
rect 6924 8192 7244 8193
rect 6924 8128 6932 8192
rect 6996 8128 7012 8192
rect 7076 8128 7092 8192
rect 7156 8128 7172 8192
rect 7236 8128 7244 8192
rect 6924 8127 7244 8128
rect 12904 8192 13224 8193
rect 12904 8128 12912 8192
rect 12976 8128 12992 8192
rect 13056 8128 13072 8192
rect 13136 8128 13152 8192
rect 13216 8128 13224 8192
rect 12904 8127 13224 8128
rect 3934 7648 4254 7649
rect 3934 7584 3942 7648
rect 4006 7584 4022 7648
rect 4086 7584 4102 7648
rect 4166 7584 4182 7648
rect 4246 7584 4254 7648
rect 3934 7583 4254 7584
rect 9914 7648 10234 7649
rect 9914 7584 9922 7648
rect 9986 7584 10002 7648
rect 10066 7584 10082 7648
rect 10146 7584 10162 7648
rect 10226 7584 10234 7648
rect 9914 7583 10234 7584
rect 15894 7648 16214 7649
rect 15894 7584 15902 7648
rect 15966 7584 15982 7648
rect 16046 7584 16062 7648
rect 16126 7584 16142 7648
rect 16206 7584 16214 7648
rect 15894 7583 16214 7584
rect 6924 7104 7244 7105
rect 6924 7040 6932 7104
rect 6996 7040 7012 7104
rect 7076 7040 7092 7104
rect 7156 7040 7172 7104
rect 7236 7040 7244 7104
rect 6924 7039 7244 7040
rect 12904 7104 13224 7105
rect 12904 7040 12912 7104
rect 12976 7040 12992 7104
rect 13056 7040 13072 7104
rect 13136 7040 13152 7104
rect 13216 7040 13224 7104
rect 12904 7039 13224 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 18689 6898 18755 6901
rect 19396 6898 20196 6928
rect 18689 6896 20196 6898
rect 18689 6840 18694 6896
rect 18750 6840 20196 6896
rect 18689 6838 20196 6840
rect 18689 6835 18755 6838
rect 19396 6808 20196 6838
rect 3934 6560 4254 6561
rect 3934 6496 3942 6560
rect 4006 6496 4022 6560
rect 4086 6496 4102 6560
rect 4166 6496 4182 6560
rect 4246 6496 4254 6560
rect 3934 6495 4254 6496
rect 9914 6560 10234 6561
rect 9914 6496 9922 6560
rect 9986 6496 10002 6560
rect 10066 6496 10082 6560
rect 10146 6496 10162 6560
rect 10226 6496 10234 6560
rect 9914 6495 10234 6496
rect 15894 6560 16214 6561
rect 15894 6496 15902 6560
rect 15966 6496 15982 6560
rect 16046 6496 16062 6560
rect 16126 6496 16142 6560
rect 16206 6496 16214 6560
rect 15894 6495 16214 6496
rect 6924 6016 7244 6017
rect 6924 5952 6932 6016
rect 6996 5952 7012 6016
rect 7076 5952 7092 6016
rect 7156 5952 7172 6016
rect 7236 5952 7244 6016
rect 6924 5951 7244 5952
rect 12904 6016 13224 6017
rect 12904 5952 12912 6016
rect 12976 5952 12992 6016
rect 13056 5952 13072 6016
rect 13136 5952 13152 6016
rect 13216 5952 13224 6016
rect 12904 5951 13224 5952
rect 3934 5472 4254 5473
rect 3934 5408 3942 5472
rect 4006 5408 4022 5472
rect 4086 5408 4102 5472
rect 4166 5408 4182 5472
rect 4246 5408 4254 5472
rect 3934 5407 4254 5408
rect 9914 5472 10234 5473
rect 9914 5408 9922 5472
rect 9986 5408 10002 5472
rect 10066 5408 10082 5472
rect 10146 5408 10162 5472
rect 10226 5408 10234 5472
rect 9914 5407 10234 5408
rect 15894 5472 16214 5473
rect 15894 5408 15902 5472
rect 15966 5408 15982 5472
rect 16046 5408 16062 5472
rect 16126 5408 16142 5472
rect 16206 5408 16214 5472
rect 15894 5407 16214 5408
rect 6924 4928 7244 4929
rect 0 4858 800 4888
rect 6924 4864 6932 4928
rect 6996 4864 7012 4928
rect 7076 4864 7092 4928
rect 7156 4864 7172 4928
rect 7236 4864 7244 4928
rect 6924 4863 7244 4864
rect 12904 4928 13224 4929
rect 12904 4864 12912 4928
rect 12976 4864 12992 4928
rect 13056 4864 13072 4928
rect 13136 4864 13152 4928
rect 13216 4864 13224 4928
rect 12904 4863 13224 4864
rect 1485 4858 1551 4861
rect 0 4856 1551 4858
rect 0 4800 1490 4856
rect 1546 4800 1551 4856
rect 0 4798 1551 4800
rect 0 4768 800 4798
rect 1485 4795 1551 4798
rect 18689 4858 18755 4861
rect 19396 4858 20196 4888
rect 18689 4856 20196 4858
rect 18689 4800 18694 4856
rect 18750 4800 20196 4856
rect 18689 4798 20196 4800
rect 18689 4795 18755 4798
rect 19396 4768 20196 4798
rect 3934 4384 4254 4385
rect 3934 4320 3942 4384
rect 4006 4320 4022 4384
rect 4086 4320 4102 4384
rect 4166 4320 4182 4384
rect 4246 4320 4254 4384
rect 3934 4319 4254 4320
rect 9914 4384 10234 4385
rect 9914 4320 9922 4384
rect 9986 4320 10002 4384
rect 10066 4320 10082 4384
rect 10146 4320 10162 4384
rect 10226 4320 10234 4384
rect 9914 4319 10234 4320
rect 15894 4384 16214 4385
rect 15894 4320 15902 4384
rect 15966 4320 15982 4384
rect 16046 4320 16062 4384
rect 16126 4320 16142 4384
rect 16206 4320 16214 4384
rect 15894 4319 16214 4320
rect 6924 3840 7244 3841
rect 6924 3776 6932 3840
rect 6996 3776 7012 3840
rect 7076 3776 7092 3840
rect 7156 3776 7172 3840
rect 7236 3776 7244 3840
rect 6924 3775 7244 3776
rect 12904 3840 13224 3841
rect 12904 3776 12912 3840
rect 12976 3776 12992 3840
rect 13056 3776 13072 3840
rect 13136 3776 13152 3840
rect 13216 3776 13224 3840
rect 12904 3775 13224 3776
rect 3934 3296 4254 3297
rect 3934 3232 3942 3296
rect 4006 3232 4022 3296
rect 4086 3232 4102 3296
rect 4166 3232 4182 3296
rect 4246 3232 4254 3296
rect 3934 3231 4254 3232
rect 9914 3296 10234 3297
rect 9914 3232 9922 3296
rect 9986 3232 10002 3296
rect 10066 3232 10082 3296
rect 10146 3232 10162 3296
rect 10226 3232 10234 3296
rect 9914 3231 10234 3232
rect 15894 3296 16214 3297
rect 15894 3232 15902 3296
rect 15966 3232 15982 3296
rect 16046 3232 16062 3296
rect 16126 3232 16142 3296
rect 16206 3232 16214 3296
rect 15894 3231 16214 3232
rect 0 2818 800 2848
rect 1393 2818 1459 2821
rect 0 2816 1459 2818
rect 0 2760 1398 2816
rect 1454 2760 1459 2816
rect 0 2758 1459 2760
rect 0 2728 800 2758
rect 1393 2755 1459 2758
rect 18689 2818 18755 2821
rect 19396 2818 20196 2848
rect 18689 2816 20196 2818
rect 18689 2760 18694 2816
rect 18750 2760 20196 2816
rect 18689 2758 20196 2760
rect 18689 2755 18755 2758
rect 6924 2752 7244 2753
rect 6924 2688 6932 2752
rect 6996 2688 7012 2752
rect 7076 2688 7092 2752
rect 7156 2688 7172 2752
rect 7236 2688 7244 2752
rect 6924 2687 7244 2688
rect 12904 2752 13224 2753
rect 12904 2688 12912 2752
rect 12976 2688 12992 2752
rect 13056 2688 13072 2752
rect 13136 2688 13152 2752
rect 13216 2688 13224 2752
rect 19396 2728 20196 2758
rect 12904 2687 13224 2688
rect 3934 2208 4254 2209
rect 3934 2144 3942 2208
rect 4006 2144 4022 2208
rect 4086 2144 4102 2208
rect 4166 2144 4182 2208
rect 4246 2144 4254 2208
rect 3934 2143 4254 2144
rect 9914 2208 10234 2209
rect 9914 2144 9922 2208
rect 9986 2144 10002 2208
rect 10066 2144 10082 2208
rect 10146 2144 10162 2208
rect 10226 2144 10234 2208
rect 9914 2143 10234 2144
rect 15894 2208 16214 2209
rect 15894 2144 15902 2208
rect 15966 2144 15982 2208
rect 16046 2144 16062 2208
rect 16126 2144 16142 2208
rect 16206 2144 16214 2208
rect 15894 2143 16214 2144
rect 19149 778 19215 781
rect 19396 778 20196 808
rect 19149 776 20196 778
rect 19149 720 19154 776
rect 19210 720 20196 776
rect 19149 718 20196 720
rect 19149 715 19215 718
rect 19396 688 20196 718
<< via3 >>
rect 6932 20156 6996 20160
rect 6932 20100 6936 20156
rect 6936 20100 6992 20156
rect 6992 20100 6996 20156
rect 6932 20096 6996 20100
rect 7012 20156 7076 20160
rect 7012 20100 7016 20156
rect 7016 20100 7072 20156
rect 7072 20100 7076 20156
rect 7012 20096 7076 20100
rect 7092 20156 7156 20160
rect 7092 20100 7096 20156
rect 7096 20100 7152 20156
rect 7152 20100 7156 20156
rect 7092 20096 7156 20100
rect 7172 20156 7236 20160
rect 7172 20100 7176 20156
rect 7176 20100 7232 20156
rect 7232 20100 7236 20156
rect 7172 20096 7236 20100
rect 12912 20156 12976 20160
rect 12912 20100 12916 20156
rect 12916 20100 12972 20156
rect 12972 20100 12976 20156
rect 12912 20096 12976 20100
rect 12992 20156 13056 20160
rect 12992 20100 12996 20156
rect 12996 20100 13052 20156
rect 13052 20100 13056 20156
rect 12992 20096 13056 20100
rect 13072 20156 13136 20160
rect 13072 20100 13076 20156
rect 13076 20100 13132 20156
rect 13132 20100 13136 20156
rect 13072 20096 13136 20100
rect 13152 20156 13216 20160
rect 13152 20100 13156 20156
rect 13156 20100 13212 20156
rect 13212 20100 13216 20156
rect 13152 20096 13216 20100
rect 3942 19612 4006 19616
rect 3942 19556 3946 19612
rect 3946 19556 4002 19612
rect 4002 19556 4006 19612
rect 3942 19552 4006 19556
rect 4022 19612 4086 19616
rect 4022 19556 4026 19612
rect 4026 19556 4082 19612
rect 4082 19556 4086 19612
rect 4022 19552 4086 19556
rect 4102 19612 4166 19616
rect 4102 19556 4106 19612
rect 4106 19556 4162 19612
rect 4162 19556 4166 19612
rect 4102 19552 4166 19556
rect 4182 19612 4246 19616
rect 4182 19556 4186 19612
rect 4186 19556 4242 19612
rect 4242 19556 4246 19612
rect 4182 19552 4246 19556
rect 9922 19612 9986 19616
rect 9922 19556 9926 19612
rect 9926 19556 9982 19612
rect 9982 19556 9986 19612
rect 9922 19552 9986 19556
rect 10002 19612 10066 19616
rect 10002 19556 10006 19612
rect 10006 19556 10062 19612
rect 10062 19556 10066 19612
rect 10002 19552 10066 19556
rect 10082 19612 10146 19616
rect 10082 19556 10086 19612
rect 10086 19556 10142 19612
rect 10142 19556 10146 19612
rect 10082 19552 10146 19556
rect 10162 19612 10226 19616
rect 10162 19556 10166 19612
rect 10166 19556 10222 19612
rect 10222 19556 10226 19612
rect 10162 19552 10226 19556
rect 15902 19612 15966 19616
rect 15902 19556 15906 19612
rect 15906 19556 15962 19612
rect 15962 19556 15966 19612
rect 15902 19552 15966 19556
rect 15982 19612 16046 19616
rect 15982 19556 15986 19612
rect 15986 19556 16042 19612
rect 16042 19556 16046 19612
rect 15982 19552 16046 19556
rect 16062 19612 16126 19616
rect 16062 19556 16066 19612
rect 16066 19556 16122 19612
rect 16122 19556 16126 19612
rect 16062 19552 16126 19556
rect 16142 19612 16206 19616
rect 16142 19556 16146 19612
rect 16146 19556 16202 19612
rect 16202 19556 16206 19612
rect 16142 19552 16206 19556
rect 6932 19068 6996 19072
rect 6932 19012 6936 19068
rect 6936 19012 6992 19068
rect 6992 19012 6996 19068
rect 6932 19008 6996 19012
rect 7012 19068 7076 19072
rect 7012 19012 7016 19068
rect 7016 19012 7072 19068
rect 7072 19012 7076 19068
rect 7012 19008 7076 19012
rect 7092 19068 7156 19072
rect 7092 19012 7096 19068
rect 7096 19012 7152 19068
rect 7152 19012 7156 19068
rect 7092 19008 7156 19012
rect 7172 19068 7236 19072
rect 7172 19012 7176 19068
rect 7176 19012 7232 19068
rect 7232 19012 7236 19068
rect 7172 19008 7236 19012
rect 12912 19068 12976 19072
rect 12912 19012 12916 19068
rect 12916 19012 12972 19068
rect 12972 19012 12976 19068
rect 12912 19008 12976 19012
rect 12992 19068 13056 19072
rect 12992 19012 12996 19068
rect 12996 19012 13052 19068
rect 13052 19012 13056 19068
rect 12992 19008 13056 19012
rect 13072 19068 13136 19072
rect 13072 19012 13076 19068
rect 13076 19012 13132 19068
rect 13132 19012 13136 19068
rect 13072 19008 13136 19012
rect 13152 19068 13216 19072
rect 13152 19012 13156 19068
rect 13156 19012 13212 19068
rect 13212 19012 13216 19068
rect 13152 19008 13216 19012
rect 3942 18524 4006 18528
rect 3942 18468 3946 18524
rect 3946 18468 4002 18524
rect 4002 18468 4006 18524
rect 3942 18464 4006 18468
rect 4022 18524 4086 18528
rect 4022 18468 4026 18524
rect 4026 18468 4082 18524
rect 4082 18468 4086 18524
rect 4022 18464 4086 18468
rect 4102 18524 4166 18528
rect 4102 18468 4106 18524
rect 4106 18468 4162 18524
rect 4162 18468 4166 18524
rect 4102 18464 4166 18468
rect 4182 18524 4246 18528
rect 4182 18468 4186 18524
rect 4186 18468 4242 18524
rect 4242 18468 4246 18524
rect 4182 18464 4246 18468
rect 9922 18524 9986 18528
rect 9922 18468 9926 18524
rect 9926 18468 9982 18524
rect 9982 18468 9986 18524
rect 9922 18464 9986 18468
rect 10002 18524 10066 18528
rect 10002 18468 10006 18524
rect 10006 18468 10062 18524
rect 10062 18468 10066 18524
rect 10002 18464 10066 18468
rect 10082 18524 10146 18528
rect 10082 18468 10086 18524
rect 10086 18468 10142 18524
rect 10142 18468 10146 18524
rect 10082 18464 10146 18468
rect 10162 18524 10226 18528
rect 10162 18468 10166 18524
rect 10166 18468 10222 18524
rect 10222 18468 10226 18524
rect 10162 18464 10226 18468
rect 15902 18524 15966 18528
rect 15902 18468 15906 18524
rect 15906 18468 15962 18524
rect 15962 18468 15966 18524
rect 15902 18464 15966 18468
rect 15982 18524 16046 18528
rect 15982 18468 15986 18524
rect 15986 18468 16042 18524
rect 16042 18468 16046 18524
rect 15982 18464 16046 18468
rect 16062 18524 16126 18528
rect 16062 18468 16066 18524
rect 16066 18468 16122 18524
rect 16122 18468 16126 18524
rect 16062 18464 16126 18468
rect 16142 18524 16206 18528
rect 16142 18468 16146 18524
rect 16146 18468 16202 18524
rect 16202 18468 16206 18524
rect 16142 18464 16206 18468
rect 6932 17980 6996 17984
rect 6932 17924 6936 17980
rect 6936 17924 6992 17980
rect 6992 17924 6996 17980
rect 6932 17920 6996 17924
rect 7012 17980 7076 17984
rect 7012 17924 7016 17980
rect 7016 17924 7072 17980
rect 7072 17924 7076 17980
rect 7012 17920 7076 17924
rect 7092 17980 7156 17984
rect 7092 17924 7096 17980
rect 7096 17924 7152 17980
rect 7152 17924 7156 17980
rect 7092 17920 7156 17924
rect 7172 17980 7236 17984
rect 7172 17924 7176 17980
rect 7176 17924 7232 17980
rect 7232 17924 7236 17980
rect 7172 17920 7236 17924
rect 12912 17980 12976 17984
rect 12912 17924 12916 17980
rect 12916 17924 12972 17980
rect 12972 17924 12976 17980
rect 12912 17920 12976 17924
rect 12992 17980 13056 17984
rect 12992 17924 12996 17980
rect 12996 17924 13052 17980
rect 13052 17924 13056 17980
rect 12992 17920 13056 17924
rect 13072 17980 13136 17984
rect 13072 17924 13076 17980
rect 13076 17924 13132 17980
rect 13132 17924 13136 17980
rect 13072 17920 13136 17924
rect 13152 17980 13216 17984
rect 13152 17924 13156 17980
rect 13156 17924 13212 17980
rect 13212 17924 13216 17980
rect 13152 17920 13216 17924
rect 3942 17436 4006 17440
rect 3942 17380 3946 17436
rect 3946 17380 4002 17436
rect 4002 17380 4006 17436
rect 3942 17376 4006 17380
rect 4022 17436 4086 17440
rect 4022 17380 4026 17436
rect 4026 17380 4082 17436
rect 4082 17380 4086 17436
rect 4022 17376 4086 17380
rect 4102 17436 4166 17440
rect 4102 17380 4106 17436
rect 4106 17380 4162 17436
rect 4162 17380 4166 17436
rect 4102 17376 4166 17380
rect 4182 17436 4246 17440
rect 4182 17380 4186 17436
rect 4186 17380 4242 17436
rect 4242 17380 4246 17436
rect 4182 17376 4246 17380
rect 9922 17436 9986 17440
rect 9922 17380 9926 17436
rect 9926 17380 9982 17436
rect 9982 17380 9986 17436
rect 9922 17376 9986 17380
rect 10002 17436 10066 17440
rect 10002 17380 10006 17436
rect 10006 17380 10062 17436
rect 10062 17380 10066 17436
rect 10002 17376 10066 17380
rect 10082 17436 10146 17440
rect 10082 17380 10086 17436
rect 10086 17380 10142 17436
rect 10142 17380 10146 17436
rect 10082 17376 10146 17380
rect 10162 17436 10226 17440
rect 10162 17380 10166 17436
rect 10166 17380 10222 17436
rect 10222 17380 10226 17436
rect 10162 17376 10226 17380
rect 15902 17436 15966 17440
rect 15902 17380 15906 17436
rect 15906 17380 15962 17436
rect 15962 17380 15966 17436
rect 15902 17376 15966 17380
rect 15982 17436 16046 17440
rect 15982 17380 15986 17436
rect 15986 17380 16042 17436
rect 16042 17380 16046 17436
rect 15982 17376 16046 17380
rect 16062 17436 16126 17440
rect 16062 17380 16066 17436
rect 16066 17380 16122 17436
rect 16122 17380 16126 17436
rect 16062 17376 16126 17380
rect 16142 17436 16206 17440
rect 16142 17380 16146 17436
rect 16146 17380 16202 17436
rect 16202 17380 16206 17436
rect 16142 17376 16206 17380
rect 6932 16892 6996 16896
rect 6932 16836 6936 16892
rect 6936 16836 6992 16892
rect 6992 16836 6996 16892
rect 6932 16832 6996 16836
rect 7012 16892 7076 16896
rect 7012 16836 7016 16892
rect 7016 16836 7072 16892
rect 7072 16836 7076 16892
rect 7012 16832 7076 16836
rect 7092 16892 7156 16896
rect 7092 16836 7096 16892
rect 7096 16836 7152 16892
rect 7152 16836 7156 16892
rect 7092 16832 7156 16836
rect 7172 16892 7236 16896
rect 7172 16836 7176 16892
rect 7176 16836 7232 16892
rect 7232 16836 7236 16892
rect 7172 16832 7236 16836
rect 12912 16892 12976 16896
rect 12912 16836 12916 16892
rect 12916 16836 12972 16892
rect 12972 16836 12976 16892
rect 12912 16832 12976 16836
rect 12992 16892 13056 16896
rect 12992 16836 12996 16892
rect 12996 16836 13052 16892
rect 13052 16836 13056 16892
rect 12992 16832 13056 16836
rect 13072 16892 13136 16896
rect 13072 16836 13076 16892
rect 13076 16836 13132 16892
rect 13132 16836 13136 16892
rect 13072 16832 13136 16836
rect 13152 16892 13216 16896
rect 13152 16836 13156 16892
rect 13156 16836 13212 16892
rect 13212 16836 13216 16892
rect 13152 16832 13216 16836
rect 3942 16348 4006 16352
rect 3942 16292 3946 16348
rect 3946 16292 4002 16348
rect 4002 16292 4006 16348
rect 3942 16288 4006 16292
rect 4022 16348 4086 16352
rect 4022 16292 4026 16348
rect 4026 16292 4082 16348
rect 4082 16292 4086 16348
rect 4022 16288 4086 16292
rect 4102 16348 4166 16352
rect 4102 16292 4106 16348
rect 4106 16292 4162 16348
rect 4162 16292 4166 16348
rect 4102 16288 4166 16292
rect 4182 16348 4246 16352
rect 4182 16292 4186 16348
rect 4186 16292 4242 16348
rect 4242 16292 4246 16348
rect 4182 16288 4246 16292
rect 9922 16348 9986 16352
rect 9922 16292 9926 16348
rect 9926 16292 9982 16348
rect 9982 16292 9986 16348
rect 9922 16288 9986 16292
rect 10002 16348 10066 16352
rect 10002 16292 10006 16348
rect 10006 16292 10062 16348
rect 10062 16292 10066 16348
rect 10002 16288 10066 16292
rect 10082 16348 10146 16352
rect 10082 16292 10086 16348
rect 10086 16292 10142 16348
rect 10142 16292 10146 16348
rect 10082 16288 10146 16292
rect 10162 16348 10226 16352
rect 10162 16292 10166 16348
rect 10166 16292 10222 16348
rect 10222 16292 10226 16348
rect 10162 16288 10226 16292
rect 15902 16348 15966 16352
rect 15902 16292 15906 16348
rect 15906 16292 15962 16348
rect 15962 16292 15966 16348
rect 15902 16288 15966 16292
rect 15982 16348 16046 16352
rect 15982 16292 15986 16348
rect 15986 16292 16042 16348
rect 16042 16292 16046 16348
rect 15982 16288 16046 16292
rect 16062 16348 16126 16352
rect 16062 16292 16066 16348
rect 16066 16292 16122 16348
rect 16122 16292 16126 16348
rect 16062 16288 16126 16292
rect 16142 16348 16206 16352
rect 16142 16292 16146 16348
rect 16146 16292 16202 16348
rect 16202 16292 16206 16348
rect 16142 16288 16206 16292
rect 6932 15804 6996 15808
rect 6932 15748 6936 15804
rect 6936 15748 6992 15804
rect 6992 15748 6996 15804
rect 6932 15744 6996 15748
rect 7012 15804 7076 15808
rect 7012 15748 7016 15804
rect 7016 15748 7072 15804
rect 7072 15748 7076 15804
rect 7012 15744 7076 15748
rect 7092 15804 7156 15808
rect 7092 15748 7096 15804
rect 7096 15748 7152 15804
rect 7152 15748 7156 15804
rect 7092 15744 7156 15748
rect 7172 15804 7236 15808
rect 7172 15748 7176 15804
rect 7176 15748 7232 15804
rect 7232 15748 7236 15804
rect 7172 15744 7236 15748
rect 12912 15804 12976 15808
rect 12912 15748 12916 15804
rect 12916 15748 12972 15804
rect 12972 15748 12976 15804
rect 12912 15744 12976 15748
rect 12992 15804 13056 15808
rect 12992 15748 12996 15804
rect 12996 15748 13052 15804
rect 13052 15748 13056 15804
rect 12992 15744 13056 15748
rect 13072 15804 13136 15808
rect 13072 15748 13076 15804
rect 13076 15748 13132 15804
rect 13132 15748 13136 15804
rect 13072 15744 13136 15748
rect 13152 15804 13216 15808
rect 13152 15748 13156 15804
rect 13156 15748 13212 15804
rect 13212 15748 13216 15804
rect 13152 15744 13216 15748
rect 3942 15260 4006 15264
rect 3942 15204 3946 15260
rect 3946 15204 4002 15260
rect 4002 15204 4006 15260
rect 3942 15200 4006 15204
rect 4022 15260 4086 15264
rect 4022 15204 4026 15260
rect 4026 15204 4082 15260
rect 4082 15204 4086 15260
rect 4022 15200 4086 15204
rect 4102 15260 4166 15264
rect 4102 15204 4106 15260
rect 4106 15204 4162 15260
rect 4162 15204 4166 15260
rect 4102 15200 4166 15204
rect 4182 15260 4246 15264
rect 4182 15204 4186 15260
rect 4186 15204 4242 15260
rect 4242 15204 4246 15260
rect 4182 15200 4246 15204
rect 9922 15260 9986 15264
rect 9922 15204 9926 15260
rect 9926 15204 9982 15260
rect 9982 15204 9986 15260
rect 9922 15200 9986 15204
rect 10002 15260 10066 15264
rect 10002 15204 10006 15260
rect 10006 15204 10062 15260
rect 10062 15204 10066 15260
rect 10002 15200 10066 15204
rect 10082 15260 10146 15264
rect 10082 15204 10086 15260
rect 10086 15204 10142 15260
rect 10142 15204 10146 15260
rect 10082 15200 10146 15204
rect 10162 15260 10226 15264
rect 10162 15204 10166 15260
rect 10166 15204 10222 15260
rect 10222 15204 10226 15260
rect 10162 15200 10226 15204
rect 15902 15260 15966 15264
rect 15902 15204 15906 15260
rect 15906 15204 15962 15260
rect 15962 15204 15966 15260
rect 15902 15200 15966 15204
rect 15982 15260 16046 15264
rect 15982 15204 15986 15260
rect 15986 15204 16042 15260
rect 16042 15204 16046 15260
rect 15982 15200 16046 15204
rect 16062 15260 16126 15264
rect 16062 15204 16066 15260
rect 16066 15204 16122 15260
rect 16122 15204 16126 15260
rect 16062 15200 16126 15204
rect 16142 15260 16206 15264
rect 16142 15204 16146 15260
rect 16146 15204 16202 15260
rect 16202 15204 16206 15260
rect 16142 15200 16206 15204
rect 6932 14716 6996 14720
rect 6932 14660 6936 14716
rect 6936 14660 6992 14716
rect 6992 14660 6996 14716
rect 6932 14656 6996 14660
rect 7012 14716 7076 14720
rect 7012 14660 7016 14716
rect 7016 14660 7072 14716
rect 7072 14660 7076 14716
rect 7012 14656 7076 14660
rect 7092 14716 7156 14720
rect 7092 14660 7096 14716
rect 7096 14660 7152 14716
rect 7152 14660 7156 14716
rect 7092 14656 7156 14660
rect 7172 14716 7236 14720
rect 7172 14660 7176 14716
rect 7176 14660 7232 14716
rect 7232 14660 7236 14716
rect 7172 14656 7236 14660
rect 12912 14716 12976 14720
rect 12912 14660 12916 14716
rect 12916 14660 12972 14716
rect 12972 14660 12976 14716
rect 12912 14656 12976 14660
rect 12992 14716 13056 14720
rect 12992 14660 12996 14716
rect 12996 14660 13052 14716
rect 13052 14660 13056 14716
rect 12992 14656 13056 14660
rect 13072 14716 13136 14720
rect 13072 14660 13076 14716
rect 13076 14660 13132 14716
rect 13132 14660 13136 14716
rect 13072 14656 13136 14660
rect 13152 14716 13216 14720
rect 13152 14660 13156 14716
rect 13156 14660 13212 14716
rect 13212 14660 13216 14716
rect 13152 14656 13216 14660
rect 3942 14172 4006 14176
rect 3942 14116 3946 14172
rect 3946 14116 4002 14172
rect 4002 14116 4006 14172
rect 3942 14112 4006 14116
rect 4022 14172 4086 14176
rect 4022 14116 4026 14172
rect 4026 14116 4082 14172
rect 4082 14116 4086 14172
rect 4022 14112 4086 14116
rect 4102 14172 4166 14176
rect 4102 14116 4106 14172
rect 4106 14116 4162 14172
rect 4162 14116 4166 14172
rect 4102 14112 4166 14116
rect 4182 14172 4246 14176
rect 4182 14116 4186 14172
rect 4186 14116 4242 14172
rect 4242 14116 4246 14172
rect 4182 14112 4246 14116
rect 9922 14172 9986 14176
rect 9922 14116 9926 14172
rect 9926 14116 9982 14172
rect 9982 14116 9986 14172
rect 9922 14112 9986 14116
rect 10002 14172 10066 14176
rect 10002 14116 10006 14172
rect 10006 14116 10062 14172
rect 10062 14116 10066 14172
rect 10002 14112 10066 14116
rect 10082 14172 10146 14176
rect 10082 14116 10086 14172
rect 10086 14116 10142 14172
rect 10142 14116 10146 14172
rect 10082 14112 10146 14116
rect 10162 14172 10226 14176
rect 10162 14116 10166 14172
rect 10166 14116 10222 14172
rect 10222 14116 10226 14172
rect 10162 14112 10226 14116
rect 15902 14172 15966 14176
rect 15902 14116 15906 14172
rect 15906 14116 15962 14172
rect 15962 14116 15966 14172
rect 15902 14112 15966 14116
rect 15982 14172 16046 14176
rect 15982 14116 15986 14172
rect 15986 14116 16042 14172
rect 16042 14116 16046 14172
rect 15982 14112 16046 14116
rect 16062 14172 16126 14176
rect 16062 14116 16066 14172
rect 16066 14116 16122 14172
rect 16122 14116 16126 14172
rect 16062 14112 16126 14116
rect 16142 14172 16206 14176
rect 16142 14116 16146 14172
rect 16146 14116 16202 14172
rect 16202 14116 16206 14172
rect 16142 14112 16206 14116
rect 6932 13628 6996 13632
rect 6932 13572 6936 13628
rect 6936 13572 6992 13628
rect 6992 13572 6996 13628
rect 6932 13568 6996 13572
rect 7012 13628 7076 13632
rect 7012 13572 7016 13628
rect 7016 13572 7072 13628
rect 7072 13572 7076 13628
rect 7012 13568 7076 13572
rect 7092 13628 7156 13632
rect 7092 13572 7096 13628
rect 7096 13572 7152 13628
rect 7152 13572 7156 13628
rect 7092 13568 7156 13572
rect 7172 13628 7236 13632
rect 7172 13572 7176 13628
rect 7176 13572 7232 13628
rect 7232 13572 7236 13628
rect 7172 13568 7236 13572
rect 12912 13628 12976 13632
rect 12912 13572 12916 13628
rect 12916 13572 12972 13628
rect 12972 13572 12976 13628
rect 12912 13568 12976 13572
rect 12992 13628 13056 13632
rect 12992 13572 12996 13628
rect 12996 13572 13052 13628
rect 13052 13572 13056 13628
rect 12992 13568 13056 13572
rect 13072 13628 13136 13632
rect 13072 13572 13076 13628
rect 13076 13572 13132 13628
rect 13132 13572 13136 13628
rect 13072 13568 13136 13572
rect 13152 13628 13216 13632
rect 13152 13572 13156 13628
rect 13156 13572 13212 13628
rect 13212 13572 13216 13628
rect 13152 13568 13216 13572
rect 3942 13084 4006 13088
rect 3942 13028 3946 13084
rect 3946 13028 4002 13084
rect 4002 13028 4006 13084
rect 3942 13024 4006 13028
rect 4022 13084 4086 13088
rect 4022 13028 4026 13084
rect 4026 13028 4082 13084
rect 4082 13028 4086 13084
rect 4022 13024 4086 13028
rect 4102 13084 4166 13088
rect 4102 13028 4106 13084
rect 4106 13028 4162 13084
rect 4162 13028 4166 13084
rect 4102 13024 4166 13028
rect 4182 13084 4246 13088
rect 4182 13028 4186 13084
rect 4186 13028 4242 13084
rect 4242 13028 4246 13084
rect 4182 13024 4246 13028
rect 9922 13084 9986 13088
rect 9922 13028 9926 13084
rect 9926 13028 9982 13084
rect 9982 13028 9986 13084
rect 9922 13024 9986 13028
rect 10002 13084 10066 13088
rect 10002 13028 10006 13084
rect 10006 13028 10062 13084
rect 10062 13028 10066 13084
rect 10002 13024 10066 13028
rect 10082 13084 10146 13088
rect 10082 13028 10086 13084
rect 10086 13028 10142 13084
rect 10142 13028 10146 13084
rect 10082 13024 10146 13028
rect 10162 13084 10226 13088
rect 10162 13028 10166 13084
rect 10166 13028 10222 13084
rect 10222 13028 10226 13084
rect 10162 13024 10226 13028
rect 15902 13084 15966 13088
rect 15902 13028 15906 13084
rect 15906 13028 15962 13084
rect 15962 13028 15966 13084
rect 15902 13024 15966 13028
rect 15982 13084 16046 13088
rect 15982 13028 15986 13084
rect 15986 13028 16042 13084
rect 16042 13028 16046 13084
rect 15982 13024 16046 13028
rect 16062 13084 16126 13088
rect 16062 13028 16066 13084
rect 16066 13028 16122 13084
rect 16122 13028 16126 13084
rect 16062 13024 16126 13028
rect 16142 13084 16206 13088
rect 16142 13028 16146 13084
rect 16146 13028 16202 13084
rect 16202 13028 16206 13084
rect 16142 13024 16206 13028
rect 6932 12540 6996 12544
rect 6932 12484 6936 12540
rect 6936 12484 6992 12540
rect 6992 12484 6996 12540
rect 6932 12480 6996 12484
rect 7012 12540 7076 12544
rect 7012 12484 7016 12540
rect 7016 12484 7072 12540
rect 7072 12484 7076 12540
rect 7012 12480 7076 12484
rect 7092 12540 7156 12544
rect 7092 12484 7096 12540
rect 7096 12484 7152 12540
rect 7152 12484 7156 12540
rect 7092 12480 7156 12484
rect 7172 12540 7236 12544
rect 7172 12484 7176 12540
rect 7176 12484 7232 12540
rect 7232 12484 7236 12540
rect 7172 12480 7236 12484
rect 12912 12540 12976 12544
rect 12912 12484 12916 12540
rect 12916 12484 12972 12540
rect 12972 12484 12976 12540
rect 12912 12480 12976 12484
rect 12992 12540 13056 12544
rect 12992 12484 12996 12540
rect 12996 12484 13052 12540
rect 13052 12484 13056 12540
rect 12992 12480 13056 12484
rect 13072 12540 13136 12544
rect 13072 12484 13076 12540
rect 13076 12484 13132 12540
rect 13132 12484 13136 12540
rect 13072 12480 13136 12484
rect 13152 12540 13216 12544
rect 13152 12484 13156 12540
rect 13156 12484 13212 12540
rect 13212 12484 13216 12540
rect 13152 12480 13216 12484
rect 3942 11996 4006 12000
rect 3942 11940 3946 11996
rect 3946 11940 4002 11996
rect 4002 11940 4006 11996
rect 3942 11936 4006 11940
rect 4022 11996 4086 12000
rect 4022 11940 4026 11996
rect 4026 11940 4082 11996
rect 4082 11940 4086 11996
rect 4022 11936 4086 11940
rect 4102 11996 4166 12000
rect 4102 11940 4106 11996
rect 4106 11940 4162 11996
rect 4162 11940 4166 11996
rect 4102 11936 4166 11940
rect 4182 11996 4246 12000
rect 4182 11940 4186 11996
rect 4186 11940 4242 11996
rect 4242 11940 4246 11996
rect 4182 11936 4246 11940
rect 9922 11996 9986 12000
rect 9922 11940 9926 11996
rect 9926 11940 9982 11996
rect 9982 11940 9986 11996
rect 9922 11936 9986 11940
rect 10002 11996 10066 12000
rect 10002 11940 10006 11996
rect 10006 11940 10062 11996
rect 10062 11940 10066 11996
rect 10002 11936 10066 11940
rect 10082 11996 10146 12000
rect 10082 11940 10086 11996
rect 10086 11940 10142 11996
rect 10142 11940 10146 11996
rect 10082 11936 10146 11940
rect 10162 11996 10226 12000
rect 10162 11940 10166 11996
rect 10166 11940 10222 11996
rect 10222 11940 10226 11996
rect 10162 11936 10226 11940
rect 15902 11996 15966 12000
rect 15902 11940 15906 11996
rect 15906 11940 15962 11996
rect 15962 11940 15966 11996
rect 15902 11936 15966 11940
rect 15982 11996 16046 12000
rect 15982 11940 15986 11996
rect 15986 11940 16042 11996
rect 16042 11940 16046 11996
rect 15982 11936 16046 11940
rect 16062 11996 16126 12000
rect 16062 11940 16066 11996
rect 16066 11940 16122 11996
rect 16122 11940 16126 11996
rect 16062 11936 16126 11940
rect 16142 11996 16206 12000
rect 16142 11940 16146 11996
rect 16146 11940 16202 11996
rect 16202 11940 16206 11996
rect 16142 11936 16206 11940
rect 6932 11452 6996 11456
rect 6932 11396 6936 11452
rect 6936 11396 6992 11452
rect 6992 11396 6996 11452
rect 6932 11392 6996 11396
rect 7012 11452 7076 11456
rect 7012 11396 7016 11452
rect 7016 11396 7072 11452
rect 7072 11396 7076 11452
rect 7012 11392 7076 11396
rect 7092 11452 7156 11456
rect 7092 11396 7096 11452
rect 7096 11396 7152 11452
rect 7152 11396 7156 11452
rect 7092 11392 7156 11396
rect 7172 11452 7236 11456
rect 7172 11396 7176 11452
rect 7176 11396 7232 11452
rect 7232 11396 7236 11452
rect 7172 11392 7236 11396
rect 12912 11452 12976 11456
rect 12912 11396 12916 11452
rect 12916 11396 12972 11452
rect 12972 11396 12976 11452
rect 12912 11392 12976 11396
rect 12992 11452 13056 11456
rect 12992 11396 12996 11452
rect 12996 11396 13052 11452
rect 13052 11396 13056 11452
rect 12992 11392 13056 11396
rect 13072 11452 13136 11456
rect 13072 11396 13076 11452
rect 13076 11396 13132 11452
rect 13132 11396 13136 11452
rect 13072 11392 13136 11396
rect 13152 11452 13216 11456
rect 13152 11396 13156 11452
rect 13156 11396 13212 11452
rect 13212 11396 13216 11452
rect 13152 11392 13216 11396
rect 3942 10908 4006 10912
rect 3942 10852 3946 10908
rect 3946 10852 4002 10908
rect 4002 10852 4006 10908
rect 3942 10848 4006 10852
rect 4022 10908 4086 10912
rect 4022 10852 4026 10908
rect 4026 10852 4082 10908
rect 4082 10852 4086 10908
rect 4022 10848 4086 10852
rect 4102 10908 4166 10912
rect 4102 10852 4106 10908
rect 4106 10852 4162 10908
rect 4162 10852 4166 10908
rect 4102 10848 4166 10852
rect 4182 10908 4246 10912
rect 4182 10852 4186 10908
rect 4186 10852 4242 10908
rect 4242 10852 4246 10908
rect 4182 10848 4246 10852
rect 9922 10908 9986 10912
rect 9922 10852 9926 10908
rect 9926 10852 9982 10908
rect 9982 10852 9986 10908
rect 9922 10848 9986 10852
rect 10002 10908 10066 10912
rect 10002 10852 10006 10908
rect 10006 10852 10062 10908
rect 10062 10852 10066 10908
rect 10002 10848 10066 10852
rect 10082 10908 10146 10912
rect 10082 10852 10086 10908
rect 10086 10852 10142 10908
rect 10142 10852 10146 10908
rect 10082 10848 10146 10852
rect 10162 10908 10226 10912
rect 10162 10852 10166 10908
rect 10166 10852 10222 10908
rect 10222 10852 10226 10908
rect 10162 10848 10226 10852
rect 15902 10908 15966 10912
rect 15902 10852 15906 10908
rect 15906 10852 15962 10908
rect 15962 10852 15966 10908
rect 15902 10848 15966 10852
rect 15982 10908 16046 10912
rect 15982 10852 15986 10908
rect 15986 10852 16042 10908
rect 16042 10852 16046 10908
rect 15982 10848 16046 10852
rect 16062 10908 16126 10912
rect 16062 10852 16066 10908
rect 16066 10852 16122 10908
rect 16122 10852 16126 10908
rect 16062 10848 16126 10852
rect 16142 10908 16206 10912
rect 16142 10852 16146 10908
rect 16146 10852 16202 10908
rect 16202 10852 16206 10908
rect 16142 10848 16206 10852
rect 6932 10364 6996 10368
rect 6932 10308 6936 10364
rect 6936 10308 6992 10364
rect 6992 10308 6996 10364
rect 6932 10304 6996 10308
rect 7012 10364 7076 10368
rect 7012 10308 7016 10364
rect 7016 10308 7072 10364
rect 7072 10308 7076 10364
rect 7012 10304 7076 10308
rect 7092 10364 7156 10368
rect 7092 10308 7096 10364
rect 7096 10308 7152 10364
rect 7152 10308 7156 10364
rect 7092 10304 7156 10308
rect 7172 10364 7236 10368
rect 7172 10308 7176 10364
rect 7176 10308 7232 10364
rect 7232 10308 7236 10364
rect 7172 10304 7236 10308
rect 12912 10364 12976 10368
rect 12912 10308 12916 10364
rect 12916 10308 12972 10364
rect 12972 10308 12976 10364
rect 12912 10304 12976 10308
rect 12992 10364 13056 10368
rect 12992 10308 12996 10364
rect 12996 10308 13052 10364
rect 13052 10308 13056 10364
rect 12992 10304 13056 10308
rect 13072 10364 13136 10368
rect 13072 10308 13076 10364
rect 13076 10308 13132 10364
rect 13132 10308 13136 10364
rect 13072 10304 13136 10308
rect 13152 10364 13216 10368
rect 13152 10308 13156 10364
rect 13156 10308 13212 10364
rect 13212 10308 13216 10364
rect 13152 10304 13216 10308
rect 3942 9820 4006 9824
rect 3942 9764 3946 9820
rect 3946 9764 4002 9820
rect 4002 9764 4006 9820
rect 3942 9760 4006 9764
rect 4022 9820 4086 9824
rect 4022 9764 4026 9820
rect 4026 9764 4082 9820
rect 4082 9764 4086 9820
rect 4022 9760 4086 9764
rect 4102 9820 4166 9824
rect 4102 9764 4106 9820
rect 4106 9764 4162 9820
rect 4162 9764 4166 9820
rect 4102 9760 4166 9764
rect 4182 9820 4246 9824
rect 4182 9764 4186 9820
rect 4186 9764 4242 9820
rect 4242 9764 4246 9820
rect 4182 9760 4246 9764
rect 9922 9820 9986 9824
rect 9922 9764 9926 9820
rect 9926 9764 9982 9820
rect 9982 9764 9986 9820
rect 9922 9760 9986 9764
rect 10002 9820 10066 9824
rect 10002 9764 10006 9820
rect 10006 9764 10062 9820
rect 10062 9764 10066 9820
rect 10002 9760 10066 9764
rect 10082 9820 10146 9824
rect 10082 9764 10086 9820
rect 10086 9764 10142 9820
rect 10142 9764 10146 9820
rect 10082 9760 10146 9764
rect 10162 9820 10226 9824
rect 10162 9764 10166 9820
rect 10166 9764 10222 9820
rect 10222 9764 10226 9820
rect 10162 9760 10226 9764
rect 15902 9820 15966 9824
rect 15902 9764 15906 9820
rect 15906 9764 15962 9820
rect 15962 9764 15966 9820
rect 15902 9760 15966 9764
rect 15982 9820 16046 9824
rect 15982 9764 15986 9820
rect 15986 9764 16042 9820
rect 16042 9764 16046 9820
rect 15982 9760 16046 9764
rect 16062 9820 16126 9824
rect 16062 9764 16066 9820
rect 16066 9764 16122 9820
rect 16122 9764 16126 9820
rect 16062 9760 16126 9764
rect 16142 9820 16206 9824
rect 16142 9764 16146 9820
rect 16146 9764 16202 9820
rect 16202 9764 16206 9820
rect 16142 9760 16206 9764
rect 6932 9276 6996 9280
rect 6932 9220 6936 9276
rect 6936 9220 6992 9276
rect 6992 9220 6996 9276
rect 6932 9216 6996 9220
rect 7012 9276 7076 9280
rect 7012 9220 7016 9276
rect 7016 9220 7072 9276
rect 7072 9220 7076 9276
rect 7012 9216 7076 9220
rect 7092 9276 7156 9280
rect 7092 9220 7096 9276
rect 7096 9220 7152 9276
rect 7152 9220 7156 9276
rect 7092 9216 7156 9220
rect 7172 9276 7236 9280
rect 7172 9220 7176 9276
rect 7176 9220 7232 9276
rect 7232 9220 7236 9276
rect 7172 9216 7236 9220
rect 12912 9276 12976 9280
rect 12912 9220 12916 9276
rect 12916 9220 12972 9276
rect 12972 9220 12976 9276
rect 12912 9216 12976 9220
rect 12992 9276 13056 9280
rect 12992 9220 12996 9276
rect 12996 9220 13052 9276
rect 13052 9220 13056 9276
rect 12992 9216 13056 9220
rect 13072 9276 13136 9280
rect 13072 9220 13076 9276
rect 13076 9220 13132 9276
rect 13132 9220 13136 9276
rect 13072 9216 13136 9220
rect 13152 9276 13216 9280
rect 13152 9220 13156 9276
rect 13156 9220 13212 9276
rect 13212 9220 13216 9276
rect 13152 9216 13216 9220
rect 3942 8732 4006 8736
rect 3942 8676 3946 8732
rect 3946 8676 4002 8732
rect 4002 8676 4006 8732
rect 3942 8672 4006 8676
rect 4022 8732 4086 8736
rect 4022 8676 4026 8732
rect 4026 8676 4082 8732
rect 4082 8676 4086 8732
rect 4022 8672 4086 8676
rect 4102 8732 4166 8736
rect 4102 8676 4106 8732
rect 4106 8676 4162 8732
rect 4162 8676 4166 8732
rect 4102 8672 4166 8676
rect 4182 8732 4246 8736
rect 4182 8676 4186 8732
rect 4186 8676 4242 8732
rect 4242 8676 4246 8732
rect 4182 8672 4246 8676
rect 9922 8732 9986 8736
rect 9922 8676 9926 8732
rect 9926 8676 9982 8732
rect 9982 8676 9986 8732
rect 9922 8672 9986 8676
rect 10002 8732 10066 8736
rect 10002 8676 10006 8732
rect 10006 8676 10062 8732
rect 10062 8676 10066 8732
rect 10002 8672 10066 8676
rect 10082 8732 10146 8736
rect 10082 8676 10086 8732
rect 10086 8676 10142 8732
rect 10142 8676 10146 8732
rect 10082 8672 10146 8676
rect 10162 8732 10226 8736
rect 10162 8676 10166 8732
rect 10166 8676 10222 8732
rect 10222 8676 10226 8732
rect 10162 8672 10226 8676
rect 15902 8732 15966 8736
rect 15902 8676 15906 8732
rect 15906 8676 15962 8732
rect 15962 8676 15966 8732
rect 15902 8672 15966 8676
rect 15982 8732 16046 8736
rect 15982 8676 15986 8732
rect 15986 8676 16042 8732
rect 16042 8676 16046 8732
rect 15982 8672 16046 8676
rect 16062 8732 16126 8736
rect 16062 8676 16066 8732
rect 16066 8676 16122 8732
rect 16122 8676 16126 8732
rect 16062 8672 16126 8676
rect 16142 8732 16206 8736
rect 16142 8676 16146 8732
rect 16146 8676 16202 8732
rect 16202 8676 16206 8732
rect 16142 8672 16206 8676
rect 6932 8188 6996 8192
rect 6932 8132 6936 8188
rect 6936 8132 6992 8188
rect 6992 8132 6996 8188
rect 6932 8128 6996 8132
rect 7012 8188 7076 8192
rect 7012 8132 7016 8188
rect 7016 8132 7072 8188
rect 7072 8132 7076 8188
rect 7012 8128 7076 8132
rect 7092 8188 7156 8192
rect 7092 8132 7096 8188
rect 7096 8132 7152 8188
rect 7152 8132 7156 8188
rect 7092 8128 7156 8132
rect 7172 8188 7236 8192
rect 7172 8132 7176 8188
rect 7176 8132 7232 8188
rect 7232 8132 7236 8188
rect 7172 8128 7236 8132
rect 12912 8188 12976 8192
rect 12912 8132 12916 8188
rect 12916 8132 12972 8188
rect 12972 8132 12976 8188
rect 12912 8128 12976 8132
rect 12992 8188 13056 8192
rect 12992 8132 12996 8188
rect 12996 8132 13052 8188
rect 13052 8132 13056 8188
rect 12992 8128 13056 8132
rect 13072 8188 13136 8192
rect 13072 8132 13076 8188
rect 13076 8132 13132 8188
rect 13132 8132 13136 8188
rect 13072 8128 13136 8132
rect 13152 8188 13216 8192
rect 13152 8132 13156 8188
rect 13156 8132 13212 8188
rect 13212 8132 13216 8188
rect 13152 8128 13216 8132
rect 3942 7644 4006 7648
rect 3942 7588 3946 7644
rect 3946 7588 4002 7644
rect 4002 7588 4006 7644
rect 3942 7584 4006 7588
rect 4022 7644 4086 7648
rect 4022 7588 4026 7644
rect 4026 7588 4082 7644
rect 4082 7588 4086 7644
rect 4022 7584 4086 7588
rect 4102 7644 4166 7648
rect 4102 7588 4106 7644
rect 4106 7588 4162 7644
rect 4162 7588 4166 7644
rect 4102 7584 4166 7588
rect 4182 7644 4246 7648
rect 4182 7588 4186 7644
rect 4186 7588 4242 7644
rect 4242 7588 4246 7644
rect 4182 7584 4246 7588
rect 9922 7644 9986 7648
rect 9922 7588 9926 7644
rect 9926 7588 9982 7644
rect 9982 7588 9986 7644
rect 9922 7584 9986 7588
rect 10002 7644 10066 7648
rect 10002 7588 10006 7644
rect 10006 7588 10062 7644
rect 10062 7588 10066 7644
rect 10002 7584 10066 7588
rect 10082 7644 10146 7648
rect 10082 7588 10086 7644
rect 10086 7588 10142 7644
rect 10142 7588 10146 7644
rect 10082 7584 10146 7588
rect 10162 7644 10226 7648
rect 10162 7588 10166 7644
rect 10166 7588 10222 7644
rect 10222 7588 10226 7644
rect 10162 7584 10226 7588
rect 15902 7644 15966 7648
rect 15902 7588 15906 7644
rect 15906 7588 15962 7644
rect 15962 7588 15966 7644
rect 15902 7584 15966 7588
rect 15982 7644 16046 7648
rect 15982 7588 15986 7644
rect 15986 7588 16042 7644
rect 16042 7588 16046 7644
rect 15982 7584 16046 7588
rect 16062 7644 16126 7648
rect 16062 7588 16066 7644
rect 16066 7588 16122 7644
rect 16122 7588 16126 7644
rect 16062 7584 16126 7588
rect 16142 7644 16206 7648
rect 16142 7588 16146 7644
rect 16146 7588 16202 7644
rect 16202 7588 16206 7644
rect 16142 7584 16206 7588
rect 6932 7100 6996 7104
rect 6932 7044 6936 7100
rect 6936 7044 6992 7100
rect 6992 7044 6996 7100
rect 6932 7040 6996 7044
rect 7012 7100 7076 7104
rect 7012 7044 7016 7100
rect 7016 7044 7072 7100
rect 7072 7044 7076 7100
rect 7012 7040 7076 7044
rect 7092 7100 7156 7104
rect 7092 7044 7096 7100
rect 7096 7044 7152 7100
rect 7152 7044 7156 7100
rect 7092 7040 7156 7044
rect 7172 7100 7236 7104
rect 7172 7044 7176 7100
rect 7176 7044 7232 7100
rect 7232 7044 7236 7100
rect 7172 7040 7236 7044
rect 12912 7100 12976 7104
rect 12912 7044 12916 7100
rect 12916 7044 12972 7100
rect 12972 7044 12976 7100
rect 12912 7040 12976 7044
rect 12992 7100 13056 7104
rect 12992 7044 12996 7100
rect 12996 7044 13052 7100
rect 13052 7044 13056 7100
rect 12992 7040 13056 7044
rect 13072 7100 13136 7104
rect 13072 7044 13076 7100
rect 13076 7044 13132 7100
rect 13132 7044 13136 7100
rect 13072 7040 13136 7044
rect 13152 7100 13216 7104
rect 13152 7044 13156 7100
rect 13156 7044 13212 7100
rect 13212 7044 13216 7100
rect 13152 7040 13216 7044
rect 3942 6556 4006 6560
rect 3942 6500 3946 6556
rect 3946 6500 4002 6556
rect 4002 6500 4006 6556
rect 3942 6496 4006 6500
rect 4022 6556 4086 6560
rect 4022 6500 4026 6556
rect 4026 6500 4082 6556
rect 4082 6500 4086 6556
rect 4022 6496 4086 6500
rect 4102 6556 4166 6560
rect 4102 6500 4106 6556
rect 4106 6500 4162 6556
rect 4162 6500 4166 6556
rect 4102 6496 4166 6500
rect 4182 6556 4246 6560
rect 4182 6500 4186 6556
rect 4186 6500 4242 6556
rect 4242 6500 4246 6556
rect 4182 6496 4246 6500
rect 9922 6556 9986 6560
rect 9922 6500 9926 6556
rect 9926 6500 9982 6556
rect 9982 6500 9986 6556
rect 9922 6496 9986 6500
rect 10002 6556 10066 6560
rect 10002 6500 10006 6556
rect 10006 6500 10062 6556
rect 10062 6500 10066 6556
rect 10002 6496 10066 6500
rect 10082 6556 10146 6560
rect 10082 6500 10086 6556
rect 10086 6500 10142 6556
rect 10142 6500 10146 6556
rect 10082 6496 10146 6500
rect 10162 6556 10226 6560
rect 10162 6500 10166 6556
rect 10166 6500 10222 6556
rect 10222 6500 10226 6556
rect 10162 6496 10226 6500
rect 15902 6556 15966 6560
rect 15902 6500 15906 6556
rect 15906 6500 15962 6556
rect 15962 6500 15966 6556
rect 15902 6496 15966 6500
rect 15982 6556 16046 6560
rect 15982 6500 15986 6556
rect 15986 6500 16042 6556
rect 16042 6500 16046 6556
rect 15982 6496 16046 6500
rect 16062 6556 16126 6560
rect 16062 6500 16066 6556
rect 16066 6500 16122 6556
rect 16122 6500 16126 6556
rect 16062 6496 16126 6500
rect 16142 6556 16206 6560
rect 16142 6500 16146 6556
rect 16146 6500 16202 6556
rect 16202 6500 16206 6556
rect 16142 6496 16206 6500
rect 6932 6012 6996 6016
rect 6932 5956 6936 6012
rect 6936 5956 6992 6012
rect 6992 5956 6996 6012
rect 6932 5952 6996 5956
rect 7012 6012 7076 6016
rect 7012 5956 7016 6012
rect 7016 5956 7072 6012
rect 7072 5956 7076 6012
rect 7012 5952 7076 5956
rect 7092 6012 7156 6016
rect 7092 5956 7096 6012
rect 7096 5956 7152 6012
rect 7152 5956 7156 6012
rect 7092 5952 7156 5956
rect 7172 6012 7236 6016
rect 7172 5956 7176 6012
rect 7176 5956 7232 6012
rect 7232 5956 7236 6012
rect 7172 5952 7236 5956
rect 12912 6012 12976 6016
rect 12912 5956 12916 6012
rect 12916 5956 12972 6012
rect 12972 5956 12976 6012
rect 12912 5952 12976 5956
rect 12992 6012 13056 6016
rect 12992 5956 12996 6012
rect 12996 5956 13052 6012
rect 13052 5956 13056 6012
rect 12992 5952 13056 5956
rect 13072 6012 13136 6016
rect 13072 5956 13076 6012
rect 13076 5956 13132 6012
rect 13132 5956 13136 6012
rect 13072 5952 13136 5956
rect 13152 6012 13216 6016
rect 13152 5956 13156 6012
rect 13156 5956 13212 6012
rect 13212 5956 13216 6012
rect 13152 5952 13216 5956
rect 3942 5468 4006 5472
rect 3942 5412 3946 5468
rect 3946 5412 4002 5468
rect 4002 5412 4006 5468
rect 3942 5408 4006 5412
rect 4022 5468 4086 5472
rect 4022 5412 4026 5468
rect 4026 5412 4082 5468
rect 4082 5412 4086 5468
rect 4022 5408 4086 5412
rect 4102 5468 4166 5472
rect 4102 5412 4106 5468
rect 4106 5412 4162 5468
rect 4162 5412 4166 5468
rect 4102 5408 4166 5412
rect 4182 5468 4246 5472
rect 4182 5412 4186 5468
rect 4186 5412 4242 5468
rect 4242 5412 4246 5468
rect 4182 5408 4246 5412
rect 9922 5468 9986 5472
rect 9922 5412 9926 5468
rect 9926 5412 9982 5468
rect 9982 5412 9986 5468
rect 9922 5408 9986 5412
rect 10002 5468 10066 5472
rect 10002 5412 10006 5468
rect 10006 5412 10062 5468
rect 10062 5412 10066 5468
rect 10002 5408 10066 5412
rect 10082 5468 10146 5472
rect 10082 5412 10086 5468
rect 10086 5412 10142 5468
rect 10142 5412 10146 5468
rect 10082 5408 10146 5412
rect 10162 5468 10226 5472
rect 10162 5412 10166 5468
rect 10166 5412 10222 5468
rect 10222 5412 10226 5468
rect 10162 5408 10226 5412
rect 15902 5468 15966 5472
rect 15902 5412 15906 5468
rect 15906 5412 15962 5468
rect 15962 5412 15966 5468
rect 15902 5408 15966 5412
rect 15982 5468 16046 5472
rect 15982 5412 15986 5468
rect 15986 5412 16042 5468
rect 16042 5412 16046 5468
rect 15982 5408 16046 5412
rect 16062 5468 16126 5472
rect 16062 5412 16066 5468
rect 16066 5412 16122 5468
rect 16122 5412 16126 5468
rect 16062 5408 16126 5412
rect 16142 5468 16206 5472
rect 16142 5412 16146 5468
rect 16146 5412 16202 5468
rect 16202 5412 16206 5468
rect 16142 5408 16206 5412
rect 6932 4924 6996 4928
rect 6932 4868 6936 4924
rect 6936 4868 6992 4924
rect 6992 4868 6996 4924
rect 6932 4864 6996 4868
rect 7012 4924 7076 4928
rect 7012 4868 7016 4924
rect 7016 4868 7072 4924
rect 7072 4868 7076 4924
rect 7012 4864 7076 4868
rect 7092 4924 7156 4928
rect 7092 4868 7096 4924
rect 7096 4868 7152 4924
rect 7152 4868 7156 4924
rect 7092 4864 7156 4868
rect 7172 4924 7236 4928
rect 7172 4868 7176 4924
rect 7176 4868 7232 4924
rect 7232 4868 7236 4924
rect 7172 4864 7236 4868
rect 12912 4924 12976 4928
rect 12912 4868 12916 4924
rect 12916 4868 12972 4924
rect 12972 4868 12976 4924
rect 12912 4864 12976 4868
rect 12992 4924 13056 4928
rect 12992 4868 12996 4924
rect 12996 4868 13052 4924
rect 13052 4868 13056 4924
rect 12992 4864 13056 4868
rect 13072 4924 13136 4928
rect 13072 4868 13076 4924
rect 13076 4868 13132 4924
rect 13132 4868 13136 4924
rect 13072 4864 13136 4868
rect 13152 4924 13216 4928
rect 13152 4868 13156 4924
rect 13156 4868 13212 4924
rect 13212 4868 13216 4924
rect 13152 4864 13216 4868
rect 3942 4380 4006 4384
rect 3942 4324 3946 4380
rect 3946 4324 4002 4380
rect 4002 4324 4006 4380
rect 3942 4320 4006 4324
rect 4022 4380 4086 4384
rect 4022 4324 4026 4380
rect 4026 4324 4082 4380
rect 4082 4324 4086 4380
rect 4022 4320 4086 4324
rect 4102 4380 4166 4384
rect 4102 4324 4106 4380
rect 4106 4324 4162 4380
rect 4162 4324 4166 4380
rect 4102 4320 4166 4324
rect 4182 4380 4246 4384
rect 4182 4324 4186 4380
rect 4186 4324 4242 4380
rect 4242 4324 4246 4380
rect 4182 4320 4246 4324
rect 9922 4380 9986 4384
rect 9922 4324 9926 4380
rect 9926 4324 9982 4380
rect 9982 4324 9986 4380
rect 9922 4320 9986 4324
rect 10002 4380 10066 4384
rect 10002 4324 10006 4380
rect 10006 4324 10062 4380
rect 10062 4324 10066 4380
rect 10002 4320 10066 4324
rect 10082 4380 10146 4384
rect 10082 4324 10086 4380
rect 10086 4324 10142 4380
rect 10142 4324 10146 4380
rect 10082 4320 10146 4324
rect 10162 4380 10226 4384
rect 10162 4324 10166 4380
rect 10166 4324 10222 4380
rect 10222 4324 10226 4380
rect 10162 4320 10226 4324
rect 15902 4380 15966 4384
rect 15902 4324 15906 4380
rect 15906 4324 15962 4380
rect 15962 4324 15966 4380
rect 15902 4320 15966 4324
rect 15982 4380 16046 4384
rect 15982 4324 15986 4380
rect 15986 4324 16042 4380
rect 16042 4324 16046 4380
rect 15982 4320 16046 4324
rect 16062 4380 16126 4384
rect 16062 4324 16066 4380
rect 16066 4324 16122 4380
rect 16122 4324 16126 4380
rect 16062 4320 16126 4324
rect 16142 4380 16206 4384
rect 16142 4324 16146 4380
rect 16146 4324 16202 4380
rect 16202 4324 16206 4380
rect 16142 4320 16206 4324
rect 6932 3836 6996 3840
rect 6932 3780 6936 3836
rect 6936 3780 6992 3836
rect 6992 3780 6996 3836
rect 6932 3776 6996 3780
rect 7012 3836 7076 3840
rect 7012 3780 7016 3836
rect 7016 3780 7072 3836
rect 7072 3780 7076 3836
rect 7012 3776 7076 3780
rect 7092 3836 7156 3840
rect 7092 3780 7096 3836
rect 7096 3780 7152 3836
rect 7152 3780 7156 3836
rect 7092 3776 7156 3780
rect 7172 3836 7236 3840
rect 7172 3780 7176 3836
rect 7176 3780 7232 3836
rect 7232 3780 7236 3836
rect 7172 3776 7236 3780
rect 12912 3836 12976 3840
rect 12912 3780 12916 3836
rect 12916 3780 12972 3836
rect 12972 3780 12976 3836
rect 12912 3776 12976 3780
rect 12992 3836 13056 3840
rect 12992 3780 12996 3836
rect 12996 3780 13052 3836
rect 13052 3780 13056 3836
rect 12992 3776 13056 3780
rect 13072 3836 13136 3840
rect 13072 3780 13076 3836
rect 13076 3780 13132 3836
rect 13132 3780 13136 3836
rect 13072 3776 13136 3780
rect 13152 3836 13216 3840
rect 13152 3780 13156 3836
rect 13156 3780 13212 3836
rect 13212 3780 13216 3836
rect 13152 3776 13216 3780
rect 3942 3292 4006 3296
rect 3942 3236 3946 3292
rect 3946 3236 4002 3292
rect 4002 3236 4006 3292
rect 3942 3232 4006 3236
rect 4022 3292 4086 3296
rect 4022 3236 4026 3292
rect 4026 3236 4082 3292
rect 4082 3236 4086 3292
rect 4022 3232 4086 3236
rect 4102 3292 4166 3296
rect 4102 3236 4106 3292
rect 4106 3236 4162 3292
rect 4162 3236 4166 3292
rect 4102 3232 4166 3236
rect 4182 3292 4246 3296
rect 4182 3236 4186 3292
rect 4186 3236 4242 3292
rect 4242 3236 4246 3292
rect 4182 3232 4246 3236
rect 9922 3292 9986 3296
rect 9922 3236 9926 3292
rect 9926 3236 9982 3292
rect 9982 3236 9986 3292
rect 9922 3232 9986 3236
rect 10002 3292 10066 3296
rect 10002 3236 10006 3292
rect 10006 3236 10062 3292
rect 10062 3236 10066 3292
rect 10002 3232 10066 3236
rect 10082 3292 10146 3296
rect 10082 3236 10086 3292
rect 10086 3236 10142 3292
rect 10142 3236 10146 3292
rect 10082 3232 10146 3236
rect 10162 3292 10226 3296
rect 10162 3236 10166 3292
rect 10166 3236 10222 3292
rect 10222 3236 10226 3292
rect 10162 3232 10226 3236
rect 15902 3292 15966 3296
rect 15902 3236 15906 3292
rect 15906 3236 15962 3292
rect 15962 3236 15966 3292
rect 15902 3232 15966 3236
rect 15982 3292 16046 3296
rect 15982 3236 15986 3292
rect 15986 3236 16042 3292
rect 16042 3236 16046 3292
rect 15982 3232 16046 3236
rect 16062 3292 16126 3296
rect 16062 3236 16066 3292
rect 16066 3236 16122 3292
rect 16122 3236 16126 3292
rect 16062 3232 16126 3236
rect 16142 3292 16206 3296
rect 16142 3236 16146 3292
rect 16146 3236 16202 3292
rect 16202 3236 16206 3292
rect 16142 3232 16206 3236
rect 6932 2748 6996 2752
rect 6932 2692 6936 2748
rect 6936 2692 6992 2748
rect 6992 2692 6996 2748
rect 6932 2688 6996 2692
rect 7012 2748 7076 2752
rect 7012 2692 7016 2748
rect 7016 2692 7072 2748
rect 7072 2692 7076 2748
rect 7012 2688 7076 2692
rect 7092 2748 7156 2752
rect 7092 2692 7096 2748
rect 7096 2692 7152 2748
rect 7152 2692 7156 2748
rect 7092 2688 7156 2692
rect 7172 2748 7236 2752
rect 7172 2692 7176 2748
rect 7176 2692 7232 2748
rect 7232 2692 7236 2748
rect 7172 2688 7236 2692
rect 12912 2748 12976 2752
rect 12912 2692 12916 2748
rect 12916 2692 12972 2748
rect 12972 2692 12976 2748
rect 12912 2688 12976 2692
rect 12992 2748 13056 2752
rect 12992 2692 12996 2748
rect 12996 2692 13052 2748
rect 13052 2692 13056 2748
rect 12992 2688 13056 2692
rect 13072 2748 13136 2752
rect 13072 2692 13076 2748
rect 13076 2692 13132 2748
rect 13132 2692 13136 2748
rect 13072 2688 13136 2692
rect 13152 2748 13216 2752
rect 13152 2692 13156 2748
rect 13156 2692 13212 2748
rect 13212 2692 13216 2748
rect 13152 2688 13216 2692
rect 3942 2204 4006 2208
rect 3942 2148 3946 2204
rect 3946 2148 4002 2204
rect 4002 2148 4006 2204
rect 3942 2144 4006 2148
rect 4022 2204 4086 2208
rect 4022 2148 4026 2204
rect 4026 2148 4082 2204
rect 4082 2148 4086 2204
rect 4022 2144 4086 2148
rect 4102 2204 4166 2208
rect 4102 2148 4106 2204
rect 4106 2148 4162 2204
rect 4162 2148 4166 2204
rect 4102 2144 4166 2148
rect 4182 2204 4246 2208
rect 4182 2148 4186 2204
rect 4186 2148 4242 2204
rect 4242 2148 4246 2204
rect 4182 2144 4246 2148
rect 9922 2204 9986 2208
rect 9922 2148 9926 2204
rect 9926 2148 9982 2204
rect 9982 2148 9986 2204
rect 9922 2144 9986 2148
rect 10002 2204 10066 2208
rect 10002 2148 10006 2204
rect 10006 2148 10062 2204
rect 10062 2148 10066 2204
rect 10002 2144 10066 2148
rect 10082 2204 10146 2208
rect 10082 2148 10086 2204
rect 10086 2148 10142 2204
rect 10142 2148 10146 2204
rect 10082 2144 10146 2148
rect 10162 2204 10226 2208
rect 10162 2148 10166 2204
rect 10166 2148 10222 2204
rect 10222 2148 10226 2204
rect 10162 2144 10226 2148
rect 15902 2204 15966 2208
rect 15902 2148 15906 2204
rect 15906 2148 15962 2204
rect 15962 2148 15966 2204
rect 15902 2144 15966 2148
rect 15982 2204 16046 2208
rect 15982 2148 15986 2204
rect 15986 2148 16042 2204
rect 16042 2148 16046 2204
rect 15982 2144 16046 2148
rect 16062 2204 16126 2208
rect 16062 2148 16066 2204
rect 16066 2148 16122 2204
rect 16122 2148 16126 2204
rect 16062 2144 16126 2148
rect 16142 2204 16206 2208
rect 16142 2148 16146 2204
rect 16146 2148 16202 2204
rect 16202 2148 16206 2204
rect 16142 2144 16206 2148
<< metal4 >>
rect 3934 19616 4254 20176
rect 3934 19552 3942 19616
rect 4006 19552 4022 19616
rect 4086 19552 4102 19616
rect 4166 19552 4182 19616
rect 4246 19552 4254 19616
rect 3934 18528 4254 19552
rect 3934 18464 3942 18528
rect 4006 18464 4022 18528
rect 4086 18464 4102 18528
rect 4166 18464 4182 18528
rect 4246 18464 4254 18528
rect 3934 17440 4254 18464
rect 3934 17376 3942 17440
rect 4006 17376 4022 17440
rect 4086 17376 4102 17440
rect 4166 17376 4182 17440
rect 4246 17376 4254 17440
rect 3934 17206 4254 17376
rect 3934 16970 3976 17206
rect 4212 16970 4254 17206
rect 3934 16352 4254 16970
rect 3934 16288 3942 16352
rect 4006 16288 4022 16352
rect 4086 16288 4102 16352
rect 4166 16288 4182 16352
rect 4246 16288 4254 16352
rect 3934 15264 4254 16288
rect 3934 15200 3942 15264
rect 4006 15200 4022 15264
rect 4086 15200 4102 15264
rect 4166 15200 4182 15264
rect 4246 15200 4254 15264
rect 3934 14176 4254 15200
rect 3934 14112 3942 14176
rect 4006 14112 4022 14176
rect 4086 14112 4102 14176
rect 4166 14112 4182 14176
rect 4246 14112 4254 14176
rect 3934 13088 4254 14112
rect 3934 13024 3942 13088
rect 4006 13024 4022 13088
rect 4086 13024 4102 13088
rect 4166 13024 4182 13088
rect 4246 13024 4254 13088
rect 3934 12000 4254 13024
rect 3934 11936 3942 12000
rect 4006 11936 4022 12000
rect 4086 11936 4102 12000
rect 4166 11936 4182 12000
rect 4246 11936 4254 12000
rect 3934 11222 4254 11936
rect 3934 10986 3976 11222
rect 4212 10986 4254 11222
rect 3934 10912 4254 10986
rect 3934 10848 3942 10912
rect 4006 10848 4022 10912
rect 4086 10848 4102 10912
rect 4166 10848 4182 10912
rect 4246 10848 4254 10912
rect 3934 9824 4254 10848
rect 3934 9760 3942 9824
rect 4006 9760 4022 9824
rect 4086 9760 4102 9824
rect 4166 9760 4182 9824
rect 4246 9760 4254 9824
rect 3934 8736 4254 9760
rect 3934 8672 3942 8736
rect 4006 8672 4022 8736
rect 4086 8672 4102 8736
rect 4166 8672 4182 8736
rect 4246 8672 4254 8736
rect 3934 7648 4254 8672
rect 3934 7584 3942 7648
rect 4006 7584 4022 7648
rect 4086 7584 4102 7648
rect 4166 7584 4182 7648
rect 4246 7584 4254 7648
rect 3934 6560 4254 7584
rect 3934 6496 3942 6560
rect 4006 6496 4022 6560
rect 4086 6496 4102 6560
rect 4166 6496 4182 6560
rect 4246 6496 4254 6560
rect 3934 5472 4254 6496
rect 3934 5408 3942 5472
rect 4006 5408 4022 5472
rect 4086 5408 4102 5472
rect 4166 5408 4182 5472
rect 4246 5408 4254 5472
rect 3934 5238 4254 5408
rect 3934 5002 3976 5238
rect 4212 5002 4254 5238
rect 3934 4384 4254 5002
rect 3934 4320 3942 4384
rect 4006 4320 4022 4384
rect 4086 4320 4102 4384
rect 4166 4320 4182 4384
rect 4246 4320 4254 4384
rect 3934 3296 4254 4320
rect 3934 3232 3942 3296
rect 4006 3232 4022 3296
rect 4086 3232 4102 3296
rect 4166 3232 4182 3296
rect 4246 3232 4254 3296
rect 3934 2208 4254 3232
rect 3934 2144 3942 2208
rect 4006 2144 4022 2208
rect 4086 2144 4102 2208
rect 4166 2144 4182 2208
rect 4246 2144 4254 2208
rect 3934 2128 4254 2144
rect 6924 20160 7244 20176
rect 6924 20096 6932 20160
rect 6996 20096 7012 20160
rect 7076 20096 7092 20160
rect 7156 20096 7172 20160
rect 7236 20096 7244 20160
rect 6924 19072 7244 20096
rect 6924 19008 6932 19072
rect 6996 19008 7012 19072
rect 7076 19008 7092 19072
rect 7156 19008 7172 19072
rect 7236 19008 7244 19072
rect 6924 17984 7244 19008
rect 6924 17920 6932 17984
rect 6996 17920 7012 17984
rect 7076 17920 7092 17984
rect 7156 17920 7172 17984
rect 7236 17920 7244 17984
rect 6924 16896 7244 17920
rect 6924 16832 6932 16896
rect 6996 16832 7012 16896
rect 7076 16832 7092 16896
rect 7156 16832 7172 16896
rect 7236 16832 7244 16896
rect 6924 15808 7244 16832
rect 6924 15744 6932 15808
rect 6996 15744 7012 15808
rect 7076 15744 7092 15808
rect 7156 15744 7172 15808
rect 7236 15744 7244 15808
rect 6924 14720 7244 15744
rect 6924 14656 6932 14720
rect 6996 14656 7012 14720
rect 7076 14656 7092 14720
rect 7156 14656 7172 14720
rect 7236 14656 7244 14720
rect 6924 14214 7244 14656
rect 6924 13978 6966 14214
rect 7202 13978 7244 14214
rect 6924 13632 7244 13978
rect 6924 13568 6932 13632
rect 6996 13568 7012 13632
rect 7076 13568 7092 13632
rect 7156 13568 7172 13632
rect 7236 13568 7244 13632
rect 6924 12544 7244 13568
rect 6924 12480 6932 12544
rect 6996 12480 7012 12544
rect 7076 12480 7092 12544
rect 7156 12480 7172 12544
rect 7236 12480 7244 12544
rect 6924 11456 7244 12480
rect 6924 11392 6932 11456
rect 6996 11392 7012 11456
rect 7076 11392 7092 11456
rect 7156 11392 7172 11456
rect 7236 11392 7244 11456
rect 6924 10368 7244 11392
rect 6924 10304 6932 10368
rect 6996 10304 7012 10368
rect 7076 10304 7092 10368
rect 7156 10304 7172 10368
rect 7236 10304 7244 10368
rect 6924 9280 7244 10304
rect 6924 9216 6932 9280
rect 6996 9216 7012 9280
rect 7076 9216 7092 9280
rect 7156 9216 7172 9280
rect 7236 9216 7244 9280
rect 6924 8230 7244 9216
rect 6924 8192 6966 8230
rect 7202 8192 7244 8230
rect 6924 8128 6932 8192
rect 7236 8128 7244 8192
rect 6924 7994 6966 8128
rect 7202 7994 7244 8128
rect 6924 7104 7244 7994
rect 6924 7040 6932 7104
rect 6996 7040 7012 7104
rect 7076 7040 7092 7104
rect 7156 7040 7172 7104
rect 7236 7040 7244 7104
rect 6924 6016 7244 7040
rect 6924 5952 6932 6016
rect 6996 5952 7012 6016
rect 7076 5952 7092 6016
rect 7156 5952 7172 6016
rect 7236 5952 7244 6016
rect 6924 4928 7244 5952
rect 6924 4864 6932 4928
rect 6996 4864 7012 4928
rect 7076 4864 7092 4928
rect 7156 4864 7172 4928
rect 7236 4864 7244 4928
rect 6924 3840 7244 4864
rect 6924 3776 6932 3840
rect 6996 3776 7012 3840
rect 7076 3776 7092 3840
rect 7156 3776 7172 3840
rect 7236 3776 7244 3840
rect 6924 2752 7244 3776
rect 6924 2688 6932 2752
rect 6996 2688 7012 2752
rect 7076 2688 7092 2752
rect 7156 2688 7172 2752
rect 7236 2688 7244 2752
rect 6924 2128 7244 2688
rect 9914 19616 10234 20176
rect 9914 19552 9922 19616
rect 9986 19552 10002 19616
rect 10066 19552 10082 19616
rect 10146 19552 10162 19616
rect 10226 19552 10234 19616
rect 9914 18528 10234 19552
rect 9914 18464 9922 18528
rect 9986 18464 10002 18528
rect 10066 18464 10082 18528
rect 10146 18464 10162 18528
rect 10226 18464 10234 18528
rect 9914 17440 10234 18464
rect 9914 17376 9922 17440
rect 9986 17376 10002 17440
rect 10066 17376 10082 17440
rect 10146 17376 10162 17440
rect 10226 17376 10234 17440
rect 9914 17206 10234 17376
rect 9914 16970 9956 17206
rect 10192 16970 10234 17206
rect 9914 16352 10234 16970
rect 9914 16288 9922 16352
rect 9986 16288 10002 16352
rect 10066 16288 10082 16352
rect 10146 16288 10162 16352
rect 10226 16288 10234 16352
rect 9914 15264 10234 16288
rect 9914 15200 9922 15264
rect 9986 15200 10002 15264
rect 10066 15200 10082 15264
rect 10146 15200 10162 15264
rect 10226 15200 10234 15264
rect 9914 14176 10234 15200
rect 9914 14112 9922 14176
rect 9986 14112 10002 14176
rect 10066 14112 10082 14176
rect 10146 14112 10162 14176
rect 10226 14112 10234 14176
rect 9914 13088 10234 14112
rect 9914 13024 9922 13088
rect 9986 13024 10002 13088
rect 10066 13024 10082 13088
rect 10146 13024 10162 13088
rect 10226 13024 10234 13088
rect 9914 12000 10234 13024
rect 9914 11936 9922 12000
rect 9986 11936 10002 12000
rect 10066 11936 10082 12000
rect 10146 11936 10162 12000
rect 10226 11936 10234 12000
rect 9914 11222 10234 11936
rect 9914 10986 9956 11222
rect 10192 10986 10234 11222
rect 9914 10912 10234 10986
rect 9914 10848 9922 10912
rect 9986 10848 10002 10912
rect 10066 10848 10082 10912
rect 10146 10848 10162 10912
rect 10226 10848 10234 10912
rect 9914 9824 10234 10848
rect 9914 9760 9922 9824
rect 9986 9760 10002 9824
rect 10066 9760 10082 9824
rect 10146 9760 10162 9824
rect 10226 9760 10234 9824
rect 9914 8736 10234 9760
rect 9914 8672 9922 8736
rect 9986 8672 10002 8736
rect 10066 8672 10082 8736
rect 10146 8672 10162 8736
rect 10226 8672 10234 8736
rect 9914 7648 10234 8672
rect 9914 7584 9922 7648
rect 9986 7584 10002 7648
rect 10066 7584 10082 7648
rect 10146 7584 10162 7648
rect 10226 7584 10234 7648
rect 9914 6560 10234 7584
rect 9914 6496 9922 6560
rect 9986 6496 10002 6560
rect 10066 6496 10082 6560
rect 10146 6496 10162 6560
rect 10226 6496 10234 6560
rect 9914 5472 10234 6496
rect 9914 5408 9922 5472
rect 9986 5408 10002 5472
rect 10066 5408 10082 5472
rect 10146 5408 10162 5472
rect 10226 5408 10234 5472
rect 9914 5238 10234 5408
rect 9914 5002 9956 5238
rect 10192 5002 10234 5238
rect 9914 4384 10234 5002
rect 9914 4320 9922 4384
rect 9986 4320 10002 4384
rect 10066 4320 10082 4384
rect 10146 4320 10162 4384
rect 10226 4320 10234 4384
rect 9914 3296 10234 4320
rect 9914 3232 9922 3296
rect 9986 3232 10002 3296
rect 10066 3232 10082 3296
rect 10146 3232 10162 3296
rect 10226 3232 10234 3296
rect 9914 2208 10234 3232
rect 9914 2144 9922 2208
rect 9986 2144 10002 2208
rect 10066 2144 10082 2208
rect 10146 2144 10162 2208
rect 10226 2144 10234 2208
rect 9914 2128 10234 2144
rect 12904 20160 13224 20176
rect 12904 20096 12912 20160
rect 12976 20096 12992 20160
rect 13056 20096 13072 20160
rect 13136 20096 13152 20160
rect 13216 20096 13224 20160
rect 12904 19072 13224 20096
rect 12904 19008 12912 19072
rect 12976 19008 12992 19072
rect 13056 19008 13072 19072
rect 13136 19008 13152 19072
rect 13216 19008 13224 19072
rect 12904 17984 13224 19008
rect 12904 17920 12912 17984
rect 12976 17920 12992 17984
rect 13056 17920 13072 17984
rect 13136 17920 13152 17984
rect 13216 17920 13224 17984
rect 12904 16896 13224 17920
rect 12904 16832 12912 16896
rect 12976 16832 12992 16896
rect 13056 16832 13072 16896
rect 13136 16832 13152 16896
rect 13216 16832 13224 16896
rect 12904 15808 13224 16832
rect 12904 15744 12912 15808
rect 12976 15744 12992 15808
rect 13056 15744 13072 15808
rect 13136 15744 13152 15808
rect 13216 15744 13224 15808
rect 12904 14720 13224 15744
rect 12904 14656 12912 14720
rect 12976 14656 12992 14720
rect 13056 14656 13072 14720
rect 13136 14656 13152 14720
rect 13216 14656 13224 14720
rect 12904 14214 13224 14656
rect 12904 13978 12946 14214
rect 13182 13978 13224 14214
rect 12904 13632 13224 13978
rect 12904 13568 12912 13632
rect 12976 13568 12992 13632
rect 13056 13568 13072 13632
rect 13136 13568 13152 13632
rect 13216 13568 13224 13632
rect 12904 12544 13224 13568
rect 12904 12480 12912 12544
rect 12976 12480 12992 12544
rect 13056 12480 13072 12544
rect 13136 12480 13152 12544
rect 13216 12480 13224 12544
rect 12904 11456 13224 12480
rect 12904 11392 12912 11456
rect 12976 11392 12992 11456
rect 13056 11392 13072 11456
rect 13136 11392 13152 11456
rect 13216 11392 13224 11456
rect 12904 10368 13224 11392
rect 12904 10304 12912 10368
rect 12976 10304 12992 10368
rect 13056 10304 13072 10368
rect 13136 10304 13152 10368
rect 13216 10304 13224 10368
rect 12904 9280 13224 10304
rect 12904 9216 12912 9280
rect 12976 9216 12992 9280
rect 13056 9216 13072 9280
rect 13136 9216 13152 9280
rect 13216 9216 13224 9280
rect 12904 8230 13224 9216
rect 12904 8192 12946 8230
rect 13182 8192 13224 8230
rect 12904 8128 12912 8192
rect 13216 8128 13224 8192
rect 12904 7994 12946 8128
rect 13182 7994 13224 8128
rect 12904 7104 13224 7994
rect 12904 7040 12912 7104
rect 12976 7040 12992 7104
rect 13056 7040 13072 7104
rect 13136 7040 13152 7104
rect 13216 7040 13224 7104
rect 12904 6016 13224 7040
rect 12904 5952 12912 6016
rect 12976 5952 12992 6016
rect 13056 5952 13072 6016
rect 13136 5952 13152 6016
rect 13216 5952 13224 6016
rect 12904 4928 13224 5952
rect 12904 4864 12912 4928
rect 12976 4864 12992 4928
rect 13056 4864 13072 4928
rect 13136 4864 13152 4928
rect 13216 4864 13224 4928
rect 12904 3840 13224 4864
rect 12904 3776 12912 3840
rect 12976 3776 12992 3840
rect 13056 3776 13072 3840
rect 13136 3776 13152 3840
rect 13216 3776 13224 3840
rect 12904 2752 13224 3776
rect 12904 2688 12912 2752
rect 12976 2688 12992 2752
rect 13056 2688 13072 2752
rect 13136 2688 13152 2752
rect 13216 2688 13224 2752
rect 12904 2128 13224 2688
rect 15894 19616 16214 20176
rect 15894 19552 15902 19616
rect 15966 19552 15982 19616
rect 16046 19552 16062 19616
rect 16126 19552 16142 19616
rect 16206 19552 16214 19616
rect 15894 18528 16214 19552
rect 15894 18464 15902 18528
rect 15966 18464 15982 18528
rect 16046 18464 16062 18528
rect 16126 18464 16142 18528
rect 16206 18464 16214 18528
rect 15894 17440 16214 18464
rect 15894 17376 15902 17440
rect 15966 17376 15982 17440
rect 16046 17376 16062 17440
rect 16126 17376 16142 17440
rect 16206 17376 16214 17440
rect 15894 17206 16214 17376
rect 15894 16970 15936 17206
rect 16172 16970 16214 17206
rect 15894 16352 16214 16970
rect 15894 16288 15902 16352
rect 15966 16288 15982 16352
rect 16046 16288 16062 16352
rect 16126 16288 16142 16352
rect 16206 16288 16214 16352
rect 15894 15264 16214 16288
rect 15894 15200 15902 15264
rect 15966 15200 15982 15264
rect 16046 15200 16062 15264
rect 16126 15200 16142 15264
rect 16206 15200 16214 15264
rect 15894 14176 16214 15200
rect 15894 14112 15902 14176
rect 15966 14112 15982 14176
rect 16046 14112 16062 14176
rect 16126 14112 16142 14176
rect 16206 14112 16214 14176
rect 15894 13088 16214 14112
rect 15894 13024 15902 13088
rect 15966 13024 15982 13088
rect 16046 13024 16062 13088
rect 16126 13024 16142 13088
rect 16206 13024 16214 13088
rect 15894 12000 16214 13024
rect 15894 11936 15902 12000
rect 15966 11936 15982 12000
rect 16046 11936 16062 12000
rect 16126 11936 16142 12000
rect 16206 11936 16214 12000
rect 15894 11222 16214 11936
rect 15894 10986 15936 11222
rect 16172 10986 16214 11222
rect 15894 10912 16214 10986
rect 15894 10848 15902 10912
rect 15966 10848 15982 10912
rect 16046 10848 16062 10912
rect 16126 10848 16142 10912
rect 16206 10848 16214 10912
rect 15894 9824 16214 10848
rect 15894 9760 15902 9824
rect 15966 9760 15982 9824
rect 16046 9760 16062 9824
rect 16126 9760 16142 9824
rect 16206 9760 16214 9824
rect 15894 8736 16214 9760
rect 15894 8672 15902 8736
rect 15966 8672 15982 8736
rect 16046 8672 16062 8736
rect 16126 8672 16142 8736
rect 16206 8672 16214 8736
rect 15894 7648 16214 8672
rect 15894 7584 15902 7648
rect 15966 7584 15982 7648
rect 16046 7584 16062 7648
rect 16126 7584 16142 7648
rect 16206 7584 16214 7648
rect 15894 6560 16214 7584
rect 15894 6496 15902 6560
rect 15966 6496 15982 6560
rect 16046 6496 16062 6560
rect 16126 6496 16142 6560
rect 16206 6496 16214 6560
rect 15894 5472 16214 6496
rect 15894 5408 15902 5472
rect 15966 5408 15982 5472
rect 16046 5408 16062 5472
rect 16126 5408 16142 5472
rect 16206 5408 16214 5472
rect 15894 5238 16214 5408
rect 15894 5002 15936 5238
rect 16172 5002 16214 5238
rect 15894 4384 16214 5002
rect 15894 4320 15902 4384
rect 15966 4320 15982 4384
rect 16046 4320 16062 4384
rect 16126 4320 16142 4384
rect 16206 4320 16214 4384
rect 15894 3296 16214 4320
rect 15894 3232 15902 3296
rect 15966 3232 15982 3296
rect 16046 3232 16062 3296
rect 16126 3232 16142 3296
rect 16206 3232 16214 3296
rect 15894 2208 16214 3232
rect 15894 2144 15902 2208
rect 15966 2144 15982 2208
rect 16046 2144 16062 2208
rect 16126 2144 16142 2208
rect 16206 2144 16214 2208
rect 15894 2128 16214 2144
<< via4 >>
rect 3976 16970 4212 17206
rect 3976 10986 4212 11222
rect 3976 5002 4212 5238
rect 6966 13978 7202 14214
rect 6966 8192 7202 8230
rect 6966 8128 6996 8192
rect 6996 8128 7012 8192
rect 7012 8128 7076 8192
rect 7076 8128 7092 8192
rect 7092 8128 7156 8192
rect 7156 8128 7172 8192
rect 7172 8128 7202 8192
rect 6966 7994 7202 8128
rect 9956 16970 10192 17206
rect 9956 10986 10192 11222
rect 9956 5002 10192 5238
rect 12946 13978 13182 14214
rect 12946 8192 13182 8230
rect 12946 8128 12976 8192
rect 12976 8128 12992 8192
rect 12992 8128 13056 8192
rect 13056 8128 13072 8192
rect 13072 8128 13136 8192
rect 13136 8128 13152 8192
rect 13152 8128 13182 8192
rect 12946 7994 13182 8128
rect 15936 16970 16172 17206
rect 15936 10986 16172 11222
rect 15936 5002 16172 5238
<< metal5 >>
rect 1104 17206 19044 17248
rect 1104 16970 3976 17206
rect 4212 16970 9956 17206
rect 10192 16970 15936 17206
rect 16172 16970 19044 17206
rect 1104 16928 19044 16970
rect 1104 14214 19044 14256
rect 1104 13978 6966 14214
rect 7202 13978 12946 14214
rect 13182 13978 19044 14214
rect 1104 13936 19044 13978
rect 1104 11222 19044 11264
rect 1104 10986 3976 11222
rect 4212 10986 9956 11222
rect 10192 10986 15936 11222
rect 16172 10986 19044 11222
rect 1104 10944 19044 10986
rect 1104 8230 19044 8272
rect 1104 7994 6966 8230
rect 7202 7994 12946 8230
rect 13182 7994 19044 8230
rect 1104 7952 19044 7994
rect 1104 5238 19044 5280
rect 1104 5002 3976 5238
rect 4212 5002 9956 5238
rect 10192 5002 15936 5238
rect 16172 5002 19044 5238
rect 1104 4960 19044 5002
use sky130_fd_sc_hd__decap_8  FILLER_0_12
timestamp 1619617919
transform 1 0 2208 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6
timestamp 1619617919
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output45
timestamp 1619617919
transform -1 0 2208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1619617919
transform -1 0 1656 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1619617919
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1619617919
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1619617919
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_18
timestamp 1619617919
transform 1 0 2760 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20
timestamp 1619617919
transform 1 0 2944 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1619617919
transform -1 0 3496 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_6
timestamp 1619617919
transform 1 0 1656 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrbp_2  idiv2
timestamp 1619617919
transform 1 0 3036 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1619617919
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1619617919
transform -1 0 4876 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26
timestamp 1619617919
transform 1 0 3496 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30
timestamp 1619617919
transform 1 0 3864 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1619617919
transform 1 0 4876 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_45
timestamp 1619617919
transform 1 0 5244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_56
timestamp 1619617919
transform 1 0 6256 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56
timestamp 1619617919
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1619617919
transform -1 0 6256 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1619617919
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1619617919
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  irb
timestamp 1619617919
transform 1 0 5796 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_1_70
timestamp 1619617919
transform 1 0 7544 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb1
timestamp 1619617919
transform 1 0 7820 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _369_
timestamp 1619617919
transform -1 0 8464 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_1_58
timestamp 1619617919
transform 1 0 6440 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_59
timestamp 1619617919
transform 1 0 6532 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1619617919
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1619617919
transform -1 0 8740 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen1
timestamp 1619617919
transform 1 0 8464 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_1_94
timestamp 1619617919
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_88
timestamp 1619617919
transform 1 0 9200 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1619617919
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1619617919
transform 1 0 8924 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _356_
timestamp 1619617919
transform -1 0 10028 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1619617919
transform 1 0 9476 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1619617919
transform 1 0 10028 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb0
timestamp 1619617919
transform 1 0 9936 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_1_108
timestamp 1619617919
transform 1 0 11040 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106
timestamp 1619617919
transform 1 0 10856 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101
timestamp 1619617919
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1619617919
transform 1 0 10580 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen0
timestamp 1619617919
transform 1 0 10580 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_1_115
timestamp 1619617919
transform 1 0 11684 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1619617919
transform 1 0 11868 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1619617919
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1619617919
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1619617919
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1619617919
transform -1 0 12052 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_121
timestamp 1619617919
transform 1 0 12236 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1619617919
transform -1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb1
timestamp 1619617919
transform -1 0 12696 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_1_131
timestamp 1619617919
transform 1 0 13156 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130
timestamp 1619617919
transform 1 0 13064 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen1
timestamp 1619617919
transform 1 0 12696 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1619617919
transform -1 0 13064 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1619617919
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_6  input1
timestamp 1619617919
transform 1 0 14536 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1619617919
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb0
timestamp 1619617919
transform -1 0 14352 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen0
timestamp 1619617919
transform -1 0 14444 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1619617919
transform -1 0 14720 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfrbp_1  idiv16
timestamp 1619617919
transform -1 0 16836 0 1 2720
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1619617919
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1619617919
transform 1 0 16560 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1619617919
transform 1 0 15364 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_159
timestamp 1619617919
transform 1 0 15732 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1619617919
transform 1 0 16468 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_171
timestamp 1619617919
transform 1 0 16836 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_172
timestamp 1619617919
transform 1 0 16928 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_175
timestamp 1619617919
transform 1 0 17204 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1619617919
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_188
timestamp 1619617919
transform 1 0 18400 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_184
timestamp 1619617919
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 1619617919
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output43
timestamp 1619617919
transform -1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1619617919
transform 1 0 18492 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1619617919
transform -1 0 18768 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1619617919
transform -1 0 19044 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1619617919
transform -1 0 19044 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1619617919
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1619617919
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1619617919
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrbp_2  idiv4
timestamp 1619617919
transform -1 0 6348 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1619617919
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1619617919
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_30
timestamp 1619617919
transform 1 0 3864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_57
timestamp 1619617919
transform 1 0 6348 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_69
timestamp 1619617919
transform 1 0 7452 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1619617919
transform -1 0 8372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1619617919
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_75
timestamp 1619617919
transform 1 0 8004 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_79
timestamp 1619617919
transform 1 0 8372 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1619617919
transform 1 0 8924 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_87
timestamp 1619617919
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_99
timestamp 1619617919
transform 1 0 10212 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1619617919
transform 1 0 10948 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_111
timestamp 1619617919
transform 1 0 11316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1619617919
transform 1 0 12420 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1619617919
transform 1 0 14352 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1619617919
transform 1 0 13892 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1619617919
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1619617919
transform 1 0 13524 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_142
timestamp 1619617919
transform 1 0 14168 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfrbp_2  idiv8
timestamp 1619617919
transform 1 0 15548 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_4  FILLER_2_153
timestamp 1619617919
transform 1 0 15180 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1619617919
transform -1 0 19044 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_181
timestamp 1619617919
transform 1 0 17756 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_189
timestamp 1619617919
transform 1 0 18492 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1619617919
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1619617919
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1619617919
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1619617919
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1619617919
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _368_
timestamp 1619617919
transform -1 0 7728 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb0
timestamp 1619617919
transform 1 0 7728 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1619617919
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1619617919
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_58
timestamp 1619617919
transform 1 0 6440 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_62
timestamp 1619617919
transform 1 0 6808 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1619617919
transform -1 0 10672 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_79
timestamp 1619617919
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_91
timestamp 1619617919
transform 1 0 9476 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp 1619617919
transform -1 0 12512 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb1
timestamp 1619617919
transform 1 0 12512 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1619617919
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1619617919
transform 1 0 10672 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_112
timestamp 1619617919
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1619617919
transform 1 0 13616 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen1
timestamp 1619617919
transform 1 0 13156 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_3_139
timestamp 1619617919
transform 1 0 13892 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1619617919
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_151
timestamp 1619617919
transform 1 0 14996 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_163
timestamp 1619617919
transform 1 0 16100 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_172
timestamp 1619617919
transform 1 0 16928 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1619617919
transform -1 0 19044 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_184
timestamp 1619617919
transform 1 0 18032 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1619617919
transform 1 0 3220 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  ringosc.ibufp11
timestamp 1619617919
transform -1 0 2484 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1619617919
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output41
timestamp 1619617919
transform -1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_7
timestamp 1619617919
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_11
timestamp 1619617919
transform 1 0 2116 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_15
timestamp 1619617919
transform 1 0 2484 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1619617919
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1619617919
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1619617919
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1619617919
transform 1 0 4968 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen0
timestamp 1619617919
transform 1 0 7268 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1619617919
transform -1 0 6624 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_54
timestamp 1619617919
transform 1 0 6072 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_60
timestamp 1619617919
transform 1 0 6624 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_66
timestamp 1619617919
transform 1 0 7176 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_72
timestamp 1619617919
transform 1 0 7728 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[11\].id.delayenb1
timestamp 1619617919
transform 1 0 10028 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1619617919
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1619617919
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_87
timestamp 1619617919
transform 1 0 9108 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_95
timestamp 1619617919
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1619617919
transform 1 0 11132 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[11\].id.delayen1
timestamp 1619617919
transform 1 0 10672 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__buf_8  repeater46
timestamp 1619617919
transform -1 0 12512 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_124
timestamp 1619617919
transform 1 0 12512 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1619617919
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_136
timestamp 1619617919
transform 1 0 13616 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_142
timestamp 1619617919
transform 1 0 14168 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_144
timestamp 1619617919
transform 1 0 14352 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1619617919
transform 1 0 16008 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1619617919
transform 1 0 14996 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_150
timestamp 1619617919
transform 1 0 14904 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_160
timestamp 1619617919
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_171
timestamp 1619617919
transform 1 0 16836 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1619617919
transform -1 0 19044 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1619617919
transform -1 0 18768 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_183
timestamp 1619617919
transform 1 0 17940 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__inv_1  ringosc.ibufp10
timestamp 1619617919
transform -1 0 3036 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1619617919
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1619617919
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp 1619617919
transform 1 0 2484 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_21
timestamp 1619617919
transform 1 0 3036 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[5\].id.delayen1
timestamp 1619617919
transform 1 0 5520 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[5\].id.delayenb1
timestamp 1619617919
transform -1 0 5520 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_5_33
timestamp 1619617919
transform 1 0 4140 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1619617919
transform 1 0 5980 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1619617919
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_56
timestamp 1619617919
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1619617919
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_70
timestamp 1619617919
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_82
timestamp 1619617919
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_94
timestamp 1619617919
transform 1 0 9752 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1619617919
transform -1 0 12788 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1619617919
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_106
timestamp 1619617919
transform 1 0 10856 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_115
timestamp 1619617919
transform 1 0 11684 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_127
timestamp 1619617919
transform 1 0 12788 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_139
timestamp 1619617919
transform 1 0 13892 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__nor3_2  _324_
timestamp 1619617919
transform -1 0 15824 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _325_
timestamp 1619617919
transform 1 0 15824 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1619617919
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_151
timestamp 1619617919
transform 1 0 14996 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_168
timestamp 1619617919
transform 1 0 16560 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_172
timestamp 1619617919
transform 1 0 16928 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1619617919
transform -1 0 19044 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_184
timestamp 1619617919
transform 1 0 18032 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1619617919
transform -1 0 3404 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1619617919
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1619617919
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1619617919
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_15
timestamp 1619617919
transform 1 0 2484 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1619617919
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1619617919
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1619617919
transform 1 0 4876 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb0
timestamp 1619617919
transform 1 0 3864 0 -1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1619617919
transform -1 0 5796 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1619617919
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_25
timestamp 1619617919
transform 1 0 3404 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1619617919
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1619617919
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1619617919
transform 1 0 6624 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0
timestamp 1619617919
transform 1 0 6532 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.delayen0
timestamp 1619617919
transform 1 0 6992 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1619617919
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_51
timestamp 1619617919
transform 1 0 5796 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_59
timestamp 1619617919
transform 1 0 6532 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_69
timestamp 1619617919
transform 1 0 7452 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1619617919
transform 1 0 5796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_58
timestamp 1619617919
transform 1 0 6440 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_75
timestamp 1619617919
transform 1 0 8004 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_80
timestamp 1619617919
transform 1 0 8464 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1619617919
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1619617919
transform -1 0 8464 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb0
timestamp 1619617919
transform 1 0 8096 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_7_97
timestamp 1619617919
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1619617919
transform 1 0 10212 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.iss.delayenb1
timestamp 1619617919
transform 1 0 9108 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1619617919
transform 1 0 9752 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_4  ringosc.dstage\[11\].id.delayen0
timestamp 1619617919
transform 1 0 10212 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_12  FILLER_6_87
timestamp 1619617919
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1619617919
transform 1 0 10672 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen0
timestamp 1619617919
transform 1 0 12328 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb0
timestamp 1619617919
transform 1 0 12052 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1619617919
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_103
timestamp 1619617919
transform 1 0 10580 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_107
timestamp 1619617919
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_110
timestamp 1619617919
transform 1 0 11224 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_115
timestamp 1619617919
transform 1 0 11684 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1619617919
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_2  _322_
timestamp 1619617919
transform -1 0 15364 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1619617919
transform -1 0 15180 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1619617919
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_126
timestamp 1619617919
transform 1 0 12696 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_138
timestamp 1619617919
transform 1 0 13800 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_142
timestamp 1619617919
transform 1 0 14168 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1619617919
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_139
timestamp 1619617919
transform 1 0 13892 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1619617919
transform -1 0 16192 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1619617919
transform 1 0 16192 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _323_
timestamp 1619617919
transform 1 0 15180 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1619617919
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_167
timestamp 1619617919
transform 1 0 16468 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_155
timestamp 1619617919
transform 1 0 15364 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_167
timestamp 1619617919
transform 1 0 16468 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_172
timestamp 1619617919
transform 1 0 16928 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1619617919
transform -1 0 19044 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1619617919
transform -1 0 19044 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_179
timestamp 1619617919
transform 1 0 17572 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_191
timestamp 1619617919
transform 1 0 18676 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_184
timestamp 1619617919
transform 1 0 18032 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _360_
timestamp 1619617919
transform -1 0 2576 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb0
timestamp 1619617919
transform 1 0 2576 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1619617919
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1619617919
transform -1 0 1656 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6
timestamp 1619617919
transform 1 0 1656 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_23
timestamp 1619617919
transform 1 0 3220 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _372_
timestamp 1619617919
transform -1 0 5428 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1619617919
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_30
timestamp 1619617919
transform 1 0 3864 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_47
timestamp 1619617919
transform 1 0 5428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _196_
timestamp 1619617919
transform 1 0 5704 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1
timestamp 1619617919
transform 1 0 7636 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.reseten0
timestamp 1619617919
transform 1 0 6624 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  FILLER_8_57
timestamp 1619617919
transform 1 0 6348 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_74
timestamp 1619617919
transform 1 0 7912 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb0
timestamp 1619617919
transform 1 0 9936 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.delayen1
timestamp 1619617919
transform 1 0 8372 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1619617919
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_78
timestamp 1619617919
transform 1 0 8280 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1619617919
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_87
timestamp 1619617919
transform 1 0 9108 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_95
timestamp 1619617919
transform 1 0 9844 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1619617919
transform -1 0 12512 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_107
timestamp 1619617919
transform 1 0 10948 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_124
timestamp 1619617919
transform 1 0 12512 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1619617919
transform 1 0 14352 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1619617919
transform -1 0 13892 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1619617919
transform -1 0 13432 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1619617919
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_130
timestamp 1619617919
transform 1 0 13064 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_134
timestamp 1619617919
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_139
timestamp 1619617919
transform 1 0 13892 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1619617919
transform -1 0 16652 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1619617919
transform 1 0 15180 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_169
timestamp 1619617919
transform 1 0 16652 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1619617919
transform -1 0 19044 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1619617919
transform 1 0 18492 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_181
timestamp 1619617919
transform 1 0 17756 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen0
timestamp 1619617919
transform 1 0 2116 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1619617919
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1619617919
transform 1 0 1380 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_16
timestamp 1619617919
transform 1 0 2576 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _303_
timestamp 1619617919
transform 1 0 3772 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_28
timestamp 1619617919
transform 1 0 3680 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_35
timestamp 1619617919
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1619617919
transform 1 0 5428 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_8  _197_
timestamp 1619617919
transform -1 0 7912 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1619617919
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_55
timestamp 1619617919
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1619617919
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1619617919
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_98
timestamp 1619617919
transform 1 0 10120 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _291_
timestamp 1619617919
transform 1 0 10948 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1619617919
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_106
timestamp 1619617919
transform 1 0 10856 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_112
timestamp 1619617919
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_115
timestamp 1619617919
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen1
timestamp 1619617919
transform 1 0 13432 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb1
timestamp 1619617919
transform 1 0 12788 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_9_139
timestamp 1619617919
transform 1 0 13892 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen0
timestamp 1619617919
transform 1 0 16376 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb0
timestamp 1619617919
transform 1 0 15732 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1619617919
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_151
timestamp 1619617919
transform 1 0 14996 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_172
timestamp 1619617919
transform 1 0 16928 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1619617919
transform -1 0 19044 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_184
timestamp 1619617919
transform 1 0 18032 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1619617919
transform 1 0 2484 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1619617919
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1619617919
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_18
timestamp 1619617919
transform 1 0 2760 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _354_
timestamp 1619617919
transform -1 0 4968 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1619617919
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_26
timestamp 1619617919
transform 1 0 3496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_30
timestamp 1619617919
transform 1 0 3864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1619617919
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00
timestamp 1619617919
transform -1 0 7912 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01
timestamp 1619617919
transform -1 0 7544 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_10_54
timestamp 1619617919
transform 1 0 6072 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_74
timestamp 1619617919
transform 1 0 7912 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _306_
timestamp 1619617919
transform 1 0 9108 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _321_
timestamp 1619617919
transform 1 0 8464 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1619617919
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_92
timestamp 1619617919
transform 1 0 9568 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0
timestamp 1619617919
transform 1 0 10764 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_104
timestamp 1619617919
transform 1 0 10672 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1619617919
transform 1 0 11132 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1619617919
transform 1 0 12236 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1619617919
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_133
timestamp 1619617919
transform 1 0 13340 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1619617919
transform 1 0 14076 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_144
timestamp 1619617919
transform 1 0 14352 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_156
timestamp 1619617919
transform 1 0 15456 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_168
timestamp 1619617919
transform 1 0 16560 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1619617919
transform -1 0 17664 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1619617919
transform -1 0 19044 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_176
timestamp 1619617919
transform 1 0 17296 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_180
timestamp 1619617919
transform 1 0 17664 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1619617919
transform 1 0 2760 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen1
timestamp 1619617919
transform 1 0 2300 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb1
timestamp 1619617919
transform 1 0 1656 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1619617919
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1619617919
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_21
timestamp 1619617919
transform 1 0 3036 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1619617919
transform 1 0 5336 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _377_
timestamp 1619617919
transform -1 0 4600 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_38
timestamp 1619617919
transform 1 0 4600 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1619617919
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_55
timestamp 1619617919
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1619617919
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_70
timestamp 1619617919
transform 1 0 7544 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _312_
timestamp 1619617919
transform -1 0 9752 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1619617919
transform -1 0 8924 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp 1619617919
transform 1 0 8924 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_94
timestamp 1619617919
transform 1 0 9752 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1619617919
transform 1 0 12144 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen1
timestamp 1619617919
transform 1 0 11684 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb1
timestamp 1619617919
transform 1 0 10856 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1619617919
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1619617919
transform 1 0 11500 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1619617919
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 1619617919
transform 1 0 12788 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb0
timestamp 1619617919
transform 1 0 14444 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_11_130
timestamp 1619617919
transform 1 0 13064 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_142
timestamp 1619617919
transform 1 0 14168 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen0
timestamp 1619617919
transform 1 0 15088 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1619617919
transform 1 0 16376 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb1
timestamp 1619617919
transform -1 0 17664 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1619617919
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_157
timestamp 1619617919
transform 1 0 15548 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_165
timestamp 1619617919
transform 1 0 16284 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_170
timestamp 1619617919
transform 1 0 16744 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_172
timestamp 1619617919
transform 1 0 16928 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1619617919
transform 1 0 18124 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen1
timestamp 1619617919
transform 1 0 17664 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1619617919
transform -1 0 19044 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_188
timestamp 1619617919
transform 1 0 18400 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1619617919
transform 1 0 2484 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1619617919
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output39
timestamp 1619617919
transform -1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_7
timestamp 1619617919
transform 1 0 1748 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_19
timestamp 1619617919
transform 1 0 2852 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _307_
timestamp 1619617919
transform 1 0 4876 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _314_
timestamp 1619617919
transform 1 0 3864 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1619617919
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1619617919
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_36
timestamp 1619617919
transform 1 0 4416 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_40
timestamp 1619617919
transform 1 0 4784 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_48
timestamp 1619617919
transform 1 0 5520 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1619617919
transform -1 0 7360 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _302_
timestamp 1619617919
transform 1 0 6624 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_64
timestamp 1619617919
transform 1 0 6992 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_68
timestamp 1619617919
transform 1 0 7360 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1619617919
transform 1 0 9108 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _315_
timestamp 1619617919
transform 1 0 9384 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _319_
timestamp 1619617919
transform 1 0 8280 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1619617919
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_76
timestamp 1619617919
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1619617919
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_95
timestamp 1619617919
transform 1 0 9844 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1619617919
transform -1 0 11776 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb0
timestamp 1619617919
transform -1 0 13156 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_116
timestamp 1619617919
transform 1 0 11776 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen0
timestamp 1619617919
transform -1 0 13616 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1619617919
transform 1 0 14352 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1619617919
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_136
timestamp 1619617919
transform 1 0 13616 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_142
timestamp 1619617919
transform 1 0 14168 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_148
timestamp 1619617919
transform 1 0 14720 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_160
timestamp 1619617919
transform 1 0 15824 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_172
timestamp 1619617919
transform 1 0 16928 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1619617919
transform -1 0 19044 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_184
timestamp 1619617919
transform 1 0 18032 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_11
timestamp 1619617919
transform 1 0 2116 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1619617919
transform 1 0 1380 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1619617919
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1619617919
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1619617919
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb1
timestamp 1619617919
transform 1 0 2208 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1619617919
transform -1 0 2300 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen1
timestamp 1619617919
transform 1 0 2852 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1619617919
transform 1 0 3312 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_13
timestamp 1619617919
transform 1 0 2300 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_30
timestamp 1619617919
transform 1 0 3864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1619617919
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_33
timestamp 1619617919
transform 1 0 4140 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_25
timestamp 1619617919
transform 1 0 3404 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1619617919
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _366_
timestamp 1619617919
transform 1 0 4140 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _308_
timestamp 1619617919
transform 1 0 4416 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _304_
timestamp 1619617919
transform 1 0 4968 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _296_
timestamp 1619617919
transform -1 0 5520 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_14_49
timestamp 1619617919
transform 1 0 5612 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_48
timestamp 1619617919
transform 1 0 5520 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_57
timestamp 1619617919
transform 1 0 6348 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_58
timestamp 1619617919
transform 1 0 6440 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1619617919
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _301_
timestamp 1619617919
transform 1 0 6532 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _300_
timestamp 1619617919
transform -1 0 6900 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1619617919
transform 1 0 6072 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_63
timestamp 1619617919
transform 1 0 6900 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__a31o_1  _298_
timestamp 1619617919
transform -1 0 7728 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_14_63
timestamp 1619617919
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_72
timestamp 1619617919
transform 1 0 7728 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_4  _311_
timestamp 1619617919
transform 1 0 9108 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _317_
timestamp 1619617919
transform -1 0 10488 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1619617919
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_84
timestamp 1619617919
transform 1 0 8832 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_96
timestamp 1619617919
transform 1 0 9936 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_75
timestamp 1619617919
transform 1 0 8004 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_83
timestamp 1619617919
transform 1 0 8740 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _365_
timestamp 1619617919
transform 1 0 10764 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1619617919
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_108
timestamp 1619617919
transform 1 0 11040 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_115
timestamp 1619617919
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_102
timestamp 1619617919
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_114
timestamp 1619617919
transform 1 0 11592 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_122
timestamp 1619617919
transform 1 0 12328 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _347_
timestamp 1619617919
transform -1 0 12880 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _357_
timestamp 1619617919
transform 1 0 12880 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb1
timestamp 1619617919
transform -1 0 15088 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1619617919
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_127
timestamp 1619617919
transform 1 0 12788 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_139
timestamp 1619617919
transform 1 0 13892 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_137
timestamp 1619617919
transform 1 0 13708 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_144
timestamp 1619617919
transform 1 0 14352 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_161
timestamp 1619617919
transform 1 0 15916 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_155
timestamp 1619617919
transform 1 0 15364 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_151
timestamp 1619617919
transform 1 0 14996 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1619617919
transform 1 0 15732 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1619617919
transform 1 0 15456 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp 1619617919
transform 1 0 15088 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_169
timestamp 1619617919
transform 1 0 16652 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_170
timestamp 1619617919
transform 1 0 16744 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_162
timestamp 1619617919
transform 1 0 16008 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1619617919
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _373_
timestamp 1619617919
transform -1 0 17572 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1619617919
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1619617919
transform -1 0 19044 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1619617919
transform -1 0 19044 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1619617919
transform 1 0 18492 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_184
timestamp 1619617919
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_188
timestamp 1619617919
transform 1 0 18400 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_179
timestamp 1619617919
transform 1 0 17572 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_191
timestamp 1619617919
transform 1 0 18676 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1619617919
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1619617919
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1619617919
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _248_
timestamp 1619617919
transform 1 0 4600 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_15_27
timestamp 1619617919
transform 1 0 3588 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_35
timestamp 1619617919
transform 1 0 4324 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_43
timestamp 1619617919
transform 1 0 5060 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1619617919
transform 1 0 7176 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1619617919
transform 1 0 6072 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _254_
timestamp 1619617919
transform 1 0 6440 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1619617919
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_51
timestamp 1619617919
transform 1 0 5796 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_65
timestamp 1619617919
transform 1 0 7084 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_69
timestamp 1619617919
transform 1 0 7452 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1619617919
transform -1 0 9200 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _309_
timestamp 1619617919
transform 1 0 8464 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _310_
timestamp 1619617919
transform -1 0 8464 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _316_
timestamp 1619617919
transform -1 0 10028 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_97
timestamp 1619617919
transform 1 0 10028 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _292_
timestamp 1619617919
transform 1 0 12420 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _313_
timestamp 1619617919
transform -1 0 10764 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _318_
timestamp 1619617919
transform -1 0 12144 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1619617919
transform -1 0 11592 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1619617919
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_101
timestamp 1619617919
transform 1 0 10396 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_120
timestamp 1619617919
transform 1 0 12144 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1619617919
transform 1 0 12972 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_128
timestamp 1619617919
transform 1 0 12880 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_138
timestamp 1619617919
transform 1 0 13800 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen1
timestamp 1619617919
transform 1 0 14996 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1619617919
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_150
timestamp 1619617919
transform 1 0 14904 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_156
timestamp 1619617919
transform 1 0 15456 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_168
timestamp 1619617919
transform 1 0 16560 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_172
timestamp 1619617919
transform 1 0 16928 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1619617919
transform -1 0 19044 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_184
timestamp 1619617919
transform 1 0 18032 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1619617919
transform 1 0 2760 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1619617919
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1619617919
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_15
timestamp 1619617919
transform 1 0 2484 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_21
timestamp 1619617919
transform 1 0 3036 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1619617919
transform 1 0 5060 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _293_
timestamp 1619617919
transform -1 0 4600 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1619617919
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_30
timestamp 1619617919
transform 1 0 3864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_38
timestamp 1619617919
transform 1 0 4600 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_42
timestamp 1619617919
transform 1 0 4968 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_46
timestamp 1619617919
transform 1 0 5336 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _294_
timestamp 1619617919
transform 1 0 6072 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_16_59
timestamp 1619617919
transform 1 0 6532 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_71
timestamp 1619617919
transform 1 0 7636 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1619617919
transform 1 0 8096 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1619617919
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_75
timestamp 1619617919
transform 1 0 8004 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_79
timestamp 1619617919
transform 1 0 8372 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1619617919
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_87
timestamp 1619617919
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_99
timestamp 1619617919
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  _290_
timestamp 1619617919
transform 1 0 10396 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _371_
timestamp 1619617919
transform -1 0 11868 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_106
timestamp 1619617919
transform 1 0 10856 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1619617919
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1619617919
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_129
timestamp 1619617919
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1619617919
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_144
timestamp 1619617919
transform 1 0 14352 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _385_
timestamp 1619617919
transform 1 0 16100 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_16_156
timestamp 1619617919
transform 1 0 15456 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_162
timestamp 1619617919
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1619617919
transform -1 0 19044 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_184
timestamp 1619617919
transform 1 0 18032 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _364_
timestamp 1619617919
transform -1 0 2300 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen0
timestamp 1619617919
transform -1 0 3404 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb0
timestamp 1619617919
transform 1 0 2300 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1619617919
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1619617919
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _305_
timestamp 1619617919
transform 1 0 4508 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1619617919
transform 1 0 5152 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_25
timestamp 1619617919
transform 1 0 3404 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1619617919
transform 1 0 5428 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _394_
timestamp 1619617919
transform 1 0 6624 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1619617919
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_55
timestamp 1619617919
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_58
timestamp 1619617919
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__o41a_1  _320_
timestamp 1619617919
transform -1 0 9936 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_17_81
timestamp 1619617919
transform 1 0 8556 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_96
timestamp 1619617919
transform 1 0 9936 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _401_
timestamp 1619617919
transform 1 0 12328 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1619617919
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_108
timestamp 1619617919
transform 1 0 11040 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_115
timestamp 1619617919
transform 1 0 11684 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1619617919
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _386_
timestamp 1619617919
transform -1 0 16284 0 1 11424
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1619617919
transform -1 0 17296 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1619617919
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_165
timestamp 1619617919
transform 1 0 16284 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_172
timestamp 1619617919
transform 1 0 16928 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1619617919
transform -1 0 18216 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1619617919
transform -1 0 19044 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1619617919
transform -1 0 18768 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_176
timestamp 1619617919
transform 1 0 17296 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1619617919
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_186
timestamp 1619617919
transform 1 0 18216 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1619617919
transform -1 0 3220 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1619617919
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output40
timestamp 1619617919
transform -1 0 1748 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_7
timestamp 1619617919
transform 1 0 1748 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_23
timestamp 1619617919
transform 1 0 3220 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_2  _392_
timestamp 1619617919
transform 1 0 4048 0 -1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1619617919
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_30
timestamp 1619617919
transform 1 0 3864 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1619617919
transform 1 0 6164 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp 1619617919
transform -1 0 7728 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_53
timestamp 1619617919
transform 1 0 5980 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_58
timestamp 1619617919
transform 1 0 6440 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_66
timestamp 1619617919
transform 1 0 7176 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_72
timestamp 1619617919
transform 1 0 7728 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1619617919
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1619617919
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1619617919
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_99
timestamp 1619617919
transform 1 0 10212 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1619617919
transform 1 0 10488 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _199_
timestamp 1619617919
transform -1 0 13156 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1619617919
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_117
timestamp 1619617919
transform 1 0 11868 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_123
timestamp 1619617919
transform 1 0 12420 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1619617919
transform -1 0 13616 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1619617919
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_131
timestamp 1619617919
transform 1 0 13156 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_136
timestamp 1619617919
transform 1 0 13616 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_142
timestamp 1619617919
transform 1 0 14168 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_144
timestamp 1619617919
transform 1 0 14352 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _341_
timestamp 1619617919
transform 1 0 15088 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _400_
timestamp 1619617919
transform 1 0 16928 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_18_155
timestamp 1619617919
transform 1 0 15364 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_167
timestamp 1619617919
transform 1 0 16468 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_171
timestamp 1619617919
transform 1 0 16836 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1619617919
transform -1 0 19044 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1619617919
transform 1 0 1472 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen1
timestamp 1619617919
transform 1 0 3220 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb1
timestamp 1619617919
transform -1 0 3220 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1619617919
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1619617919
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1619617919
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1619617919
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1619617919
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_13
timestamp 1619617919
transform 1 0 2300 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _246_
timestamp 1619617919
transform 1 0 5152 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _273_
timestamp 1619617919
transform -1 0 5152 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1619617919
transform 1 0 3864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1619617919
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1619617919
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_39
timestamp 1619617919
transform 1 0 4692 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_28
timestamp 1619617919
transform 1 0 3680 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_33
timestamp 1619617919
transform 1 0 4140 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_45
timestamp 1619617919
transform 1 0 5244 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _252_
timestamp 1619617919
transform 1 0 7452 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _266_
timestamp 1619617919
transform -1 0 7360 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1619617919
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_51
timestamp 1619617919
transform 1 0 5796 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_58
timestamp 1619617919
transform 1 0 6440 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_68
timestamp 1619617919
transform 1 0 7360 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_57
timestamp 1619617919
transform 1 0 6348 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_69
timestamp 1619617919
transform 1 0 7452 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _258_
timestamp 1619617919
transform -1 0 9752 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _261_
timestamp 1619617919
transform -1 0 10120 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _363_
timestamp 1619617919
transform 1 0 8832 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _395_
timestamp 1619617919
transform 1 0 10120 0 -1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1619617919
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_76
timestamp 1619617919
transform 1 0 8096 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1619617919
transform 1 0 9660 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_81
timestamp 1619617919
transform 1 0 8556 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1619617919
transform 1 0 8924 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  _194_
timestamp 1619617919
transform 1 0 11684 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _212_
timestamp 1619617919
transform 1 0 12512 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1619617919
transform -1 0 11408 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1619617919
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_105
timestamp 1619617919
transform 1 0 10764 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1619617919
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_122
timestamp 1619617919
transform 1 0 12328 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_119
timestamp 1619617919
transform 1 0 12052 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_123
timestamp 1619617919
transform 1 0 12420 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _207_
timestamp 1619617919
transform 1 0 13616 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _223_
timestamp 1619617919
transform 1 0 13248 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _285_
timestamp 1619617919
transform 1 0 14352 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _286_
timestamp 1619617919
transform -1 0 15364 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1619617919
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_134
timestamp 1619617919
transform 1 0 13432 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_146
timestamp 1619617919
transform 1 0 14536 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_139
timestamp 1619617919
transform 1 0 13892 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1619617919
transform 1 0 15088 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _200_
timestamp 1619617919
transform 1 0 16928 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _287_
timestamp 1619617919
transform 1 0 15548 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _288_
timestamp 1619617919
transform 1 0 16376 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1619617919
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_155
timestamp 1619617919
transform 1 0 15364 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_167
timestamp 1619617919
transform 1 0 16468 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_155
timestamp 1619617919
transform 1 0 15364 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_171
timestamp 1619617919
transform 1 0 16836 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _209_
timestamp 1619617919
transform 1 0 17480 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1619617919
transform -1 0 19044 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1619617919
transform -1 0 19044 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_179
timestamp 1619617919
transform 1 0 17572 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_191
timestamp 1619617919
transform 1 0 18676 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_177
timestamp 1619617919
transform 1 0 17388 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_186
timestamp 1619617919
transform 1 0 18216 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1619617919
transform 1 0 2024 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1619617919
transform -1 0 3128 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1619617919
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1619617919
transform -1 0 1656 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_6
timestamp 1619617919
transform 1 0 1656 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_17
timestamp 1619617919
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_22
timestamp 1619617919
transform 1 0 3128 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1619617919
transform 1 0 5428 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _272_
timestamp 1619617919
transform -1 0 5428 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_34
timestamp 1619617919
transform 1 0 4232 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_38
timestamp 1619617919
transform 1 0 4600 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1619617919
transform -1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _265_
timestamp 1619617919
transform -1 0 7728 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1619617919
transform 1 0 5704 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1619617919
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_53
timestamp 1619617919
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_58
timestamp 1619617919
transform 1 0 6440 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1619617919
transform 1 0 9660 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1619617919
transform 1 0 9936 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _260_
timestamp 1619617919
transform 1 0 8924 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_75
timestamp 1619617919
transform 1 0 8004 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1619617919
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_99
timestamp 1619617919
transform 1 0 10212 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1619617919
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_111
timestamp 1619617919
transform 1 0 11316 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_115
timestamp 1619617919
transform 1 0 11684 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1619617919
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1619617919
transform -1 0 13616 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _224_
timestamp 1619617919
transform 1 0 12604 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1619617919
transform -1 0 15088 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_136
timestamp 1619617919
transform 1 0 13616 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_148
timestamp 1619617919
transform 1 0 14720 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1619617919
transform -1 0 16192 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1619617919
transform 1 0 16284 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _279_
timestamp 1619617919
transform -1 0 15548 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1619617919
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_157
timestamp 1619617919
transform 1 0 15548 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_164
timestamp 1619617919
transform 1 0 16192 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_168
timestamp 1619617919
transform 1 0 16560 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_172
timestamp 1619617919
transform 1 0 16928 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _210_
timestamp 1619617919
transform -1 0 17848 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1619617919
transform -1 0 19044 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1619617919
transform -1 0 18768 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_182
timestamp 1619617919
transform 1 0 17848 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_188
timestamp 1619617919
transform 1 0 18400 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb0
timestamp 1619617919
transform 1 0 1472 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1619617919
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1619617919
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_11
timestamp 1619617919
transform 1 0 2116 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_23
timestamp 1619617919
transform 1 0 3220 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _250_
timestamp 1619617919
transform -1 0 5888 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _270_
timestamp 1619617919
transform -1 0 5152 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1619617919
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_30
timestamp 1619617919
transform 1 0 3864 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_38
timestamp 1619617919
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__o32a_1  _256_
timestamp 1619617919
transform -1 0 8372 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _263_
timestamp 1619617919
transform 1 0 6992 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1619617919
transform 1 0 7360 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_52
timestamp 1619617919
transform 1 0 5888 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1619617919
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_79
timestamp 1619617919
transform 1 0 8372 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1619617919
transform 1 0 8924 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_87
timestamp 1619617919
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_99
timestamp 1619617919
transform 1 0 10212 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _220_
timestamp 1619617919
transform 1 0 10948 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_115
timestamp 1619617919
transform 1 0 11684 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1619617919
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_127
timestamp 1619617919
transform 1 0 12788 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_139
timestamp 1619617919
transform 1 0 13892 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_144
timestamp 1619617919
transform 1 0 14352 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__o2bb2ai_1  _228_
timestamp 1619617919
transform -1 0 17388 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1619617919
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_168
timestamp 1619617919
transform 1 0 16560 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1619617919
transform -1 0 19044 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1619617919
transform 1 0 17388 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_189
timestamp 1619617919
transform 1 0 18492 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1619617919
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1619617919
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1619617919
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _244_
timestamp 1619617919
transform 1 0 4692 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _269_
timestamp 1619617919
transform -1 0 5796 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1619617919
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _251_
timestamp 1619617919
transform 1 0 7268 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _262_
timestamp 1619617919
transform -1 0 8372 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1619617919
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_51
timestamp 1619617919
transform 1 0 5796 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_58
timestamp 1619617919
transform 1 0 6440 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_66
timestamp 1619617919
transform 1 0 7176 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _222_
timestamp 1619617919
transform -1 0 10396 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_79
timestamp 1619617919
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_91
timestamp 1619617919
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _206_
timestamp 1619617919
transform 1 0 12236 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _219_
timestamp 1619617919
transform 1 0 11684 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _221_
timestamp 1619617919
transform -1 0 10856 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1619617919
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_106
timestamp 1619617919
transform 1 0 10856 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_124
timestamp 1619617919
transform 1 0 12512 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _284_
timestamp 1619617919
transform 1 0 14444 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_23_136
timestamp 1619617919
transform 1 0 13616 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_144
timestamp 1619617919
transform 1 0 14352 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _208_
timestamp 1619617919
transform 1 0 16928 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1619617919
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_152
timestamp 1619617919
transform 1 0 15088 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_164
timestamp 1619617919
transform 1 0 16192 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_170
timestamp 1619617919
transform 1 0 16744 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1619617919
transform -1 0 19044 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_177
timestamp 1619617919
transform 1 0 17388 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_189
timestamp 1619617919
transform 1 0 18492 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _391_
timestamp 1619617919
transform 1 0 1840 0 -1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1619617919
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1619617919
transform -1 0 1656 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_6
timestamp 1619617919
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1619617919
transform 1 0 5152 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1619617919
transform 1 0 5428 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _274_
timestamp 1619617919
transform -1 0 5060 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _275_
timestamp 1619617919
transform 1 0 3864 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1619617919
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_43
timestamp 1619617919
transform 1 0 5060 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _267_
timestamp 1619617919
transform -1 0 7728 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_50
timestamp 1619617919
transform 1 0 5704 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_62
timestamp 1619617919
transform 1 0 6808 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_68
timestamp 1619617919
transform 1 0 7360 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_72
timestamp 1619617919
transform 1 0 7728 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1619617919
transform 1 0 9476 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1619617919
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1619617919
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_87
timestamp 1619617919
transform 1 0 9108 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_94
timestamp 1619617919
transform 1 0 9752 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__o2bb2a_1  _213_
timestamp 1619617919
transform -1 0 11960 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _402_
timestamp 1619617919
transform -1 0 13800 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_24_106
timestamp 1619617919
transform 1 0 10856 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _384_
timestamp 1619617919
transform 1 0 14352 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1619617919
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_138
timestamp 1619617919
transform 1 0 13800 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_142
timestamp 1619617919
transform 1 0 14168 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _201_
timestamp 1619617919
transform 1 0 16560 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_24_164
timestamp 1619617919
transform 1 0 16192 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1619617919
transform -1 0 18032 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _227_
timestamp 1619617919
transform 1 0 17204 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1619617919
transform -1 0 19044 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1619617919
transform 1 0 18492 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_184
timestamp 1619617919
transform 1 0 18032 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_188
timestamp 1619617919
transform 1 0 18400 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1619617919
transform -1 0 3036 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1619617919
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1619617919
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_15
timestamp 1619617919
transform 1 0 2484 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_21
timestamp 1619617919
transform 1 0 3036 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_33
timestamp 1619617919
transform 1 0 4140 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_45
timestamp 1619617919
transform 1 0 5244 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_1  _268_
timestamp 1619617919
transform 1 0 6900 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1619617919
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_58
timestamp 1619617919
transform 1 0 6440 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_62
timestamp 1619617919
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_71
timestamp 1619617919
transform 1 0 7636 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a221oi_2  _226_
timestamp 1619617919
transform 1 0 9200 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1619617919
transform 1 0 8740 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_87
timestamp 1619617919
transform 1 0 9108 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _198_
timestamp 1619617919
transform 1 0 11868 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1619617919
transform -1 0 11040 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _237_
timestamp 1619617919
transform 1 0 10304 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1619617919
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_108
timestamp 1619617919
transform 1 0 11040 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_115
timestamp 1619617919
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_124
timestamp 1619617919
transform 1 0 12512 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a311o_1  _289_
timestamp 1619617919
transform 1 0 14260 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_136
timestamp 1619617919
transform 1 0 13616 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_142
timestamp 1619617919
transform 1 0 14168 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _343_
timestamp 1619617919
transform -1 0 15272 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _399_
timestamp 1619617919
transform 1 0 16928 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1619617919
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_154
timestamp 1619617919
transform 1 0 15272 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_166
timestamp 1619617919
transform 1 0 16376 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_170
timestamp 1619617919
transform 1 0 16744 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1619617919
transform -1 0 19044 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _390_
timestamp 1619617919
transform 1 0 1564 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1619617919
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1619617919
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1619617919
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1619617919
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1619617919
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_30
timestamp 1619617919
transform 1 0 3864 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1619617919
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1619617919
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1619617919
transform 1 0 3404 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _277_
timestamp 1619617919
transform 1 0 3680 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_38
timestamp 1619617919
transform 1 0 4600 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _242_
timestamp 1619617919
transform -1 0 5060 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _240_
timestamp 1619617919
transform 1 0 4416 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_27_46
timestamp 1619617919
transform 1 0 5336 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_49
timestamp 1619617919
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_43
timestamp 1619617919
transform 1 0 5060 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1619617919
transform 1 0 5060 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1619617919
transform 1 0 5704 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1619617919
transform -1 0 7636 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _393_
timestamp 1619617919
transform 1 0 6532 0 -1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1619617919
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_53
timestamp 1619617919
transform 1 0 5980 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_54
timestamp 1619617919
transform 1 0 6072 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_58
timestamp 1619617919
transform 1 0 6440 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_66
timestamp 1619617919
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_71
timestamp 1619617919
transform 1 0 7636 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__a41o_2  _234_
timestamp 1619617919
transform 1 0 9292 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _236_
timestamp 1619617919
transform -1 0 10488 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_4  _238_
timestamp 1619617919
transform 1 0 9476 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1619617919
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_80
timestamp 1619617919
transform 1 0 8464 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1619617919
transform 1 0 9108 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_83
timestamp 1619617919
transform 1 0 8740 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _214_
timestamp 1619617919
transform 1 0 11684 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1619617919
transform -1 0 10764 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1619617919
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_108
timestamp 1619617919
transform 1 0 11040 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_120
timestamp 1619617919
transform 1 0 12144 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_105
timestamp 1619617919
transform 1 0 10764 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1619617919
transform 1 0 11500 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_120
timestamp 1619617919
transform 1 0 12144 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1619617919
transform -1 0 13524 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _387_
timestamp 1619617919
transform 1 0 13524 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1619617919
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_132
timestamp 1619617919
transform 1 0 13248 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_140
timestamp 1619617919
transform 1 0 13984 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1619617919
transform 1 0 14352 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _229_
timestamp 1619617919
transform 1 0 16928 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1619617919
transform -1 0 16652 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _231_
timestamp 1619617919
transform -1 0 17204 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _232_
timestamp 1619617919
transform 1 0 15824 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1619617919
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_156
timestamp 1619617919
transform 1 0 15456 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_164
timestamp 1619617919
transform 1 0 16192 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_156
timestamp 1619617919
transform 1 0 15456 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1619617919
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_183
timestamp 1619617919
transform 1 0 17940 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_175
timestamp 1619617919
transform 1 0 17204 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1619617919
transform 1 0 18032 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_191
timestamp 1619617919
transform 1 0 18676 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_187
timestamp 1619617919
transform 1 0 18308 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_191
timestamp 1619617919
transform 1 0 18676 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1619617919
transform 1 0 18308 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1619617919
transform -1 0 19044 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1619617919
transform -1 0 19044 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_175
timestamp 1619617919
transform 1 0 17204 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1619617919
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1619617919
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_6
timestamp 1619617919
transform 1 0 1656 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_18
timestamp 1619617919
transform 1 0 2760 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _241_
timestamp 1619617919
transform -1 0 4968 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _276_
timestamp 1619617919
transform -1 0 4692 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1619617919
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_26
timestamp 1619617919
transform 1 0 3496 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_30
timestamp 1619617919
transform 1 0 3864 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_42
timestamp 1619617919
transform 1 0 4968 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1619617919
transform -1 0 6716 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_54
timestamp 1619617919
transform 1 0 6072 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_61
timestamp 1619617919
transform 1 0 6716 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_73
timestamp 1619617919
transform 1 0 7820 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1619617919
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 1619617919
transform 1 0 8924 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_87
timestamp 1619617919
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_99
timestamp 1619617919
transform 1 0 10212 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _215_
timestamp 1619617919
transform -1 0 12880 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _216_
timestamp 1619617919
transform -1 0 12144 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _218_
timestamp 1619617919
transform -1 0 11316 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_107
timestamp 1619617919
transform 1 0 10948 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _283_
timestamp 1619617919
transform 1 0 13156 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp 1619617919
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1619617919
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_128
timestamp 1619617919
transform 1 0 12880 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_140
timestamp 1619617919
transform 1 0 13984 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_144
timestamp 1619617919
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_149
timestamp 1619617919
transform 1 0 14812 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_161
timestamp 1619617919
transform 1 0 15916 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_173
timestamp 1619617919
transform 1 0 17020 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1619617919
transform -1 0 19044 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_185
timestamp 1619617919
transform 1 0 18124 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_191
timestamp 1619617919
transform 1 0 18676 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1619617919
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1619617919
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1619617919
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1619617919
transform 1 0 4692 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1619617919
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_42
timestamp 1619617919
transform 1 0 4968 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _398_
timestamp 1619617919
transform 1 0 6440 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1619617919
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_54
timestamp 1619617919
transform 1 0 6072 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_2  _233_
timestamp 1619617919
transform 1 0 8280 0 1 17952
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_29_88
timestamp 1619617919
transform 1 0 9200 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1619617919
transform -1 0 12788 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _205_
timestamp 1619617919
transform 1 0 11684 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1619617919
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_100
timestamp 1619617919
transform 1 0 10304 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_112
timestamp 1619617919
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_122
timestamp 1619617919
transform 1 0 12328 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_1  _282_
timestamp 1619617919
transform 1 0 12788 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_131
timestamp 1619617919
transform 1 0 13156 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_143
timestamp 1619617919
transform 1 0 14260 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _383_
timestamp 1619617919
transform 1 0 16928 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1619617919
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_155
timestamp 1619617919
transform 1 0 15364 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_167
timestamp 1619617919
transform 1 0 16468 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1619617919
transform -1 0 19044 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _338_
timestamp 1619617919
transform -1 0 3496 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1619617919
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1619617919
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_15
timestamp 1619617919
transform 1 0 2484 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1619617919
transform -1 0 4784 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _278_
timestamp 1619617919
transform 1 0 3864 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1619617919
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_26
timestamp 1619617919
transform 1 0 3496 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_40
timestamp 1619617919
transform 1 0 4784 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_48
timestamp 1619617919
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _202_
timestamp 1619617919
transform -1 0 8280 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 1619617919
transform 1 0 5704 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1619617919
transform 1 0 5980 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_65
timestamp 1619617919
transform 1 0 7084 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _203_
timestamp 1619617919
transform 1 0 8280 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1619617919
transform 1 0 9108 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1619617919
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1619617919
transform 1 0 8924 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_90
timestamp 1619617919
transform 1 0 9384 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_98
timestamp 1619617919
transform 1 0 10120 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1619617919
transform -1 0 12144 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _195_
timestamp 1619617919
transform -1 0 11868 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp 1619617919
transform -1 0 10672 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_104
timestamp 1619617919
transform 1 0 10672 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_120
timestamp 1619617919
transform 1 0 12144 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _339_
timestamp 1619617919
transform -1 0 13892 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _381_
timestamp 1619617919
transform 1 0 14444 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1619617919
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_132
timestamp 1619617919
transform 1 0 13248 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_139
timestamp 1619617919
transform 1 0 13892 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_144
timestamp 1619617919
transform 1 0 14352 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _382_
timestamp 1619617919
transform 1 0 16284 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp 1619617919
transform 1 0 18124 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1619617919
transform -1 0 19044 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output42
timestamp 1619617919
transform 1 0 18400 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _349_
timestamp 1619617919
transform 1 0 1656 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _389_
timestamp 1619617919
transform 1 0 2392 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1619617919
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1619617919
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_9
timestamp 1619617919
transform 1 0 1932 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_13
timestamp 1619617919
transform 1 0 2300 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _396_
timestamp 1619617919
transform 1 0 4508 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_31_34
timestamp 1619617919
transform 1 0 4232 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _204_
timestamp 1619617919
transform -1 0 7360 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _397_
timestamp 1619617919
transform -1 0 9568 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1619617919
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_58
timestamp 1619617919
transform 1 0 6440 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_62
timestamp 1619617919
transform 1 0 6808 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_68
timestamp 1619617919
transform 1 0 7360 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _403_
timestamp 1619617919
transform 1 0 9660 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_31_92
timestamp 1619617919
transform 1 0 9568 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1619617919
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 1619617919
transform 1 0 11500 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_115
timestamp 1619617919
transform 1 0 11684 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _388_
timestamp 1619617919
transform 1 0 12788 0 1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_31_148
timestamp 1619617919
transform 1 0 14720 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _345_
timestamp 1619617919
transform -1 0 16836 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp 1619617919
transform -1 0 15548 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1619617919
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_157
timestamp 1619617919
transform 1 0 15548 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1619617919
transform 1 0 16284 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_172
timestamp 1619617919
transform 1 0 16928 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _193_
timestamp 1619617919
transform -1 0 18768 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1619617919
transform -1 0 19044 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1619617919
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1619617919
transform 1 0 2300 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1619617919
transform -1 0 2024 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output44
timestamp 1619617919
transform -1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_10
timestamp 1619617919
transform 1 0 2024 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_16
timestamp 1619617919
transform 1 0 2576 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1619617919
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1619617919
transform 1 0 3864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1619617919
transform 1 0 5520 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_28
timestamp 1619617919
transform 1 0 3680 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_33
timestamp 1619617919
transform 1 0 4140 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_45
timestamp 1619617919
transform 1 0 5244 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1619617919
transform 1 0 6440 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1619617919
transform 1 0 6900 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_51
timestamp 1619617919
transform 1 0 5796 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_57
timestamp 1619617919
transform 1 0 6348 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_59
timestamp 1619617919
transform 1 0 6532 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_66
timestamp 1619617919
transform 1 0 7176 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1619617919
transform 1 0 9108 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1619617919
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1619617919
transform 1 0 8280 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_81
timestamp 1619617919
transform 1 0 8556 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_88
timestamp 1619617919
transform 1 0 9200 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_92
timestamp 1619617919
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_96
timestamp 1619617919
transform 1 0 9936 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1619617919
transform 1 0 11776 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1619617919
transform -1 0 11776 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_108
timestamp 1619617919
transform 1 0 11040 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_112
timestamp 1619617919
transform 1 0 11408 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_117
timestamp 1619617919
transform 1 0 11868 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1619617919
transform 1 0 14444 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1619617919
transform 1 0 12880 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1619617919
transform 1 0 14536 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_125
timestamp 1619617919
transform 1 0 12604 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_131
timestamp 1619617919
transform 1 0 13156 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_143
timestamp 1619617919
transform 1 0 14260 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_149
timestamp 1619617919
transform 1 0 14812 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1619617919
transform 1 0 15640 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_157
timestamp 1619617919
transform 1 0 15548 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_161
timestamp 1619617919
transform 1 0 15916 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_173
timestamp 1619617919
transform 1 0 17020 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1619617919
transform -1 0 19044 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1619617919
transform 1 0 17112 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1619617919
transform 1 0 17480 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1619617919
transform -1 0 18400 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1619617919
transform -1 0 18768 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_175
timestamp 1619617919
transform 1 0 17204 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_181
timestamp 1619617919
transform 1 0 17756 0 -1 20128
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 8848 800 8968 6 clockc
port 0 nsew signal tristate
rlabel metal3 s 0 11568 800 11688 6 clockd[0]
port 1 nsew signal tristate
rlabel metal3 s 0 4768 800 4888 6 clockd[1]
port 2 nsew signal tristate
rlabel metal3 s 19396 18368 20196 18488 6 clockd[2]
port 3 nsew signal tristate
rlabel metal2 s 17958 0 18014 800 6 clockd[3]
port 4 nsew signal tristate
rlabel metal3 s 0 20408 800 20528 6 clockp[0]
port 5 nsew signal tristate
rlabel metal2 s 1858 0 1914 800 6 clockp[1]
port 6 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 dco
port 7 nsew signal input
rlabel metal3 s 19396 13608 20196 13728 6 div[0]
port 8 nsew signal input
rlabel metal2 s 17498 21540 17554 22340 6 div[1]
port 9 nsew signal input
rlabel metal2 s 6918 21540 6974 22340 6 div[2]
port 10 nsew signal input
rlabel metal2 s 478 0 534 800 6 div[3]
port 11 nsew signal input
rlabel metal2 s 12898 21540 12954 22340 6 div[4]
port 12 nsew signal input
rlabel metal2 s 14278 21540 14334 22340 6 ext_trim[0]
port 13 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 ext_trim[10]
port 14 nsew signal input
rlabel metal2 s 2318 21540 2374 22340 6 ext_trim[11]
port 15 nsew signal input
rlabel metal3 s 19396 4768 20196 4888 6 ext_trim[12]
port 16 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 ext_trim[13]
port 17 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 ext_trim[14]
port 18 nsew signal input
rlabel metal3 s 19396 15648 20196 15768 6 ext_trim[15]
port 19 nsew signal input
rlabel metal2 s 3698 21540 3754 22340 6 ext_trim[16]
port 20 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 ext_trim[17]
port 21 nsew signal input
rlabel metal2 s 5538 21540 5594 22340 6 ext_trim[18]
port 22 nsew signal input
rlabel metal3 s 19396 9528 20196 9648 6 ext_trim[19]
port 23 nsew signal input
rlabel metal2 s 11518 21540 11574 22340 6 ext_trim[1]
port 24 nsew signal input
rlabel metal2 s 9678 21540 9734 22340 6 ext_trim[20]
port 25 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 ext_trim[21]
port 26 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 ext_trim[22]
port 27 nsew signal input
rlabel metal3 s 19396 20408 20196 20528 6 ext_trim[23]
port 28 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 ext_trim[24]
port 29 nsew signal input
rlabel metal2 s 8298 21540 8354 22340 6 ext_trim[25]
port 30 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 ext_trim[2]
port 31 nsew signal input
rlabel metal3 s 19396 6808 20196 6928 6 ext_trim[3]
port 32 nsew signal input
rlabel metal3 s 19396 688 20196 808 6 ext_trim[4]
port 33 nsew signal input
rlabel metal3 s 19396 11568 20196 11688 6 ext_trim[5]
port 34 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 ext_trim[6]
port 35 nsew signal input
rlabel metal2 s 938 21540 994 22340 6 ext_trim[7]
port 36 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 ext_trim[8]
port 37 nsew signal input
rlabel metal3 s 19396 2728 20196 2848 6 ext_trim[9]
port 38 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 extclk_sel
port 39 nsew signal input
rlabel metal2 s 15658 21540 15714 22340 6 osc
port 40 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 reset
port 41 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 sel[0]
port 42 nsew signal input
rlabel metal2 s 18878 21540 18934 22340 6 sel[1]
port 43 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 sel[2]
port 44 nsew signal input
rlabel metal4 s 15894 2128 16214 20176 6 VPWR
port 45 nsew power bidirectional
rlabel metal4 s 9914 2128 10234 20176 6 VPWR
port 46 nsew power bidirectional
rlabel metal4 s 3934 2128 4254 20176 6 VPWR
port 47 nsew power bidirectional
rlabel metal5 s 1104 16928 19044 17248 6 VPWR
port 48 nsew power bidirectional
rlabel metal5 s 1104 10944 19044 11264 6 VPWR
port 49 nsew power bidirectional
rlabel metal5 s 1104 4960 19044 5280 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 12904 2128 13224 20176 6 VGND
port 51 nsew ground bidirectional
rlabel metal4 s 6924 2128 7244 20176 6 VGND
port 52 nsew ground bidirectional
rlabel metal5 s 1104 13936 19044 14256 6 VGND
port 53 nsew ground bidirectional
rlabel metal5 s 1104 7952 19044 8272 6 VGND
port 54 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20196 22340
<< end >>
