magic
tech sky130A
magscale 1 2
timestamp 1619516440
<< obsli1 >>
rect 1104 2159 17296 17969
<< obsm1 >>
rect 474 2128 17296 18080
<< metal2 >>
rect 478 19804 534 20604
rect 1858 19804 1914 20604
rect 3238 19804 3294 20604
rect 4618 19804 4674 20604
rect 5998 19804 6054 20604
rect 7378 19804 7434 20604
rect 8758 19804 8814 20604
rect 10138 19804 10194 20604
rect 11518 19804 11574 20604
rect 12898 19804 12954 20604
rect 14278 19804 14334 20604
rect 15658 19804 15714 20604
rect 17038 19804 17094 20604
rect 478 0 534 800
rect 1398 0 1454 800
rect 2778 0 2834 800
rect 4158 0 4214 800
rect 5538 0 5594 800
rect 6918 0 6974 800
rect 8298 0 8354 800
rect 9678 0 9734 800
rect 11058 0 11114 800
rect 12438 0 12494 800
rect 13818 0 13874 800
rect 15198 0 15254 800
rect 16578 0 16634 800
<< obsm2 >>
rect 590 19748 1802 19804
rect 1970 19748 3182 19804
rect 3350 19748 4562 19804
rect 4730 19748 5942 19804
rect 6110 19748 7322 19804
rect 7490 19748 8702 19804
rect 8870 19748 10082 19804
rect 10250 19748 11462 19804
rect 11630 19748 12842 19804
rect 13010 19748 14222 19804
rect 14390 19748 15602 19804
rect 15770 19748 16982 19804
rect 480 856 17094 19748
rect 590 711 1342 856
rect 1510 711 2722 856
rect 2890 711 4102 856
rect 4270 711 5482 856
rect 5650 711 6862 856
rect 7030 711 8242 856
rect 8410 711 9622 856
rect 9790 711 11002 856
rect 11170 711 12382 856
rect 12550 711 13762 856
rect 13930 711 15142 856
rect 15310 711 16522 856
rect 16690 711 17094 856
<< metal3 >>
rect 17660 19048 18460 19168
rect 0 18368 800 18488
rect 17660 17008 18460 17128
rect 0 16328 800 16448
rect 17660 14968 18460 15088
rect 0 14288 800 14408
rect 17660 12928 18460 13048
rect 0 12248 800 12368
rect 17660 10888 18460 11008
rect 0 10208 800 10328
rect 17660 8848 18460 8968
rect 0 8168 800 8288
rect 17660 6808 18460 6928
rect 0 6128 800 6248
rect 17660 4768 18460 4888
rect 0 4088 800 4208
rect 17660 2728 18460 2848
rect 0 2048 800 2168
rect 17660 688 18460 808
<< obsm3 >>
rect 800 18968 17580 19141
rect 800 18568 17660 18968
rect 880 18288 17660 18568
rect 800 17208 17660 18288
rect 800 16928 17580 17208
rect 800 16528 17660 16928
rect 880 16248 17660 16528
rect 800 15168 17660 16248
rect 800 14888 17580 15168
rect 800 14488 17660 14888
rect 880 14208 17660 14488
rect 800 13128 17660 14208
rect 800 12848 17580 13128
rect 800 12448 17660 12848
rect 880 12168 17660 12448
rect 800 11088 17660 12168
rect 800 10808 17580 11088
rect 800 10408 17660 10808
rect 880 10128 17660 10408
rect 800 9048 17660 10128
rect 800 8768 17580 9048
rect 800 8368 17660 8768
rect 880 8088 17660 8368
rect 800 7008 17660 8088
rect 800 6728 17580 7008
rect 800 6328 17660 6728
rect 880 6048 17660 6328
rect 800 4968 17660 6048
rect 800 4688 17580 4968
rect 800 4288 17660 4688
rect 880 4008 17660 4288
rect 800 2928 17660 4008
rect 800 2648 17580 2928
rect 800 2248 17660 2648
rect 880 1968 17660 2248
rect 800 888 17660 1968
rect 800 715 17580 888
<< metal4 >>
rect -916 156 -596 19972
rect -256 816 64 19312
rect 3643 156 3963 19972
rect 6341 156 6661 19972
rect 9040 156 9360 19972
rect 11739 156 12059 19972
rect 14437 156 14757 19972
rect 18336 816 18656 19312
rect 18996 156 19316 19972
<< obsm4 >>
rect 4043 156 6261 19972
rect 6741 156 8960 19972
rect 9440 156 11659 19972
<< metal5 >>
rect -916 19652 19316 19972
rect -256 18992 18656 19312
rect -916 15115 19316 15435
rect -916 12485 19316 12805
rect -916 9856 19316 10176
rect -916 7227 19316 7547
rect -916 4597 19316 4917
rect -256 816 18656 1136
rect -916 156 19316 476
<< obsm5 >>
rect -916 15114 19316 15115
rect 0 13125 18460 14795
rect 0 10496 18460 12165
rect 0 7867 18460 9536
rect -916 7226 19316 7227
<< labels >>
rlabel metal3 s 0 8168 800 8288 6 clockc
port 1 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 clockd[0]
port 2 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 clockd[1]
port 3 nsew signal output
rlabel metal3 s 17660 17008 18460 17128 6 clockd[2]
port 4 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 clockd[3]
port 5 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 clockp[0]
port 6 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 clockp[1]
port 7 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 dco
port 8 nsew signal input
rlabel metal3 s 17660 12928 18460 13048 6 div[0]
port 9 nsew signal input
rlabel metal2 s 15658 19804 15714 20604 6 div[1]
port 10 nsew signal input
rlabel metal2 s 5998 19804 6054 20604 6 div[2]
port 11 nsew signal input
rlabel metal2 s 478 0 534 800 6 div[3]
port 12 nsew signal input
rlabel metal2 s 11518 19804 11574 20604 6 div[4]
port 13 nsew signal input
rlabel metal2 s 12898 19804 12954 20604 6 ext_trim[0]
port 14 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 ext_trim[10]
port 15 nsew signal input
rlabel metal2 s 1858 19804 1914 20604 6 ext_trim[11]
port 16 nsew signal input
rlabel metal3 s 17660 4768 18460 4888 6 ext_trim[12]
port 17 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 ext_trim[13]
port 18 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 ext_trim[14]
port 19 nsew signal input
rlabel metal3 s 17660 14968 18460 15088 6 ext_trim[15]
port 20 nsew signal input
rlabel metal2 s 3238 19804 3294 20604 6 ext_trim[16]
port 21 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 ext_trim[17]
port 22 nsew signal input
rlabel metal2 s 4618 19804 4674 20604 6 ext_trim[18]
port 23 nsew signal input
rlabel metal3 s 17660 8848 18460 8968 6 ext_trim[19]
port 24 nsew signal input
rlabel metal2 s 10138 19804 10194 20604 6 ext_trim[1]
port 25 nsew signal input
rlabel metal2 s 8758 19804 8814 20604 6 ext_trim[20]
port 26 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 ext_trim[21]
port 27 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 ext_trim[22]
port 28 nsew signal input
rlabel metal3 s 17660 19048 18460 19168 6 ext_trim[23]
port 29 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 ext_trim[24]
port 30 nsew signal input
rlabel metal2 s 7378 19804 7434 20604 6 ext_trim[25]
port 31 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 ext_trim[2]
port 32 nsew signal input
rlabel metal3 s 17660 6808 18460 6928 6 ext_trim[3]
port 33 nsew signal input
rlabel metal3 s 17660 688 18460 808 6 ext_trim[4]
port 34 nsew signal input
rlabel metal3 s 17660 10888 18460 11008 6 ext_trim[5]
port 35 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 ext_trim[6]
port 36 nsew signal input
rlabel metal2 s 478 19804 534 20604 6 ext_trim[7]
port 37 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 ext_trim[8]
port 38 nsew signal input
rlabel metal3 s 17660 2728 18460 2848 6 ext_trim[9]
port 39 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 extclk_sel
port 40 nsew signal input
rlabel metal2 s 14278 19804 14334 20604 6 osc
port 41 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 reset
port 42 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 sel[0]
port 43 nsew signal input
rlabel metal2 s 17038 19804 17094 20604 6 sel[1]
port 44 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 sel[2]
port 45 nsew signal input
rlabel metal4 s 14437 156 14757 19972 6 VPWR
port 46 nsew power bidirectional
rlabel metal4 s 9040 156 9360 19972 6 VPWR
port 47 nsew power bidirectional
rlabel metal4 s 3643 156 3963 19972 6 VPWR
port 48 nsew power bidirectional
rlabel metal4 s 18336 816 18656 19312 6 VPWR
port 49 nsew power bidirectional
rlabel metal4 s -256 816 64 19312 4 VPWR
port 50 nsew power bidirectional
rlabel metal5 s -256 18992 18656 19312 6 VPWR
port 51 nsew power bidirectional
rlabel metal5 s -916 15115 19316 15435 6 VPWR
port 52 nsew power bidirectional
rlabel metal5 s -916 9856 19316 10176 6 VPWR
port 53 nsew power bidirectional
rlabel metal5 s -916 4597 19316 4917 6 VPWR
port 54 nsew power bidirectional
rlabel metal5 s -256 816 18656 1136 6 VPWR
port 55 nsew power bidirectional
rlabel metal4 s 18996 156 19316 19972 6 VGND
port 56 nsew ground bidirectional
rlabel metal4 s 11739 156 12059 19972 6 VGND
port 57 nsew ground bidirectional
rlabel metal4 s 6341 156 6661 19972 6 VGND
port 58 nsew ground bidirectional
rlabel metal4 s -916 156 -596 19972 4 VGND
port 59 nsew ground bidirectional
rlabel metal5 s -916 19652 19316 19972 6 VGND
port 60 nsew ground bidirectional
rlabel metal5 s -916 12485 19316 12805 6 VGND
port 61 nsew ground bidirectional
rlabel metal5 s -916 7227 19316 7547 6 VGND
port 62 nsew ground bidirectional
rlabel metal5 s -916 156 19316 476 6 VGND
port 63 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 18460 20604
string LEFview TRUE
string GDS_FILE /openLANE_flow/designs/digital_pll/runs/fifth_run/results/magic/digital_pll.gds
string GDS_END 1425158
string GDS_START 514058
<< end >>

