magic
tech sky130A
magscale 1 2
timestamp 1619632572
<< locali >>
rect 8401 16031 8435 16201
rect 9873 15555 9907 15657
rect 7113 13923 7147 14025
rect 19441 13379 19475 13481
rect 17141 11067 17175 11169
rect 21925 5899 21959 6681
<< viali >>
rect 1501 22729 1535 22763
rect 2973 22661 3007 22695
rect 8033 22661 8067 22695
rect 1777 22525 1811 22559
rect 2789 22525 2823 22559
rect 4629 22525 4663 22559
rect 6009 22525 6043 22559
rect 7849 22525 7883 22559
rect 9689 22525 9723 22559
rect 11713 22525 11747 22559
rect 12909 22525 12943 22559
rect 14933 22525 14967 22559
rect 16773 22525 16807 22559
rect 18153 22525 18187 22559
rect 20085 22525 20119 22559
rect 21097 22525 21131 22559
rect 21465 22525 21499 22559
rect 1593 22457 1627 22491
rect 1961 22389 1995 22423
rect 4813 22389 4847 22423
rect 6193 22389 6227 22423
rect 9873 22389 9907 22423
rect 11529 22389 11563 22423
rect 13093 22389 13127 22423
rect 14749 22389 14783 22423
rect 16589 22389 16623 22423
rect 17969 22389 18003 22423
rect 19901 22389 19935 22423
rect 20913 22389 20947 22423
rect 21281 22389 21315 22423
rect 4997 22049 5031 22083
rect 5089 22049 5123 22083
rect 5365 22049 5399 22083
rect 5641 22049 5675 22083
rect 7573 22049 7607 22083
rect 9873 22049 9907 22083
rect 11713 22049 11747 22083
rect 11897 22049 11931 22083
rect 11989 22049 12023 22083
rect 12127 22049 12161 22083
rect 12725 22049 12759 22083
rect 15209 22049 15243 22083
rect 18337 22049 18371 22083
rect 19993 22049 20027 22083
rect 4813 21845 4847 21879
rect 5273 21845 5307 21879
rect 5457 21845 5491 21879
rect 7757 21845 7791 21879
rect 10057 21845 10091 21879
rect 12265 21845 12299 21879
rect 12909 21845 12943 21879
rect 15393 21845 15427 21879
rect 18521 21845 18555 21879
rect 20177 21845 20211 21879
rect 1777 21641 1811 21675
rect 5641 21641 5675 21675
rect 5825 21641 5859 21675
rect 4169 21505 4203 21539
rect 9045 21505 9079 21539
rect 9321 21505 9355 21539
rect 10885 21505 10919 21539
rect 12081 21505 12115 21539
rect 14289 21505 14323 21539
rect 16037 21505 16071 21539
rect 17417 21505 17451 21539
rect 19165 21505 19199 21539
rect 19533 21505 19567 21539
rect 1961 21437 1995 21471
rect 3893 21437 3927 21471
rect 5733 21437 5767 21471
rect 6653 21437 6687 21471
rect 11805 21437 11839 21471
rect 17141 21437 17175 21471
rect 19257 21437 19291 21471
rect 6929 21369 6963 21403
rect 11069 21369 11103 21403
rect 11253 21369 11287 21403
rect 14565 21369 14599 21403
rect 17693 21369 17727 21403
rect 8401 21301 8435 21335
rect 10793 21301 10827 21335
rect 13553 21301 13587 21335
rect 17325 21301 17359 21335
rect 21005 21301 21039 21335
rect 7205 21097 7239 21131
rect 14657 21097 14691 21131
rect 7481 21029 7515 21063
rect 7573 21029 7607 21063
rect 7711 21029 7745 21063
rect 12081 21029 12115 21063
rect 14933 21029 14967 21063
rect 7389 20961 7423 20995
rect 7849 20961 7883 20995
rect 8217 20961 8251 20995
rect 11989 20961 12023 20995
rect 12173 20961 12207 20995
rect 12357 20961 12391 20995
rect 14841 20961 14875 20995
rect 15025 20961 15059 20995
rect 15209 20961 15243 20995
rect 16221 20961 16255 20995
rect 21281 20961 21315 20995
rect 16497 20893 16531 20927
rect 8309 20757 8343 20791
rect 11805 20757 11839 20791
rect 17969 20757 18003 20791
rect 21373 20757 21407 20791
rect 9597 20417 9631 20451
rect 9873 20417 9907 20451
rect 11345 20417 11379 20451
rect 1409 20349 1443 20383
rect 2513 20349 2547 20383
rect 5273 20349 5307 20383
rect 5457 20349 5491 20383
rect 11897 20349 11931 20383
rect 12081 20349 12115 20383
rect 12357 20349 12391 20383
rect 12541 20349 12575 20383
rect 12633 20349 12667 20383
rect 15117 20349 15151 20383
rect 20729 20349 20763 20383
rect 20821 20349 20855 20383
rect 21189 20349 21223 20383
rect 21281 20349 21315 20383
rect 2789 20281 2823 20315
rect 20177 20281 20211 20315
rect 1593 20213 1627 20247
rect 4261 20213 4295 20247
rect 5365 20213 5399 20247
rect 15025 20213 15059 20247
rect 3525 20009 3559 20043
rect 4721 20009 4755 20043
rect 7757 20009 7791 20043
rect 8217 20009 8251 20043
rect 10517 20009 10551 20043
rect 21373 20009 21407 20043
rect 5825 19941 5859 19975
rect 7941 19941 7975 19975
rect 15301 19941 15335 19975
rect 15393 19941 15427 19975
rect 3709 19873 3743 19907
rect 4905 19873 4939 19907
rect 4997 19873 5031 19907
rect 5089 19873 5123 19907
rect 5207 19873 5241 19907
rect 5457 19873 5491 19907
rect 5641 19873 5675 19907
rect 5917 19873 5951 19907
rect 8125 19873 8159 19907
rect 8217 19873 8251 19907
rect 8401 19873 8435 19907
rect 10333 19873 10367 19907
rect 15117 19873 15151 19907
rect 15485 19873 15519 19907
rect 15761 19873 15795 19907
rect 16129 19873 16163 19907
rect 16221 19873 16255 19907
rect 16405 19873 16439 19907
rect 19625 19873 19659 19907
rect 5365 19805 5399 19839
rect 14565 19805 14599 19839
rect 14657 19805 14691 19839
rect 15025 19805 15059 19839
rect 19901 19805 19935 19839
rect 16405 19737 16439 19771
rect 6009 19669 6043 19703
rect 14381 19669 14415 19703
rect 15669 19669 15703 19703
rect 15853 19669 15887 19703
rect 5181 19465 5215 19499
rect 5641 19465 5675 19499
rect 7941 19465 7975 19499
rect 20637 19465 20671 19499
rect 6009 19397 6043 19431
rect 5825 19329 5859 19363
rect 8033 19329 8067 19363
rect 8217 19329 8251 19363
rect 14657 19329 14691 19363
rect 5365 19261 5399 19295
rect 5457 19261 5491 19295
rect 5733 19261 5767 19295
rect 6101 19261 6135 19295
rect 7389 19261 7423 19295
rect 7573 19261 7607 19295
rect 7757 19261 7791 19295
rect 8309 19261 8343 19295
rect 8585 19261 8619 19295
rect 12725 19261 12759 19295
rect 13829 19261 13863 19295
rect 14013 19261 14047 19295
rect 14381 19261 14415 19295
rect 14565 19261 14599 19295
rect 14749 19261 14783 19295
rect 14933 19261 14967 19295
rect 15393 19261 15427 19295
rect 17601 19261 17635 19295
rect 20453 19261 20487 19295
rect 7665 19193 7699 19227
rect 8033 19193 8067 19227
rect 14197 19193 14231 19227
rect 15025 19193 15059 19227
rect 15209 19193 15243 19227
rect 5825 19125 5859 19159
rect 8677 19125 8711 19159
rect 12633 19125 12667 19159
rect 13829 19125 13863 19159
rect 17785 19125 17819 19159
rect 19073 18921 19107 18955
rect 8769 18853 8803 18887
rect 9505 18853 9539 18887
rect 13001 18853 13035 18887
rect 16589 18853 16623 18887
rect 16957 18853 16991 18887
rect 6561 18785 6595 18819
rect 8677 18785 8711 18819
rect 9137 18785 9171 18819
rect 9230 18785 9264 18819
rect 9413 18785 9447 18819
rect 9602 18785 9636 18819
rect 12541 18785 12575 18819
rect 12633 18785 12667 18819
rect 12909 18785 12943 18819
rect 13369 18785 13403 18819
rect 15853 18785 15887 18819
rect 16037 18785 16071 18819
rect 16129 18785 16163 18819
rect 16405 18785 16439 18819
rect 19165 18785 19199 18819
rect 19257 18785 19291 18819
rect 19625 18785 19659 18819
rect 19809 18785 19843 18819
rect 12817 18717 12851 18751
rect 13093 18717 13127 18751
rect 16221 18717 16255 18751
rect 16681 18717 16715 18751
rect 18429 18717 18463 18751
rect 18797 18717 18831 18751
rect 12357 18649 12391 18683
rect 6653 18581 6687 18615
rect 9781 18581 9815 18615
rect 13185 18581 13219 18615
rect 13277 18581 13311 18615
rect 19717 18581 19751 18615
rect 8493 18377 8527 18411
rect 8953 18377 8987 18411
rect 16681 18377 16715 18411
rect 18705 18309 18739 18343
rect 2697 18241 2731 18275
rect 2973 18241 3007 18275
rect 9413 18241 9447 18275
rect 19533 18241 19567 18275
rect 8677 18173 8711 18207
rect 8799 18173 8833 18207
rect 9045 18173 9079 18207
rect 9137 18173 9171 18207
rect 9229 18173 9263 18207
rect 10333 18173 10367 18207
rect 12633 18173 12667 18207
rect 12817 18173 12851 18207
rect 13001 18173 13035 18207
rect 13277 18173 13311 18207
rect 13461 18173 13495 18207
rect 16589 18173 16623 18207
rect 16773 18173 16807 18207
rect 18797 18173 18831 18207
rect 19257 18173 19291 18207
rect 19441 18173 19475 18207
rect 19625 18173 19659 18207
rect 19809 18173 19843 18207
rect 12173 18105 12207 18139
rect 4445 18037 4479 18071
rect 9413 18037 9447 18071
rect 10517 18037 10551 18071
rect 19073 18037 19107 18071
rect 3893 17833 3927 17867
rect 4629 17833 4663 17867
rect 6009 17833 6043 17867
rect 4905 17765 4939 17799
rect 4997 17765 5031 17799
rect 5549 17765 5583 17799
rect 9597 17765 9631 17799
rect 14841 17765 14875 17799
rect 1409 17697 1443 17731
rect 4077 17697 4111 17731
rect 4813 17697 4847 17731
rect 5135 17697 5169 17731
rect 5273 17697 5307 17731
rect 5733 17697 5767 17731
rect 6193 17697 6227 17731
rect 6377 17697 6411 17731
rect 6469 17697 6503 17731
rect 8033 17697 8067 17731
rect 8493 17697 8527 17731
rect 9321 17697 9355 17731
rect 12173 17697 12207 17731
rect 12541 17697 12575 17731
rect 14749 17697 14783 17731
rect 14933 17697 14967 17731
rect 15117 17697 15151 17731
rect 20729 17697 20763 17731
rect 21465 17697 21499 17731
rect 6561 17629 6595 17663
rect 8217 17629 8251 17663
rect 8309 17629 8343 17663
rect 8125 17561 8159 17595
rect 12265 17561 12299 17595
rect 1593 17493 1627 17527
rect 5365 17493 5399 17527
rect 7849 17493 7883 17527
rect 11069 17493 11103 17527
rect 12633 17493 12667 17527
rect 14565 17493 14599 17527
rect 20913 17493 20947 17527
rect 21281 17493 21315 17527
rect 7113 17289 7147 17323
rect 10241 17289 10275 17323
rect 13001 17289 13035 17323
rect 13369 17289 13403 17323
rect 16221 17289 16255 17323
rect 5825 17221 5859 17255
rect 11989 17221 12023 17255
rect 6745 17153 6779 17187
rect 12449 17153 12483 17187
rect 12633 17153 12667 17187
rect 13093 17153 13127 17187
rect 14473 17153 14507 17187
rect 14749 17153 14783 17187
rect 19717 17153 19751 17187
rect 5549 17085 5583 17119
rect 5641 17085 5675 17119
rect 5917 17085 5951 17119
rect 6009 17085 6043 17119
rect 6469 17085 6503 17119
rect 6653 17085 6687 17119
rect 6837 17085 6871 17119
rect 6929 17085 6963 17119
rect 10149 17085 10183 17119
rect 11897 17085 11931 17119
rect 12357 17085 12391 17119
rect 12725 17085 12759 17119
rect 13001 17085 13035 17119
rect 5365 17017 5399 17051
rect 6101 17017 6135 17051
rect 19993 17017 20027 17051
rect 21465 16949 21499 16983
rect 17785 16745 17819 16779
rect 20177 16745 20211 16779
rect 6101 16677 6135 16711
rect 17141 16677 17175 16711
rect 17233 16677 17267 16711
rect 19809 16677 19843 16711
rect 19901 16677 19935 16711
rect 5825 16609 5859 16643
rect 6285 16609 6319 16643
rect 8125 16609 8159 16643
rect 8217 16609 8251 16643
rect 17049 16609 17083 16643
rect 17417 16609 17451 16643
rect 17509 16609 17543 16643
rect 17601 16609 17635 16643
rect 19625 16609 19659 16643
rect 19993 16609 20027 16643
rect 20453 16609 20487 16643
rect 6101 16541 6135 16575
rect 5917 16473 5951 16507
rect 6377 16405 6411 16439
rect 16865 16405 16899 16439
rect 20361 16405 20395 16439
rect 8401 16201 8435 16235
rect 14473 16201 14507 16235
rect 18705 16201 18739 16235
rect 19073 16201 19107 16235
rect 15025 16133 15059 16167
rect 16957 16065 16991 16099
rect 17233 16065 17267 16099
rect 1593 15997 1627 16031
rect 2145 15997 2179 16031
rect 6469 15997 6503 16031
rect 6562 15997 6596 16031
rect 6745 15997 6779 16031
rect 6934 15997 6968 16031
rect 7205 15997 7239 16031
rect 8309 15997 8343 16031
rect 8401 15997 8435 16031
rect 8493 15997 8527 16031
rect 8586 15997 8620 16031
rect 8861 15997 8895 16031
rect 8958 15997 8992 16031
rect 10977 15997 11011 16031
rect 14654 15997 14688 16031
rect 15117 15997 15151 16031
rect 15393 15997 15427 16031
rect 15669 15997 15703 16031
rect 15761 15997 15795 16031
rect 15945 15997 15979 16031
rect 19257 15997 19291 16031
rect 19533 15997 19567 16031
rect 19717 15997 19751 16031
rect 19901 15997 19935 16031
rect 2053 15929 2087 15963
rect 6837 15929 6871 15963
rect 7297 15929 7331 15963
rect 8217 15929 8251 15963
rect 8769 15929 8803 15963
rect 15853 15929 15887 15963
rect 19441 15929 19475 15963
rect 19993 15929 20027 15963
rect 7113 15861 7147 15895
rect 9137 15861 9171 15895
rect 11161 15861 11195 15895
rect 14657 15861 14691 15895
rect 15209 15861 15243 15895
rect 15577 15861 15611 15895
rect 8861 15657 8895 15691
rect 9873 15657 9907 15691
rect 12173 15657 12207 15691
rect 12817 15657 12851 15691
rect 12909 15657 12943 15691
rect 14381 15657 14415 15691
rect 14565 15657 14599 15691
rect 17141 15657 17175 15691
rect 17325 15657 17359 15691
rect 19901 15657 19935 15691
rect 20085 15657 20119 15691
rect 21281 15657 21315 15691
rect 9137 15589 9171 15623
rect 10241 15589 10275 15623
rect 13277 15589 13311 15623
rect 16957 15589 16991 15623
rect 17233 15589 17267 15623
rect 1409 15521 1443 15555
rect 2605 15521 2639 15555
rect 3065 15521 3099 15555
rect 3249 15521 3283 15555
rect 8309 15521 8343 15555
rect 8585 15521 8619 15555
rect 8677 15521 8711 15555
rect 9413 15521 9447 15555
rect 9873 15521 9907 15555
rect 9965 15521 9999 15555
rect 12357 15521 12391 15555
rect 13093 15521 13127 15555
rect 14562 15521 14596 15555
rect 14933 15521 14967 15555
rect 19625 15521 19659 15555
rect 19809 15521 19843 15555
rect 20177 15521 20211 15555
rect 21465 15521 21499 15555
rect 2053 15453 2087 15487
rect 9137 15453 9171 15487
rect 9321 15453 9355 15487
rect 12449 15453 12483 15487
rect 15025 15453 15059 15487
rect 2513 15385 2547 15419
rect 1593 15317 1627 15351
rect 8401 15317 8435 15351
rect 11713 15317 11747 15351
rect 17509 15317 17543 15351
rect 1593 15113 1627 15147
rect 6653 15113 6687 15147
rect 6837 15113 6871 15147
rect 7297 15113 7331 15147
rect 13093 15113 13127 15147
rect 3893 15045 3927 15079
rect 3985 15045 4019 15079
rect 9505 15045 9539 15079
rect 10333 15045 10367 15079
rect 14289 15045 14323 15079
rect 2053 14977 2087 15011
rect 2145 14977 2179 15011
rect 3525 14977 3559 15011
rect 6469 14977 6503 15011
rect 10057 14977 10091 15011
rect 13645 14977 13679 15011
rect 13737 14977 13771 15011
rect 2881 14909 2915 14943
rect 3433 14909 3467 14943
rect 4169 14909 4203 14943
rect 5089 14909 5123 14943
rect 6745 14909 6779 14943
rect 7021 14909 7055 14943
rect 7113 14909 7147 14943
rect 7389 14909 7423 14943
rect 10241 14909 10275 14943
rect 13277 14909 13311 14943
rect 13369 14909 13403 14943
rect 14565 14909 14599 14943
rect 19809 14909 19843 14943
rect 19993 14909 20027 14943
rect 20177 14909 20211 14943
rect 2973 14841 3007 14875
rect 9781 14841 9815 14875
rect 14289 14841 14323 14875
rect 19901 14841 19935 14875
rect 1961 14773 1995 14807
rect 3893 14773 3927 14807
rect 4905 14773 4939 14807
rect 6469 14773 6503 14807
rect 9965 14773 9999 14807
rect 14473 14773 14507 14807
rect 19625 14773 19659 14807
rect 14565 14569 14599 14603
rect 14749 14569 14783 14603
rect 17325 14569 17359 14603
rect 18981 14569 19015 14603
rect 20177 14569 20211 14603
rect 20361 14569 20395 14603
rect 5641 14501 5675 14535
rect 15393 14501 15427 14535
rect 5917 14433 5951 14467
rect 12817 14433 12851 14467
rect 14746 14433 14780 14467
rect 15209 14433 15243 14467
rect 15301 14433 15335 14467
rect 15485 14433 15519 14467
rect 15761 14433 15795 14467
rect 17417 14433 17451 14467
rect 18889 14433 18923 14467
rect 20302 14433 20336 14467
rect 20821 14433 20855 14467
rect 12909 14365 12943 14399
rect 15117 14297 15151 14331
rect 15669 14297 15703 14331
rect 4169 14229 4203 14263
rect 20729 14229 20763 14263
rect 6469 14025 6503 14059
rect 7113 14025 7147 14059
rect 8125 14025 8159 14059
rect 10241 14025 10275 14059
rect 17877 14025 17911 14059
rect 18153 14025 18187 14059
rect 6193 13957 6227 13991
rect 7849 13957 7883 13991
rect 9873 13957 9907 13991
rect 17509 13957 17543 13991
rect 6745 13889 6779 13923
rect 7113 13889 7147 13923
rect 9781 13889 9815 13923
rect 17969 13889 18003 13923
rect 6101 13821 6135 13855
rect 6653 13821 6687 13855
rect 6837 13821 6871 13855
rect 6929 13821 6963 13855
rect 7297 13821 7331 13855
rect 7481 13821 7515 13855
rect 7757 13821 7791 13855
rect 8033 13821 8067 13855
rect 9505 13821 9539 13855
rect 9689 13821 9723 13855
rect 9965 13821 9999 13855
rect 17785 13821 17819 13855
rect 17877 13821 17911 13855
rect 18245 13821 18279 13855
rect 18797 13821 18831 13855
rect 18889 13753 18923 13787
rect 7665 13685 7699 13719
rect 17969 13685 18003 13719
rect 1869 13481 1903 13515
rect 3341 13481 3375 13515
rect 7389 13481 7423 13515
rect 8309 13481 8343 13515
rect 17785 13481 17819 13515
rect 19441 13481 19475 13515
rect 12081 13413 12115 13447
rect 12173 13413 12207 13447
rect 14657 13413 14691 13447
rect 17417 13413 17451 13447
rect 19901 13413 19935 13447
rect 1961 13345 1995 13379
rect 3249 13345 3283 13379
rect 7297 13345 7331 13379
rect 8217 13345 8251 13379
rect 12817 13345 12851 13379
rect 13001 13345 13035 13379
rect 14565 13345 14599 13379
rect 14749 13345 14783 13379
rect 14933 13345 14967 13379
rect 18061 13345 18095 13379
rect 18153 13345 18187 13379
rect 18705 13345 18739 13379
rect 18889 13345 18923 13379
rect 19073 13345 19107 13379
rect 19257 13345 19291 13379
rect 19441 13345 19475 13379
rect 19625 13345 19659 13379
rect 19809 13345 19843 13379
rect 19993 13345 20027 13379
rect 20637 13345 20671 13379
rect 21465 13345 21499 13379
rect 1777 13277 1811 13311
rect 12173 13277 12207 13311
rect 15669 13277 15703 13311
rect 17693 13277 17727 13311
rect 17969 13277 18003 13311
rect 18245 13277 18279 13311
rect 18981 13277 19015 13311
rect 12633 13209 12667 13243
rect 21281 13209 21315 13243
rect 2329 13141 2363 13175
rect 13185 13141 13219 13175
rect 14381 13141 14415 13175
rect 18521 13141 18555 13175
rect 20177 13141 20211 13175
rect 20821 13141 20855 13175
rect 1501 12937 1535 12971
rect 2697 12937 2731 12971
rect 3157 12937 3191 12971
rect 4905 12937 4939 12971
rect 5273 12937 5307 12971
rect 6745 12937 6779 12971
rect 9229 12937 9263 12971
rect 9873 12937 9907 12971
rect 10057 12937 10091 12971
rect 16589 12937 16623 12971
rect 17417 12937 17451 12971
rect 21465 12937 21499 12971
rect 9965 12869 9999 12903
rect 11437 12869 11471 12903
rect 2789 12801 2823 12835
rect 8125 12801 8159 12835
rect 9321 12801 9355 12835
rect 10425 12801 10459 12835
rect 12173 12801 12207 12835
rect 12265 12801 12299 12835
rect 13461 12801 13495 12835
rect 19717 12801 19751 12835
rect 19993 12801 20027 12835
rect 2145 12733 2179 12767
rect 2697 12733 2731 12767
rect 3157 12733 3191 12767
rect 5181 12733 5215 12767
rect 5273 12733 5307 12767
rect 6469 12733 6503 12767
rect 7757 12733 7791 12767
rect 8309 12733 8343 12767
rect 8493 12733 8527 12767
rect 9229 12733 9263 12767
rect 9689 12733 9723 12767
rect 10149 12733 10183 12767
rect 10793 12733 10827 12767
rect 10977 12733 11011 12767
rect 13277 12733 13311 12767
rect 13369 12733 13403 12767
rect 14749 12733 14783 12767
rect 16773 12733 16807 12767
rect 17325 12733 17359 12767
rect 18889 12733 18923 12767
rect 1593 12665 1627 12699
rect 6653 12665 6687 12699
rect 7573 12665 7607 12699
rect 11069 12665 11103 12699
rect 11253 12665 11287 12699
rect 19073 12665 19107 12699
rect 8493 12597 8527 12631
rect 9597 12597 9631 12631
rect 10885 12597 10919 12631
rect 11713 12597 11747 12631
rect 12081 12597 12115 12631
rect 12909 12597 12943 12631
rect 14933 12597 14967 12631
rect 19257 12597 19291 12631
rect 5549 12393 5583 12427
rect 11989 12393 12023 12427
rect 14381 12393 14415 12427
rect 3341 12325 3375 12359
rect 15853 12325 15887 12359
rect 3525 12257 3559 12291
rect 5641 12257 5675 12291
rect 6009 12257 6043 12291
rect 6285 12257 6319 12291
rect 11713 12257 11747 12291
rect 11805 12257 11839 12291
rect 16129 12257 16163 12291
rect 5549 12189 5583 12223
rect 6101 12189 6135 12223
rect 6193 12189 6227 12223
rect 5825 12121 5859 12155
rect 5089 12053 5123 12087
rect 9413 11781 9447 11815
rect 5641 11713 5675 11747
rect 5825 11713 5859 11747
rect 5917 11713 5951 11747
rect 6469 11713 6503 11747
rect 8033 11713 8067 11747
rect 8217 11713 8251 11747
rect 10149 11713 10183 11747
rect 5733 11645 5767 11679
rect 6837 11645 6871 11679
rect 7941 11645 7975 11679
rect 8125 11645 8159 11679
rect 9321 11645 9355 11679
rect 9597 11645 9631 11679
rect 10241 11645 10275 11679
rect 10425 11645 10459 11679
rect 6653 11577 6687 11611
rect 10057 11577 10091 11611
rect 5457 11509 5491 11543
rect 8401 11509 8435 11543
rect 10609 11509 10643 11543
rect 1869 11305 1903 11339
rect 4261 11305 4295 11339
rect 10425 11305 10459 11339
rect 11805 11305 11839 11339
rect 18429 11305 18463 11339
rect 3065 11237 3099 11271
rect 7021 11237 7055 11271
rect 8125 11237 8159 11271
rect 10057 11237 10091 11271
rect 10262 11237 10296 11271
rect 11897 11237 11931 11271
rect 12909 11237 12943 11271
rect 1961 11169 1995 11203
rect 2973 11169 3007 11203
rect 3525 11169 3559 11203
rect 4537 11169 4571 11203
rect 6929 11169 6963 11203
rect 7205 11169 7239 11203
rect 7297 11169 7331 11203
rect 7573 11169 7607 11203
rect 7757 11169 7791 11203
rect 8401 11169 8435 11203
rect 8493 11169 8527 11203
rect 13001 11169 13035 11203
rect 15025 11169 15059 11203
rect 17141 11169 17175 11203
rect 17233 11169 17267 11203
rect 17785 11169 17819 11203
rect 20085 11169 20119 11203
rect 1777 11101 1811 11135
rect 3893 11101 3927 11135
rect 7481 11101 7515 11135
rect 8217 11101 8251 11135
rect 11805 11101 11839 11135
rect 12725 11101 12759 11135
rect 18153 11101 18187 11135
rect 18337 11101 18371 11135
rect 2329 11033 2363 11067
rect 4261 11033 4295 11067
rect 4353 11033 4387 11067
rect 7389 11033 7423 11067
rect 7757 11033 7791 11067
rect 11345 11033 11379 11067
rect 13369 11033 13403 11067
rect 15209 11033 15243 11067
rect 17141 11033 17175 11067
rect 18797 11033 18831 11067
rect 20269 11033 20303 11067
rect 8309 10965 8343 10999
rect 10241 10965 10275 10999
rect 17233 10965 17267 10999
rect 4629 10761 4663 10795
rect 4997 10761 5031 10795
rect 7941 10761 7975 10795
rect 13461 10761 13495 10795
rect 15393 10761 15427 10795
rect 16129 10761 16163 10795
rect 17233 10761 17267 10795
rect 17693 10761 17727 10795
rect 18521 10761 18555 10795
rect 20913 10761 20947 10795
rect 6745 10625 6779 10659
rect 6929 10625 6963 10659
rect 9321 10625 9355 10659
rect 13093 10625 13127 10659
rect 15761 10625 15795 10659
rect 17601 10625 17635 10659
rect 18245 10625 18279 10659
rect 19165 10625 19199 10659
rect 19441 10625 19475 10659
rect 2697 10557 2731 10591
rect 4813 10557 4847 10591
rect 5089 10557 5123 10591
rect 6653 10557 6687 10591
rect 6837 10557 6871 10591
rect 8033 10557 8067 10591
rect 9137 10557 9171 10591
rect 9413 10557 9447 10591
rect 9505 10557 9539 10591
rect 13461 10557 13495 10591
rect 14841 10557 14875 10591
rect 15393 10557 15427 10591
rect 16129 10557 16163 10591
rect 16957 10557 16991 10591
rect 17141 10557 17175 10591
rect 17233 10557 17267 10591
rect 18705 10557 18739 10591
rect 2881 10489 2915 10523
rect 18061 10489 18095 10523
rect 6469 10421 6503 10455
rect 8953 10421 8987 10455
rect 9597 10421 9631 10455
rect 18153 10421 18187 10455
rect 1501 10217 1535 10251
rect 5273 10217 5307 10251
rect 6377 10217 6411 10251
rect 13645 10217 13679 10251
rect 21281 10217 21315 10251
rect 5457 10149 5491 10183
rect 6285 10149 6319 10183
rect 13369 10149 13403 10183
rect 1593 10081 1627 10115
rect 9781 10081 9815 10115
rect 10057 10081 10091 10115
rect 10241 10081 10275 10115
rect 12909 10081 12943 10115
rect 13461 10081 13495 10115
rect 13553 10081 13587 10115
rect 21465 10081 21499 10115
rect 5181 10013 5215 10047
rect 6469 10013 6503 10047
rect 9229 10013 9263 10047
rect 9965 10013 9999 10047
rect 5733 9945 5767 9979
rect 5917 9877 5951 9911
rect 10425 9877 10459 9911
rect 2789 9605 2823 9639
rect 2881 9605 2915 9639
rect 5273 9605 5307 9639
rect 12725 9605 12759 9639
rect 12817 9605 12851 9639
rect 2421 9537 2455 9571
rect 7389 9537 7423 9571
rect 9505 9537 9539 9571
rect 9689 9537 9723 9571
rect 10609 9537 10643 9571
rect 10701 9537 10735 9571
rect 12357 9537 12391 9571
rect 1777 9469 1811 9503
rect 2329 9469 2363 9503
rect 3065 9469 3099 9503
rect 4997 9469 5031 9503
rect 8033 9469 8067 9503
rect 8309 9469 8343 9503
rect 10425 9469 10459 9503
rect 11713 9469 11747 9503
rect 12265 9469 12299 9503
rect 13001 9469 13035 9503
rect 2237 9401 2271 9435
rect 4721 9401 4755 9435
rect 9781 9401 9815 9435
rect 10241 9401 10275 9435
rect 12173 9401 12207 9435
rect 2743 9333 2777 9367
rect 4813 9333 4847 9367
rect 10149 9333 10183 9367
rect 12725 9333 12759 9367
rect 2697 9129 2731 9163
rect 4905 9129 4939 9163
rect 14565 9129 14599 9163
rect 15209 9129 15243 9163
rect 15301 9129 15335 9163
rect 11713 9061 11747 9095
rect 16773 9061 16807 9095
rect 4721 8993 4755 9027
rect 4997 8993 5031 9027
rect 6653 8993 6687 9027
rect 6837 8993 6871 9027
rect 9505 8993 9539 9027
rect 9689 8993 9723 9027
rect 11529 8993 11563 9027
rect 14381 8993 14415 9027
rect 18429 8993 18463 9027
rect 7205 8925 7239 8959
rect 15393 8925 15427 8959
rect 2789 8789 2823 8823
rect 4537 8789 4571 8823
rect 9597 8789 9631 8823
rect 9873 8789 9907 8823
rect 14841 8789 14875 8823
rect 16865 8789 16899 8823
rect 18337 8789 18371 8823
rect 2145 8585 2179 8619
rect 16773 8585 16807 8619
rect 17325 8585 17359 8619
rect 1593 8517 1627 8551
rect 7113 8517 7147 8551
rect 19165 8517 19199 8551
rect 19257 8517 19291 8551
rect 2605 8449 2639 8483
rect 2697 8449 2731 8483
rect 2973 8449 3007 8483
rect 3525 8449 3559 8483
rect 6653 8449 6687 8483
rect 8309 8449 8343 8483
rect 16957 8449 16991 8483
rect 17325 8449 17359 8483
rect 18797 8449 18831 8483
rect 1409 8381 1443 8415
rect 2513 8381 2547 8415
rect 6561 8381 6595 8415
rect 7573 8381 7607 8415
rect 8493 8381 8527 8415
rect 8585 8381 8619 8415
rect 11897 8381 11931 8415
rect 12081 8381 12115 8415
rect 16221 8381 16255 8415
rect 16773 8381 16807 8415
rect 18153 8381 18187 8415
rect 18705 8381 18739 8415
rect 19441 8381 19475 8415
rect 21465 8381 21499 8415
rect 3433 8313 3467 8347
rect 6653 8313 6687 8347
rect 12265 8313 12299 8347
rect 18245 8313 18279 8347
rect 19165 8245 19199 8279
rect 21281 8245 21315 8279
rect 12817 8041 12851 8075
rect 15393 8041 15427 8075
rect 8033 7973 8067 8007
rect 8401 7973 8435 8007
rect 12909 7973 12943 8007
rect 16405 7973 16439 8007
rect 2145 7905 2179 7939
rect 2697 7905 2731 7939
rect 7665 7905 7699 7939
rect 8585 7905 8619 7939
rect 9873 7905 9907 7939
rect 14381 7905 14415 7939
rect 14473 7905 14507 7939
rect 14933 7905 14967 7939
rect 15025 7905 15059 7939
rect 15669 7905 15703 7939
rect 16221 7905 16255 7939
rect 13001 7837 13035 7871
rect 15393 7769 15427 7803
rect 15485 7769 15519 7803
rect 2697 7701 2731 7735
rect 8309 7701 8343 7735
rect 9781 7701 9815 7735
rect 12449 7701 12483 7735
rect 7665 7497 7699 7531
rect 12817 7497 12851 7531
rect 13277 7497 13311 7531
rect 3709 7429 3743 7463
rect 8585 7361 8619 7395
rect 12909 7361 12943 7395
rect 7849 7293 7883 7327
rect 9505 7293 9539 7327
rect 9689 7293 9723 7327
rect 10425 7293 10459 7327
rect 12265 7293 12299 7327
rect 12817 7293 12851 7327
rect 13277 7293 13311 7327
rect 14105 7293 14139 7327
rect 14289 7293 14323 7327
rect 3893 7225 3927 7259
rect 9229 7225 9263 7259
rect 10609 7225 10643 7259
rect 8309 6953 8343 6987
rect 8677 6953 8711 6987
rect 10885 6953 10919 6987
rect 10333 6885 10367 6919
rect 4261 6817 4295 6851
rect 4905 6817 4939 6851
rect 5181 6817 5215 6851
rect 5825 6817 5859 6851
rect 5917 6817 5951 6851
rect 6101 6817 6135 6851
rect 9873 6817 9907 6851
rect 10437 6817 10471 6851
rect 11161 6817 11195 6851
rect 15945 6817 15979 6851
rect 16037 6817 16071 6851
rect 5273 6749 5307 6783
rect 8125 6749 8159 6783
rect 8217 6749 8251 6783
rect 10517 6749 10551 6783
rect 16221 6749 16255 6783
rect 5733 6681 5767 6715
rect 10885 6681 10919 6715
rect 10977 6681 11011 6715
rect 21925 6681 21959 6715
rect 15577 6613 15611 6647
rect 6837 6341 6871 6375
rect 6929 6341 6963 6375
rect 17233 6273 17267 6307
rect 17417 6273 17451 6307
rect 3490 6205 3524 6239
rect 5549 6205 5583 6239
rect 6101 6205 6135 6239
rect 6469 6205 6503 6239
rect 7113 6205 7147 6239
rect 17601 6205 17635 6239
rect 17785 6205 17819 6239
rect 18153 6205 18187 6239
rect 18337 6205 18371 6239
rect 18521 6205 18555 6239
rect 5641 6137 5675 6171
rect 3387 6069 3421 6103
rect 6837 6069 6871 6103
rect 18521 6069 18555 6103
rect 6929 5865 6963 5899
rect 16129 5865 16163 5899
rect 17509 5865 17543 5899
rect 21281 5865 21315 5899
rect 21925 5865 21959 5899
rect 1593 5797 1627 5831
rect 12725 5797 12759 5831
rect 2789 5729 2823 5763
rect 7021 5729 7055 5763
rect 14565 5729 14599 5763
rect 15117 5729 15151 5763
rect 15577 5729 15611 5763
rect 16497 5729 16531 5763
rect 17417 5729 17451 5763
rect 17785 5729 17819 5763
rect 17877 5729 17911 5763
rect 18521 5729 18555 5763
rect 18705 5729 18739 5763
rect 19073 5729 19107 5763
rect 21465 5729 21499 5763
rect 15209 5661 15243 5695
rect 16589 5661 16623 5695
rect 16773 5661 16807 5695
rect 18153 5661 18187 5695
rect 18337 5661 18371 5695
rect 18981 5661 19015 5695
rect 12541 5593 12575 5627
rect 1501 5525 1535 5559
rect 2697 5525 2731 5559
rect 14565 5525 14599 5559
rect 15209 5525 15243 5559
rect 8125 5321 8159 5355
rect 8585 5321 8619 5355
rect 13001 5321 13035 5355
rect 13461 5321 13495 5355
rect 15117 5321 15151 5355
rect 16957 5321 16991 5355
rect 18061 5321 18095 5355
rect 3249 5185 3283 5219
rect 8217 5185 8251 5219
rect 17601 5185 17635 5219
rect 2973 5117 3007 5151
rect 4997 5117 5031 5151
rect 7573 5117 7607 5151
rect 8125 5117 8159 5151
rect 8585 5117 8619 5151
rect 10333 5117 10367 5151
rect 12265 5117 12299 5151
rect 12449 5117 12483 5151
rect 13001 5117 13035 5151
rect 13093 5117 13127 5151
rect 13461 5117 13495 5151
rect 14565 5117 14599 5151
rect 14749 5117 14783 5151
rect 15301 5117 15335 5151
rect 18153 5117 18187 5151
rect 11069 5049 11103 5083
rect 11253 5049 11287 5083
rect 12081 5049 12115 5083
rect 17325 4981 17359 5015
rect 17417 4981 17451 5015
rect 7849 4777 7883 4811
rect 9873 4777 9907 4811
rect 10241 4777 10275 4811
rect 17969 4777 18003 4811
rect 8217 4709 8251 4743
rect 11161 4709 11195 4743
rect 18429 4709 18463 4743
rect 4997 4641 5031 4675
rect 7021 4641 7055 4675
rect 10517 4641 10551 4675
rect 11437 4641 11471 4675
rect 18337 4641 18371 4675
rect 6745 4573 6779 4607
rect 8309 4573 8343 4607
rect 8493 4573 8527 4607
rect 9597 4573 9631 4607
rect 9781 4573 9815 4607
rect 18613 4573 18647 4607
rect 15393 4165 15427 4199
rect 15577 3961 15611 3995
rect 8861 3689 8895 3723
rect 9321 3689 9355 3723
rect 11345 3689 11379 3723
rect 11437 3689 11471 3723
rect 13921 3689 13955 3723
rect 14841 3689 14875 3723
rect 15117 3689 15151 3723
rect 3985 3621 4019 3655
rect 9137 3621 9171 3655
rect 11621 3621 11655 3655
rect 6745 3553 6779 3587
rect 7021 3553 7055 3587
rect 11897 3553 11931 3587
rect 15025 3553 15059 3587
rect 15117 3553 15151 3587
rect 8493 3485 8527 3519
rect 10977 3485 11011 3519
rect 13553 3485 13587 3519
rect 15485 3485 15519 3519
rect 4169 3417 4203 3451
rect 8861 3417 8895 3451
rect 11345 3417 11379 3451
rect 11713 3417 11747 3451
rect 13921 3417 13955 3451
rect 9045 3145 9079 3179
rect 9781 3145 9815 3179
rect 11437 3145 11471 3179
rect 12633 3145 12667 3179
rect 13829 3145 13863 3179
rect 14565 3145 14599 3179
rect 14933 3145 14967 3179
rect 15577 3145 15611 3179
rect 17220 3145 17254 3179
rect 19165 3145 19199 3179
rect 14473 3077 14507 3111
rect 8493 3009 8527 3043
rect 9505 3009 9539 3043
rect 12265 3009 12299 3043
rect 13277 3009 13311 3043
rect 16129 3009 16163 3043
rect 16957 3009 16991 3043
rect 20913 3009 20947 3043
rect 21189 3009 21223 3043
rect 1409 2941 1443 2975
rect 8677 2941 8711 2975
rect 9137 2941 9171 2975
rect 9689 2941 9723 2975
rect 9965 2941 9999 2975
rect 10885 2941 10919 2975
rect 11437 2941 11471 2975
rect 12081 2941 12115 2975
rect 12541 2941 12575 2975
rect 13461 2941 13495 2975
rect 13921 2941 13955 2975
rect 14473 2941 14507 2975
rect 14749 2941 14783 2975
rect 14933 2941 14967 2975
rect 15485 2941 15519 2975
rect 15945 2941 15979 2975
rect 18981 2941 19015 2975
rect 21465 2941 21499 2975
rect 1593 2805 1627 2839
rect 8585 2805 8619 2839
rect 11713 2805 11747 2839
rect 12173 2805 12207 2839
rect 13369 2805 13403 2839
rect 16037 2805 16071 2839
rect 21281 2805 21315 2839
rect 4077 2601 4111 2635
rect 5733 2601 5767 2635
rect 7021 2601 7055 2635
rect 8953 2601 8987 2635
rect 12173 2601 12207 2635
rect 13829 2601 13863 2635
rect 17417 2601 17451 2635
rect 18889 2601 18923 2635
rect 21281 2601 21315 2635
rect 2053 2533 2087 2567
rect 1409 2465 1443 2499
rect 3893 2465 3927 2499
rect 5549 2465 5583 2499
rect 7113 2465 7147 2499
rect 8769 2465 8803 2499
rect 10701 2465 10735 2499
rect 11989 2465 12023 2499
rect 14013 2465 14047 2499
rect 15669 2465 15703 2499
rect 17325 2465 17359 2499
rect 19073 2465 19107 2499
rect 20913 2465 20947 2499
rect 21465 2465 21499 2499
rect 16129 2397 16163 2431
rect 1593 2329 1627 2363
rect 1869 2329 1903 2363
rect 10885 2329 10919 2363
rect 20729 2329 20763 2363
<< metal1 >>
rect 1104 22874 21804 22896
rect 1104 22822 4432 22874
rect 4484 22822 4496 22874
rect 4548 22822 4560 22874
rect 4612 22822 4624 22874
rect 4676 22822 11332 22874
rect 11384 22822 11396 22874
rect 11448 22822 11460 22874
rect 11512 22822 11524 22874
rect 11576 22822 18232 22874
rect 18284 22822 18296 22874
rect 18348 22822 18360 22874
rect 18412 22822 18424 22874
rect 18476 22822 21804 22874
rect 1104 22800 21804 22822
rect 1486 22760 1492 22772
rect 1447 22732 1492 22760
rect 1486 22720 1492 22732
rect 1544 22720 1550 22772
rect 2961 22695 3019 22701
rect 2961 22661 2973 22695
rect 3007 22692 3019 22695
rect 4890 22692 4896 22704
rect 3007 22664 4896 22692
rect 3007 22661 3019 22664
rect 2961 22655 3019 22661
rect 4890 22652 4896 22664
rect 4948 22652 4954 22704
rect 8021 22695 8079 22701
rect 8021 22661 8033 22695
rect 8067 22692 8079 22695
rect 11790 22692 11796 22704
rect 8067 22664 11796 22692
rect 8067 22661 8079 22664
rect 8021 22655 8079 22661
rect 11790 22652 11796 22664
rect 11848 22652 11854 22704
rect 934 22516 940 22568
rect 992 22556 998 22568
rect 1765 22559 1823 22565
rect 1765 22556 1777 22559
rect 992 22528 1777 22556
rect 992 22516 998 22528
rect 1765 22525 1777 22528
rect 1811 22525 1823 22559
rect 2774 22556 2780 22568
rect 2735 22528 2780 22556
rect 1765 22519 1823 22525
rect 2774 22516 2780 22528
rect 2832 22516 2838 22568
rect 4617 22559 4675 22565
rect 4617 22525 4629 22559
rect 4663 22556 4675 22559
rect 4798 22556 4804 22568
rect 4663 22528 4804 22556
rect 4663 22525 4675 22528
rect 4617 22519 4675 22525
rect 4798 22516 4804 22528
rect 4856 22516 4862 22568
rect 5994 22556 6000 22568
rect 5955 22528 6000 22556
rect 5994 22516 6000 22528
rect 6052 22516 6058 22568
rect 7834 22556 7840 22568
rect 7795 22528 7840 22556
rect 7834 22516 7840 22528
rect 7892 22516 7898 22568
rect 9674 22556 9680 22568
rect 9635 22528 9680 22556
rect 9674 22516 9680 22528
rect 9732 22516 9738 22568
rect 11698 22556 11704 22568
rect 11659 22528 11704 22556
rect 11698 22516 11704 22528
rect 11756 22516 11762 22568
rect 12894 22556 12900 22568
rect 12855 22528 12900 22556
rect 12894 22516 12900 22528
rect 12952 22516 12958 22568
rect 14734 22516 14740 22568
rect 14792 22556 14798 22568
rect 14921 22559 14979 22565
rect 14921 22556 14933 22559
rect 14792 22528 14933 22556
rect 14792 22516 14798 22528
rect 14921 22525 14933 22528
rect 14967 22525 14979 22559
rect 14921 22519 14979 22525
rect 16574 22516 16580 22568
rect 16632 22556 16638 22568
rect 16761 22559 16819 22565
rect 16761 22556 16773 22559
rect 16632 22528 16773 22556
rect 16632 22516 16638 22528
rect 16761 22525 16773 22528
rect 16807 22525 16819 22559
rect 16761 22519 16819 22525
rect 17954 22516 17960 22568
rect 18012 22556 18018 22568
rect 18141 22559 18199 22565
rect 18141 22556 18153 22559
rect 18012 22528 18153 22556
rect 18012 22516 18018 22528
rect 18141 22525 18153 22528
rect 18187 22525 18199 22559
rect 18141 22519 18199 22525
rect 19794 22516 19800 22568
rect 19852 22556 19858 22568
rect 20073 22559 20131 22565
rect 20073 22556 20085 22559
rect 19852 22528 20085 22556
rect 19852 22516 19858 22528
rect 20073 22525 20085 22528
rect 20119 22525 20131 22559
rect 21082 22556 21088 22568
rect 21043 22528 21088 22556
rect 20073 22519 20131 22525
rect 21082 22516 21088 22528
rect 21140 22516 21146 22568
rect 21453 22559 21511 22565
rect 21453 22525 21465 22559
rect 21499 22556 21511 22559
rect 21634 22556 21640 22568
rect 21499 22528 21640 22556
rect 21499 22525 21511 22528
rect 21453 22519 21511 22525
rect 21634 22516 21640 22528
rect 21692 22516 21698 22568
rect 1578 22488 1584 22500
rect 1539 22460 1584 22488
rect 1578 22448 1584 22460
rect 1636 22448 1642 22500
rect 1949 22423 2007 22429
rect 1949 22389 1961 22423
rect 1995 22420 2007 22423
rect 2038 22420 2044 22432
rect 1995 22392 2044 22420
rect 1995 22389 2007 22392
rect 1949 22383 2007 22389
rect 2038 22380 2044 22392
rect 2096 22380 2102 22432
rect 4798 22420 4804 22432
rect 4759 22392 4804 22420
rect 4798 22380 4804 22392
rect 4856 22380 4862 22432
rect 6181 22423 6239 22429
rect 6181 22389 6193 22423
rect 6227 22420 6239 22423
rect 6362 22420 6368 22432
rect 6227 22392 6368 22420
rect 6227 22389 6239 22392
rect 6181 22383 6239 22389
rect 6362 22380 6368 22392
rect 6420 22380 6426 22432
rect 9674 22380 9680 22432
rect 9732 22420 9738 22432
rect 9861 22423 9919 22429
rect 9861 22420 9873 22423
rect 9732 22392 9873 22420
rect 9732 22380 9738 22392
rect 9861 22389 9873 22392
rect 9907 22389 9919 22423
rect 9861 22383 9919 22389
rect 11146 22380 11152 22432
rect 11204 22420 11210 22432
rect 11517 22423 11575 22429
rect 11517 22420 11529 22423
rect 11204 22392 11529 22420
rect 11204 22380 11210 22392
rect 11517 22389 11529 22392
rect 11563 22389 11575 22423
rect 13078 22420 13084 22432
rect 13039 22392 13084 22420
rect 11517 22383 11575 22389
rect 13078 22380 13084 22392
rect 13136 22380 13142 22432
rect 14550 22380 14556 22432
rect 14608 22420 14614 22432
rect 14737 22423 14795 22429
rect 14737 22420 14749 22423
rect 14608 22392 14749 22420
rect 14608 22380 14614 22392
rect 14737 22389 14749 22392
rect 14783 22389 14795 22423
rect 14737 22383 14795 22389
rect 16577 22423 16635 22429
rect 16577 22389 16589 22423
rect 16623 22420 16635 22423
rect 16758 22420 16764 22432
rect 16623 22392 16764 22420
rect 16623 22389 16635 22392
rect 16577 22383 16635 22389
rect 16758 22380 16764 22392
rect 16816 22380 16822 22432
rect 17954 22420 17960 22432
rect 17915 22392 17960 22420
rect 17954 22380 17960 22392
rect 18012 22380 18018 22432
rect 19610 22380 19616 22432
rect 19668 22420 19674 22432
rect 19889 22423 19947 22429
rect 19889 22420 19901 22423
rect 19668 22392 19901 22420
rect 19668 22380 19674 22392
rect 19889 22389 19901 22392
rect 19935 22389 19947 22423
rect 20898 22420 20904 22432
rect 20859 22392 20904 22420
rect 19889 22383 19947 22389
rect 20898 22380 20904 22392
rect 20956 22380 20962 22432
rect 20990 22380 20996 22432
rect 21048 22420 21054 22432
rect 21269 22423 21327 22429
rect 21269 22420 21281 22423
rect 21048 22392 21281 22420
rect 21048 22380 21054 22392
rect 21269 22389 21281 22392
rect 21315 22389 21327 22423
rect 21269 22383 21327 22389
rect 1104 22330 21804 22352
rect 1104 22278 7882 22330
rect 7934 22278 7946 22330
rect 7998 22278 8010 22330
rect 8062 22278 8074 22330
rect 8126 22278 14782 22330
rect 14834 22278 14846 22330
rect 14898 22278 14910 22330
rect 14962 22278 14974 22330
rect 15026 22278 21804 22330
rect 1104 22256 21804 22278
rect 15470 22176 15476 22228
rect 15528 22216 15534 22228
rect 20898 22216 20904 22228
rect 15528 22188 20904 22216
rect 15528 22176 15534 22188
rect 20898 22176 20904 22188
rect 20956 22176 20962 22228
rect 4908 22120 5672 22148
rect 3694 22040 3700 22092
rect 3752 22080 3758 22092
rect 4908 22080 4936 22120
rect 5644 22094 5672 22120
rect 3752 22052 4936 22080
rect 4985 22083 5043 22089
rect 3752 22040 3758 22052
rect 4985 22049 4997 22083
rect 5031 22049 5043 22083
rect 4985 22043 5043 22049
rect 5077 22083 5135 22089
rect 5077 22049 5089 22083
rect 5123 22080 5135 22083
rect 5258 22080 5264 22092
rect 5123 22052 5264 22080
rect 5123 22049 5135 22052
rect 5077 22043 5135 22049
rect 5000 22012 5028 22043
rect 5258 22040 5264 22052
rect 5316 22040 5322 22092
rect 5353 22083 5411 22089
rect 5353 22049 5365 22083
rect 5399 22080 5411 22083
rect 5534 22080 5540 22092
rect 5399 22052 5540 22080
rect 5399 22049 5411 22052
rect 5353 22043 5411 22049
rect 5534 22040 5540 22052
rect 5592 22040 5598 22092
rect 5644 22089 5709 22094
rect 5629 22083 5709 22089
rect 5629 22049 5641 22083
rect 5675 22080 5709 22083
rect 7561 22083 7619 22089
rect 7561 22080 7573 22083
rect 5675 22052 7573 22080
rect 5675 22049 5687 22052
rect 5629 22043 5687 22049
rect 7561 22049 7573 22052
rect 7607 22080 7619 22083
rect 9861 22083 9919 22089
rect 9861 22080 9873 22083
rect 7607 22052 9873 22080
rect 7607 22049 7619 22052
rect 7561 22043 7619 22049
rect 9861 22049 9873 22052
rect 9907 22080 9919 22083
rect 10318 22080 10324 22092
rect 9907 22052 10324 22080
rect 9907 22049 9919 22052
rect 9861 22043 9919 22049
rect 10318 22040 10324 22052
rect 10376 22040 10382 22092
rect 11698 22080 11704 22092
rect 11659 22052 11704 22080
rect 11698 22040 11704 22052
rect 11756 22040 11762 22092
rect 11882 22080 11888 22092
rect 11843 22052 11888 22080
rect 11882 22040 11888 22052
rect 11940 22040 11946 22092
rect 11974 22040 11980 22092
rect 12032 22080 12038 22092
rect 12115 22083 12173 22089
rect 12032 22052 12077 22080
rect 12032 22040 12038 22052
rect 12115 22049 12127 22083
rect 12161 22080 12173 22083
rect 12342 22080 12348 22092
rect 12161 22052 12348 22080
rect 12161 22049 12173 22052
rect 12115 22043 12173 22049
rect 12342 22040 12348 22052
rect 12400 22040 12406 22092
rect 12713 22083 12771 22089
rect 12713 22049 12725 22083
rect 12759 22080 12771 22083
rect 15197 22083 15255 22089
rect 15197 22080 15209 22083
rect 12759 22052 15209 22080
rect 12759 22049 12771 22052
rect 12713 22043 12771 22049
rect 15197 22049 15209 22052
rect 15243 22080 15255 22083
rect 17126 22080 17132 22092
rect 15243 22052 17132 22080
rect 15243 22049 15255 22052
rect 15197 22043 15255 22049
rect 5810 22012 5816 22024
rect 5000 21984 5816 22012
rect 5810 21972 5816 21984
rect 5868 21972 5874 22024
rect 10336 22012 10364 22040
rect 12728 22012 12756 22043
rect 17126 22040 17132 22052
rect 17184 22080 17190 22092
rect 18325 22083 18383 22089
rect 18325 22080 18337 22083
rect 17184 22052 18337 22080
rect 17184 22040 17190 22052
rect 18325 22049 18337 22052
rect 18371 22080 18383 22083
rect 19981 22083 20039 22089
rect 19981 22080 19993 22083
rect 18371 22052 19993 22080
rect 18371 22049 18383 22052
rect 18325 22043 18383 22049
rect 19981 22049 19993 22052
rect 20027 22049 20039 22083
rect 19981 22043 20039 22049
rect 10336 21984 12756 22012
rect 4154 21836 4160 21888
rect 4212 21876 4218 21888
rect 4801 21879 4859 21885
rect 4801 21876 4813 21879
rect 4212 21848 4813 21876
rect 4212 21836 4218 21848
rect 4801 21845 4813 21848
rect 4847 21845 4859 21879
rect 4801 21839 4859 21845
rect 4982 21836 4988 21888
rect 5040 21876 5046 21888
rect 5261 21879 5319 21885
rect 5261 21876 5273 21879
rect 5040 21848 5273 21876
rect 5040 21836 5046 21848
rect 5261 21845 5273 21848
rect 5307 21845 5319 21879
rect 5442 21876 5448 21888
rect 5403 21848 5448 21876
rect 5261 21839 5319 21845
rect 5442 21836 5448 21848
rect 5500 21836 5506 21888
rect 7650 21836 7656 21888
rect 7708 21876 7714 21888
rect 7745 21879 7803 21885
rect 7745 21876 7757 21879
rect 7708 21848 7757 21876
rect 7708 21836 7714 21848
rect 7745 21845 7757 21848
rect 7791 21845 7803 21879
rect 10042 21876 10048 21888
rect 10003 21848 10048 21876
rect 7745 21839 7803 21845
rect 10042 21836 10048 21848
rect 10100 21836 10106 21888
rect 12066 21836 12072 21888
rect 12124 21876 12130 21888
rect 12253 21879 12311 21885
rect 12253 21876 12265 21879
rect 12124 21848 12265 21876
rect 12124 21836 12130 21848
rect 12253 21845 12265 21848
rect 12299 21845 12311 21879
rect 12253 21839 12311 21845
rect 12802 21836 12808 21888
rect 12860 21876 12866 21888
rect 12897 21879 12955 21885
rect 12897 21876 12909 21879
rect 12860 21848 12909 21876
rect 12860 21836 12866 21848
rect 12897 21845 12909 21848
rect 12943 21845 12955 21879
rect 12897 21839 12955 21845
rect 15286 21836 15292 21888
rect 15344 21876 15350 21888
rect 15381 21879 15439 21885
rect 15381 21876 15393 21879
rect 15344 21848 15393 21876
rect 15344 21836 15350 21848
rect 15381 21845 15393 21848
rect 15427 21845 15439 21879
rect 15381 21839 15439 21845
rect 18509 21879 18567 21885
rect 18509 21845 18521 21879
rect 18555 21876 18567 21879
rect 18690 21876 18696 21888
rect 18555 21848 18696 21876
rect 18555 21845 18567 21848
rect 18509 21839 18567 21845
rect 18690 21836 18696 21848
rect 18748 21836 18754 21888
rect 20162 21876 20168 21888
rect 20123 21848 20168 21876
rect 20162 21836 20168 21848
rect 20220 21836 20226 21888
rect 1104 21786 21804 21808
rect 1104 21734 4432 21786
rect 4484 21734 4496 21786
rect 4548 21734 4560 21786
rect 4612 21734 4624 21786
rect 4676 21734 11332 21786
rect 11384 21734 11396 21786
rect 11448 21734 11460 21786
rect 11512 21734 11524 21786
rect 11576 21734 18232 21786
rect 18284 21734 18296 21786
rect 18348 21734 18360 21786
rect 18412 21734 18424 21786
rect 18476 21734 21804 21786
rect 1104 21712 21804 21734
rect 1578 21632 1584 21684
rect 1636 21672 1642 21684
rect 1765 21675 1823 21681
rect 1765 21672 1777 21675
rect 1636 21644 1777 21672
rect 1636 21632 1642 21644
rect 1765 21641 1777 21644
rect 1811 21641 1823 21675
rect 1765 21635 1823 21641
rect 5534 21632 5540 21684
rect 5592 21672 5598 21684
rect 5629 21675 5687 21681
rect 5629 21672 5641 21675
rect 5592 21644 5641 21672
rect 5592 21632 5598 21644
rect 5629 21641 5641 21644
rect 5675 21641 5687 21675
rect 5810 21672 5816 21684
rect 5771 21644 5816 21672
rect 5629 21635 5687 21641
rect 4154 21536 4160 21548
rect 4115 21508 4160 21536
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 1949 21471 2007 21477
rect 1949 21437 1961 21471
rect 1995 21468 2007 21471
rect 2498 21468 2504 21480
rect 1995 21440 2504 21468
rect 1995 21437 2007 21440
rect 1949 21431 2007 21437
rect 2498 21428 2504 21440
rect 2556 21468 2562 21480
rect 3881 21471 3939 21477
rect 3881 21468 3893 21471
rect 2556 21440 3893 21468
rect 2556 21428 2562 21440
rect 3881 21437 3893 21440
rect 3927 21437 3939 21471
rect 5644 21468 5672 21635
rect 5810 21632 5816 21644
rect 5868 21632 5874 21684
rect 16574 21672 16580 21684
rect 11808 21644 16580 21672
rect 9030 21536 9036 21548
rect 6656 21508 9036 21536
rect 6656 21477 6684 21508
rect 9030 21496 9036 21508
rect 9088 21496 9094 21548
rect 9309 21539 9367 21545
rect 9309 21505 9321 21539
rect 9355 21536 9367 21539
rect 10873 21539 10931 21545
rect 10873 21536 10885 21539
rect 9355 21508 10885 21536
rect 9355 21505 9367 21508
rect 9309 21499 9367 21505
rect 10873 21505 10885 21508
rect 10919 21505 10931 21539
rect 10873 21499 10931 21505
rect 11808 21477 11836 21644
rect 12066 21536 12072 21548
rect 12027 21508 12072 21536
rect 12066 21496 12072 21508
rect 12124 21496 12130 21548
rect 14200 21536 14228 21644
rect 16574 21632 16580 21644
rect 16632 21632 16638 21684
rect 14277 21539 14335 21545
rect 14277 21536 14289 21539
rect 14200 21508 14289 21536
rect 14277 21505 14289 21508
rect 14323 21505 14335 21539
rect 14277 21499 14335 21505
rect 15102 21496 15108 21548
rect 15160 21536 15166 21548
rect 16025 21539 16083 21545
rect 16025 21536 16037 21539
rect 15160 21508 16037 21536
rect 15160 21496 15166 21508
rect 16025 21505 16037 21508
rect 16071 21505 16083 21539
rect 16025 21499 16083 21505
rect 16574 21496 16580 21548
rect 16632 21536 16638 21548
rect 17405 21539 17463 21545
rect 17405 21536 17417 21539
rect 16632 21508 17417 21536
rect 16632 21496 16638 21508
rect 17405 21505 17417 21508
rect 17451 21536 17463 21539
rect 17770 21536 17776 21548
rect 17451 21508 17776 21536
rect 17451 21505 17463 21508
rect 17405 21499 17463 21505
rect 17770 21496 17776 21508
rect 17828 21536 17834 21548
rect 19153 21539 19211 21545
rect 17828 21508 18920 21536
rect 17828 21496 17834 21508
rect 5721 21471 5779 21477
rect 5721 21468 5733 21471
rect 5644 21440 5733 21468
rect 3881 21431 3939 21437
rect 5721 21437 5733 21440
rect 5767 21437 5779 21471
rect 6641 21471 6699 21477
rect 6641 21468 6653 21471
rect 5721 21431 5779 21437
rect 6564 21440 6653 21468
rect 3896 21332 3924 21431
rect 5442 21400 5448 21412
rect 5382 21372 5448 21400
rect 5442 21360 5448 21372
rect 5500 21360 5506 21412
rect 6564 21332 6592 21440
rect 6641 21437 6653 21440
rect 6687 21437 6699 21471
rect 11793 21471 11851 21477
rect 11793 21468 11805 21471
rect 6641 21431 6699 21437
rect 10612 21440 11805 21468
rect 6917 21403 6975 21409
rect 6917 21369 6929 21403
rect 6963 21400 6975 21403
rect 7190 21400 7196 21412
rect 6963 21372 7196 21400
rect 6963 21369 6975 21372
rect 6917 21363 6975 21369
rect 7190 21360 7196 21372
rect 7248 21360 7254 21412
rect 7650 21360 7656 21412
rect 7708 21360 7714 21412
rect 10042 21360 10048 21412
rect 10100 21360 10106 21412
rect 3896 21304 6592 21332
rect 7742 21292 7748 21344
rect 7800 21332 7806 21344
rect 8389 21335 8447 21341
rect 8389 21332 8401 21335
rect 7800 21304 8401 21332
rect 7800 21292 7806 21304
rect 8389 21301 8401 21304
rect 8435 21301 8447 21335
rect 8389 21295 8447 21301
rect 9030 21292 9036 21344
rect 9088 21332 9094 21344
rect 10612 21332 10640 21440
rect 11793 21437 11805 21440
rect 11839 21437 11851 21471
rect 17126 21468 17132 21480
rect 17087 21440 17132 21468
rect 11793 21431 11851 21437
rect 17126 21428 17132 21440
rect 17184 21428 17190 21480
rect 18892 21468 18920 21508
rect 19153 21505 19165 21539
rect 19199 21536 19211 21539
rect 19521 21539 19579 21545
rect 19521 21536 19533 21539
rect 19199 21508 19533 21536
rect 19199 21505 19211 21508
rect 19153 21499 19211 21505
rect 19521 21505 19533 21508
rect 19567 21505 19579 21539
rect 19521 21499 19579 21505
rect 19245 21471 19303 21477
rect 19245 21468 19257 21471
rect 18892 21440 19257 21468
rect 19245 21437 19257 21440
rect 19291 21437 19303 21471
rect 19245 21431 19303 21437
rect 11057 21403 11115 21409
rect 11057 21369 11069 21403
rect 11103 21369 11115 21403
rect 11238 21400 11244 21412
rect 11199 21372 11244 21400
rect 11057 21363 11115 21369
rect 9088 21304 10640 21332
rect 10781 21335 10839 21341
rect 9088 21292 9094 21304
rect 10781 21301 10793 21335
rect 10827 21332 10839 21335
rect 11072 21332 11100 21363
rect 11238 21360 11244 21372
rect 11296 21360 11302 21412
rect 12802 21360 12808 21412
rect 12860 21360 12866 21412
rect 14553 21403 14611 21409
rect 14553 21369 14565 21403
rect 14599 21400 14611 21403
rect 14642 21400 14648 21412
rect 14599 21372 14648 21400
rect 14599 21369 14611 21372
rect 14553 21363 14611 21369
rect 14642 21360 14648 21372
rect 14700 21360 14706 21412
rect 15286 21360 15292 21412
rect 15344 21360 15350 21412
rect 17681 21403 17739 21409
rect 17681 21369 17693 21403
rect 17727 21400 17739 21403
rect 17954 21400 17960 21412
rect 17727 21372 17960 21400
rect 17727 21369 17739 21372
rect 17681 21363 17739 21369
rect 17954 21360 17960 21372
rect 18012 21360 18018 21412
rect 18690 21360 18696 21412
rect 18748 21360 18754 21412
rect 20162 21360 20168 21412
rect 20220 21360 20226 21412
rect 11882 21332 11888 21344
rect 10827 21304 11888 21332
rect 10827 21301 10839 21304
rect 10781 21295 10839 21301
rect 11882 21292 11888 21304
rect 11940 21292 11946 21344
rect 13538 21332 13544 21344
rect 13499 21304 13544 21332
rect 13538 21292 13544 21304
rect 13596 21292 13602 21344
rect 17218 21292 17224 21344
rect 17276 21332 17282 21344
rect 17313 21335 17371 21341
rect 17313 21332 17325 21335
rect 17276 21304 17325 21332
rect 17276 21292 17282 21304
rect 17313 21301 17325 21304
rect 17359 21301 17371 21335
rect 17313 21295 17371 21301
rect 20898 21292 20904 21344
rect 20956 21332 20962 21344
rect 20993 21335 21051 21341
rect 20993 21332 21005 21335
rect 20956 21304 21005 21332
rect 20956 21292 20962 21304
rect 20993 21301 21005 21304
rect 21039 21301 21051 21335
rect 20993 21295 21051 21301
rect 1104 21242 21804 21264
rect 1104 21190 7882 21242
rect 7934 21190 7946 21242
rect 7998 21190 8010 21242
rect 8062 21190 8074 21242
rect 8126 21190 14782 21242
rect 14834 21190 14846 21242
rect 14898 21190 14910 21242
rect 14962 21190 14974 21242
rect 15026 21190 21804 21242
rect 1104 21168 21804 21190
rect 7190 21128 7196 21140
rect 7151 21100 7196 21128
rect 7190 21088 7196 21100
rect 7248 21088 7254 21140
rect 8294 21128 8300 21140
rect 7576 21100 8300 21128
rect 7466 21060 7472 21072
rect 7427 21032 7472 21060
rect 7466 21020 7472 21032
rect 7524 21020 7530 21072
rect 7576 21069 7604 21100
rect 8294 21088 8300 21100
rect 8352 21088 8358 21140
rect 11974 21088 11980 21140
rect 12032 21128 12038 21140
rect 14642 21128 14648 21140
rect 12032 21100 12112 21128
rect 14603 21100 14648 21128
rect 12032 21088 12038 21100
rect 7742 21069 7748 21072
rect 7561 21063 7619 21069
rect 7561 21029 7573 21063
rect 7607 21029 7619 21063
rect 7561 21023 7619 21029
rect 7699 21063 7748 21069
rect 7699 21029 7711 21063
rect 7745 21029 7748 21063
rect 7699 21023 7748 21029
rect 7742 21020 7748 21023
rect 7800 21020 7806 21072
rect 12084 21069 12112 21100
rect 14642 21088 14648 21100
rect 14700 21088 14706 21140
rect 12069 21063 12127 21069
rect 12069 21029 12081 21063
rect 12115 21060 12127 21063
rect 12618 21060 12624 21072
rect 12115 21032 12624 21060
rect 12115 21029 12127 21032
rect 12069 21023 12127 21029
rect 12618 21020 12624 21032
rect 12676 21060 12682 21072
rect 13538 21060 13544 21072
rect 12676 21032 13544 21060
rect 12676 21020 12682 21032
rect 13538 21020 13544 21032
rect 13596 21020 13602 21072
rect 14921 21063 14979 21069
rect 14921 21029 14933 21063
rect 14967 21060 14979 21063
rect 15102 21060 15108 21072
rect 14967 21032 15108 21060
rect 14967 21029 14979 21032
rect 14921 21023 14979 21029
rect 15102 21020 15108 21032
rect 15160 21020 15166 21072
rect 16574 21060 16580 21072
rect 16224 21032 16580 21060
rect 7374 20992 7380 21004
rect 7335 20964 7380 20992
rect 7374 20952 7380 20964
rect 7432 20952 7438 21004
rect 7837 20995 7895 21001
rect 7837 20961 7849 20995
rect 7883 20992 7895 20995
rect 8205 20995 8263 21001
rect 8205 20992 8217 20995
rect 7883 20964 8217 20992
rect 7883 20961 7895 20964
rect 7837 20955 7895 20961
rect 8205 20961 8217 20964
rect 8251 20992 8263 20995
rect 8846 20992 8852 21004
rect 8251 20964 8852 20992
rect 8251 20961 8263 20964
rect 8205 20955 8263 20961
rect 8846 20952 8852 20964
rect 8904 20952 8910 21004
rect 11238 20952 11244 21004
rect 11296 20992 11302 21004
rect 11698 20992 11704 21004
rect 11296 20964 11704 20992
rect 11296 20952 11302 20964
rect 11698 20952 11704 20964
rect 11756 20992 11762 21004
rect 11974 20992 11980 21004
rect 11756 20964 11980 20992
rect 11756 20952 11762 20964
rect 11974 20952 11980 20964
rect 12032 20952 12038 21004
rect 12158 20952 12164 21004
rect 12216 20992 12222 21004
rect 12342 20992 12348 21004
rect 12216 20964 12261 20992
rect 12303 20964 12348 20992
rect 12216 20952 12222 20964
rect 12342 20952 12348 20964
rect 12400 20992 12406 21004
rect 14829 20995 14887 21001
rect 14829 20992 14841 20995
rect 12400 20964 14841 20992
rect 12400 20952 12406 20964
rect 14829 20961 14841 20964
rect 14875 20961 14887 20995
rect 14829 20955 14887 20961
rect 15013 20995 15071 21001
rect 15013 20961 15025 20995
rect 15059 20961 15071 20995
rect 15194 20992 15200 21004
rect 15155 20964 15200 20992
rect 15013 20955 15071 20961
rect 14844 20856 14872 20955
rect 15028 20924 15056 20955
rect 15194 20952 15200 20964
rect 15252 20952 15258 21004
rect 16224 21001 16252 21032
rect 16574 21020 16580 21032
rect 16632 21020 16638 21072
rect 17218 21020 17224 21072
rect 17276 21020 17282 21072
rect 16209 20995 16267 21001
rect 16209 20961 16221 20995
rect 16255 20961 16267 20995
rect 16209 20955 16267 20961
rect 21082 20952 21088 21004
rect 21140 20992 21146 21004
rect 21269 20995 21327 21001
rect 21269 20992 21281 20995
rect 21140 20964 21281 20992
rect 21140 20952 21146 20964
rect 21269 20961 21281 20964
rect 21315 20961 21327 20995
rect 21269 20955 21327 20961
rect 15378 20924 15384 20936
rect 15028 20896 15384 20924
rect 15378 20884 15384 20896
rect 15436 20884 15442 20936
rect 16482 20924 16488 20936
rect 16443 20896 16488 20924
rect 16482 20884 16488 20896
rect 16540 20884 16546 20936
rect 15838 20856 15844 20868
rect 14844 20828 15844 20856
rect 15838 20816 15844 20828
rect 15896 20816 15902 20868
rect 8294 20788 8300 20800
rect 8207 20760 8300 20788
rect 8294 20748 8300 20760
rect 8352 20788 8358 20800
rect 9306 20788 9312 20800
rect 8352 20760 9312 20788
rect 8352 20748 8358 20760
rect 9306 20748 9312 20760
rect 9364 20748 9370 20800
rect 11054 20748 11060 20800
rect 11112 20788 11118 20800
rect 11793 20791 11851 20797
rect 11793 20788 11805 20791
rect 11112 20760 11805 20788
rect 11112 20748 11118 20760
rect 11793 20757 11805 20760
rect 11839 20757 11851 20791
rect 11793 20751 11851 20757
rect 15378 20748 15384 20800
rect 15436 20788 15442 20800
rect 17957 20791 18015 20797
rect 17957 20788 17969 20791
rect 15436 20760 17969 20788
rect 15436 20748 15442 20760
rect 17957 20757 17969 20760
rect 18003 20757 18015 20791
rect 21358 20788 21364 20800
rect 21319 20760 21364 20788
rect 17957 20751 18015 20757
rect 21358 20748 21364 20760
rect 21416 20748 21422 20800
rect 1104 20698 21804 20720
rect 1104 20646 4432 20698
rect 4484 20646 4496 20698
rect 4548 20646 4560 20698
rect 4612 20646 4624 20698
rect 4676 20646 11332 20698
rect 11384 20646 11396 20698
rect 11448 20646 11460 20698
rect 11512 20646 11524 20698
rect 11576 20646 18232 20698
rect 18284 20646 18296 20698
rect 18348 20646 18360 20698
rect 18412 20646 18424 20698
rect 18476 20646 21804 20698
rect 1104 20624 21804 20646
rect 11974 20476 11980 20528
rect 12032 20516 12038 20528
rect 12032 20488 12388 20516
rect 12032 20476 12038 20488
rect 9030 20408 9036 20460
rect 9088 20448 9094 20460
rect 9585 20451 9643 20457
rect 9585 20448 9597 20451
rect 9088 20420 9597 20448
rect 9088 20408 9094 20420
rect 9585 20417 9597 20420
rect 9631 20417 9643 20451
rect 9585 20411 9643 20417
rect 9861 20451 9919 20457
rect 9861 20417 9873 20451
rect 9907 20448 9919 20451
rect 11054 20448 11060 20460
rect 9907 20420 11060 20448
rect 9907 20417 9919 20420
rect 9861 20411 9919 20417
rect 11054 20408 11060 20420
rect 11112 20408 11118 20460
rect 11333 20451 11391 20457
rect 11333 20417 11345 20451
rect 11379 20448 11391 20451
rect 12360 20448 12388 20488
rect 15194 20448 15200 20460
rect 11379 20420 12112 20448
rect 11379 20417 11391 20420
rect 11333 20411 11391 20417
rect 1394 20380 1400 20392
rect 1355 20352 1400 20380
rect 1394 20340 1400 20352
rect 1452 20340 1458 20392
rect 2498 20380 2504 20392
rect 2459 20352 2504 20380
rect 2498 20340 2504 20352
rect 2556 20340 2562 20392
rect 5261 20383 5319 20389
rect 5261 20349 5273 20383
rect 5307 20349 5319 20383
rect 5261 20343 5319 20349
rect 5445 20383 5503 20389
rect 5445 20349 5457 20383
rect 5491 20380 5503 20383
rect 5534 20380 5540 20392
rect 5491 20352 5540 20380
rect 5491 20349 5503 20352
rect 5445 20343 5503 20349
rect 2777 20315 2835 20321
rect 2777 20281 2789 20315
rect 2823 20281 2835 20315
rect 2777 20275 2835 20281
rect 1486 20204 1492 20256
rect 1544 20244 1550 20256
rect 1581 20247 1639 20253
rect 1581 20244 1593 20247
rect 1544 20216 1593 20244
rect 1544 20204 1550 20216
rect 1581 20213 1593 20216
rect 1627 20213 1639 20247
rect 2792 20244 2820 20275
rect 3510 20272 3516 20324
rect 3568 20272 3574 20324
rect 5276 20312 5304 20343
rect 5534 20340 5540 20352
rect 5592 20340 5598 20392
rect 11882 20380 11888 20392
rect 11843 20352 11888 20380
rect 11882 20340 11888 20352
rect 11940 20340 11946 20392
rect 12084 20389 12112 20420
rect 12360 20420 15200 20448
rect 12069 20383 12127 20389
rect 12069 20349 12081 20383
rect 12115 20380 12127 20383
rect 12158 20380 12164 20392
rect 12115 20352 12164 20380
rect 12115 20349 12127 20352
rect 12069 20343 12127 20349
rect 12158 20340 12164 20352
rect 12216 20340 12222 20392
rect 12360 20389 12388 20420
rect 15194 20408 15200 20420
rect 15252 20448 15258 20460
rect 16390 20448 16396 20460
rect 15252 20420 16396 20448
rect 15252 20408 15258 20420
rect 16390 20408 16396 20420
rect 16448 20408 16454 20460
rect 12345 20383 12403 20389
rect 12345 20349 12357 20383
rect 12391 20349 12403 20383
rect 12526 20380 12532 20392
rect 12487 20352 12532 20380
rect 12345 20343 12403 20349
rect 12526 20340 12532 20352
rect 12584 20340 12590 20392
rect 12618 20340 12624 20392
rect 12676 20380 12682 20392
rect 15102 20380 15108 20392
rect 12676 20352 12721 20380
rect 15063 20352 15108 20380
rect 12676 20340 12682 20352
rect 15102 20340 15108 20352
rect 15160 20340 15166 20392
rect 20717 20383 20775 20389
rect 20717 20349 20729 20383
rect 20763 20349 20775 20383
rect 20717 20343 20775 20349
rect 20809 20383 20867 20389
rect 20809 20349 20821 20383
rect 20855 20380 20867 20383
rect 20898 20380 20904 20392
rect 20855 20352 20904 20380
rect 20855 20349 20867 20352
rect 20809 20343 20867 20349
rect 5276 20284 5488 20312
rect 5460 20256 5488 20284
rect 10502 20272 10508 20324
rect 10560 20272 10566 20324
rect 19702 20272 19708 20324
rect 19760 20312 19766 20324
rect 20165 20315 20223 20321
rect 20165 20312 20177 20315
rect 19760 20284 20177 20312
rect 19760 20272 19766 20284
rect 20165 20281 20177 20284
rect 20211 20281 20223 20315
rect 20732 20312 20760 20343
rect 20898 20340 20904 20352
rect 20956 20380 20962 20392
rect 21177 20383 21235 20389
rect 21177 20380 21189 20383
rect 20956 20352 21189 20380
rect 20956 20340 20962 20352
rect 21177 20349 21189 20352
rect 21223 20349 21235 20383
rect 21177 20343 21235 20349
rect 21269 20383 21327 20389
rect 21269 20349 21281 20383
rect 21315 20349 21327 20383
rect 21269 20343 21327 20349
rect 21284 20312 21312 20343
rect 21358 20312 21364 20324
rect 20732 20284 21364 20312
rect 20165 20275 20223 20281
rect 21358 20272 21364 20284
rect 21416 20272 21422 20324
rect 4154 20244 4160 20256
rect 2792 20216 4160 20244
rect 1581 20207 1639 20213
rect 4154 20204 4160 20216
rect 4212 20204 4218 20256
rect 4249 20247 4307 20253
rect 4249 20213 4261 20247
rect 4295 20244 4307 20247
rect 5166 20244 5172 20256
rect 4295 20216 5172 20244
rect 4295 20213 4307 20216
rect 4249 20207 4307 20213
rect 5166 20204 5172 20216
rect 5224 20204 5230 20256
rect 5350 20244 5356 20256
rect 5311 20216 5356 20244
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 5442 20204 5448 20256
rect 5500 20204 5506 20256
rect 15013 20247 15071 20253
rect 15013 20213 15025 20247
rect 15059 20244 15071 20247
rect 15102 20244 15108 20256
rect 15059 20216 15108 20244
rect 15059 20213 15071 20216
rect 15013 20207 15071 20213
rect 15102 20204 15108 20216
rect 15160 20204 15166 20256
rect 1104 20154 21804 20176
rect 1104 20102 7882 20154
rect 7934 20102 7946 20154
rect 7998 20102 8010 20154
rect 8062 20102 8074 20154
rect 8126 20102 14782 20154
rect 14834 20102 14846 20154
rect 14898 20102 14910 20154
rect 14962 20102 14974 20154
rect 15026 20102 21804 20154
rect 1104 20080 21804 20102
rect 3510 20040 3516 20052
rect 3471 20012 3516 20040
rect 3510 20000 3516 20012
rect 3568 20000 3574 20052
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 4709 20043 4767 20049
rect 4709 20040 4721 20043
rect 4212 20012 4721 20040
rect 4212 20000 4218 20012
rect 4709 20009 4721 20012
rect 4755 20009 4767 20043
rect 4709 20003 4767 20009
rect 5166 20000 5172 20052
rect 5224 20040 5230 20052
rect 5224 20012 5948 20040
rect 5224 20000 5230 20012
rect 5813 19975 5871 19981
rect 5813 19972 5825 19975
rect 4908 19944 5825 19972
rect 3694 19904 3700 19916
rect 3655 19876 3700 19904
rect 3694 19864 3700 19876
rect 3752 19864 3758 19916
rect 4908 19913 4936 19944
rect 5813 19941 5825 19944
rect 5859 19941 5871 19975
rect 5813 19935 5871 19941
rect 4893 19907 4951 19913
rect 4893 19873 4905 19907
rect 4939 19873 4951 19907
rect 4893 19867 4951 19873
rect 4985 19907 5043 19913
rect 4985 19873 4997 19907
rect 5031 19873 5043 19907
rect 4985 19867 5043 19873
rect 5077 19907 5135 19913
rect 5077 19873 5089 19907
rect 5123 19873 5135 19907
rect 5077 19867 5135 19873
rect 5000 19836 5028 19867
rect 4908 19808 5028 19836
rect 4908 19780 4936 19808
rect 4890 19728 4896 19780
rect 4948 19728 4954 19780
rect 4982 19728 4988 19780
rect 5040 19768 5046 19780
rect 5092 19768 5120 19867
rect 5166 19864 5172 19916
rect 5224 19913 5230 19916
rect 5224 19907 5253 19913
rect 5241 19873 5253 19907
rect 5442 19904 5448 19916
rect 5403 19876 5448 19904
rect 5224 19867 5253 19873
rect 5224 19864 5230 19867
rect 5442 19864 5448 19876
rect 5500 19864 5506 19916
rect 5534 19864 5540 19916
rect 5592 19904 5598 19916
rect 5920 19913 5948 20012
rect 7466 20000 7472 20052
rect 7524 20040 7530 20052
rect 7745 20043 7803 20049
rect 7745 20040 7757 20043
rect 7524 20012 7757 20040
rect 7524 20000 7530 20012
rect 7745 20009 7757 20012
rect 7791 20009 7803 20043
rect 8205 20043 8263 20049
rect 8205 20040 8217 20043
rect 7745 20003 7803 20009
rect 7852 20012 8217 20040
rect 7374 19932 7380 19984
rect 7432 19972 7438 19984
rect 7852 19972 7880 20012
rect 8205 20009 8217 20012
rect 8251 20009 8263 20043
rect 10502 20040 10508 20052
rect 10463 20012 10508 20040
rect 8205 20003 8263 20009
rect 10502 20000 10508 20012
rect 10560 20000 10566 20052
rect 15746 20040 15752 20052
rect 15304 20012 15752 20040
rect 15304 19981 15332 20012
rect 15746 20000 15752 20012
rect 15804 20000 15810 20052
rect 21358 20040 21364 20052
rect 21319 20012 21364 20040
rect 21358 20000 21364 20012
rect 21416 20000 21422 20052
rect 7432 19944 7880 19972
rect 7929 19975 7987 19981
rect 7432 19932 7438 19944
rect 7929 19941 7941 19975
rect 7975 19972 7987 19975
rect 15289 19975 15347 19981
rect 7975 19944 8248 19972
rect 7975 19941 7987 19944
rect 7929 19935 7987 19941
rect 8220 19916 8248 19944
rect 15289 19941 15301 19975
rect 15335 19941 15347 19975
rect 15289 19935 15347 19941
rect 15378 19932 15384 19984
rect 15436 19972 15442 19984
rect 15436 19944 15792 19972
rect 15436 19932 15442 19944
rect 5629 19907 5687 19913
rect 5629 19904 5641 19907
rect 5592 19876 5641 19904
rect 5592 19864 5598 19876
rect 5629 19873 5641 19876
rect 5675 19873 5687 19907
rect 5629 19867 5687 19873
rect 5905 19907 5963 19913
rect 5905 19873 5917 19907
rect 5951 19873 5963 19907
rect 5905 19867 5963 19873
rect 7742 19864 7748 19916
rect 7800 19904 7806 19916
rect 8113 19907 8171 19913
rect 8113 19904 8125 19907
rect 7800 19876 8125 19904
rect 7800 19864 7806 19876
rect 8113 19873 8125 19876
rect 8159 19873 8171 19907
rect 8113 19867 8171 19873
rect 5353 19839 5411 19845
rect 5353 19805 5365 19839
rect 5399 19805 5411 19839
rect 8128 19836 8156 19867
rect 8202 19864 8208 19916
rect 8260 19904 8266 19916
rect 8389 19907 8447 19913
rect 8260 19876 8305 19904
rect 8260 19864 8266 19876
rect 8389 19873 8401 19907
rect 8435 19873 8447 19907
rect 10318 19904 10324 19916
rect 10279 19876 10324 19904
rect 8389 19867 8447 19873
rect 8404 19836 8432 19867
rect 10318 19864 10324 19876
rect 10376 19864 10382 19916
rect 14458 19864 14464 19916
rect 14516 19904 14522 19916
rect 15102 19904 15108 19916
rect 14516 19876 15108 19904
rect 14516 19864 14522 19876
rect 15102 19864 15108 19876
rect 15160 19864 15166 19916
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 15764 19913 15792 19944
rect 20622 19932 20628 19984
rect 20680 19932 20686 19984
rect 15473 19907 15531 19913
rect 15473 19904 15485 19907
rect 15252 19876 15485 19904
rect 15252 19864 15258 19876
rect 15473 19873 15485 19876
rect 15519 19873 15531 19907
rect 15473 19867 15531 19873
rect 15749 19907 15807 19913
rect 15749 19873 15761 19907
rect 15795 19904 15807 19907
rect 15930 19904 15936 19916
rect 15795 19876 15936 19904
rect 15795 19873 15807 19876
rect 15749 19867 15807 19873
rect 15930 19864 15936 19876
rect 15988 19864 15994 19916
rect 16114 19904 16120 19916
rect 16075 19876 16120 19904
rect 16114 19864 16120 19876
rect 16172 19864 16178 19916
rect 16209 19907 16267 19913
rect 16209 19873 16221 19907
rect 16255 19873 16267 19907
rect 16390 19904 16396 19916
rect 16351 19876 16396 19904
rect 16209 19867 16267 19873
rect 14550 19836 14556 19848
rect 8128 19808 8432 19836
rect 14511 19808 14556 19836
rect 5353 19799 5411 19805
rect 5040 19740 5120 19768
rect 5040 19728 5046 19740
rect 5258 19728 5264 19780
rect 5316 19768 5322 19780
rect 5368 19768 5396 19799
rect 14550 19796 14556 19808
rect 14608 19796 14614 19848
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19805 14703 19839
rect 14645 19799 14703 19805
rect 8846 19768 8852 19780
rect 5316 19740 8852 19768
rect 5316 19728 5322 19740
rect 8846 19728 8852 19740
rect 8904 19728 8910 19780
rect 14660 19768 14688 19799
rect 14918 19796 14924 19848
rect 14976 19836 14982 19848
rect 15013 19839 15071 19845
rect 15013 19836 15025 19839
rect 14976 19808 15025 19836
rect 14976 19796 14982 19808
rect 15013 19805 15025 19808
rect 15059 19805 15071 19839
rect 16224 19836 16252 19867
rect 16390 19864 16396 19876
rect 16448 19864 16454 19916
rect 17770 19864 17776 19916
rect 17828 19904 17834 19916
rect 19613 19907 19671 19913
rect 19613 19904 19625 19907
rect 17828 19876 19625 19904
rect 17828 19864 17834 19876
rect 19613 19873 19625 19876
rect 19659 19873 19671 19907
rect 19613 19867 19671 19873
rect 15013 19799 15071 19805
rect 15856 19808 16252 19836
rect 19889 19839 19947 19845
rect 14660 19740 15240 19768
rect 15212 19712 15240 19740
rect 5718 19660 5724 19712
rect 5776 19700 5782 19712
rect 5997 19703 6055 19709
rect 5997 19700 6009 19703
rect 5776 19672 6009 19700
rect 5776 19660 5782 19672
rect 5997 19669 6009 19672
rect 6043 19669 6055 19703
rect 5997 19663 6055 19669
rect 14369 19703 14427 19709
rect 14369 19669 14381 19703
rect 14415 19700 14427 19703
rect 14642 19700 14648 19712
rect 14415 19672 14648 19700
rect 14415 19669 14427 19672
rect 14369 19663 14427 19669
rect 14642 19660 14648 19672
rect 14700 19660 14706 19712
rect 15194 19660 15200 19712
rect 15252 19700 15258 19712
rect 15657 19703 15715 19709
rect 15657 19700 15669 19703
rect 15252 19672 15669 19700
rect 15252 19660 15258 19672
rect 15657 19669 15669 19672
rect 15703 19669 15715 19703
rect 15657 19663 15715 19669
rect 15746 19660 15752 19712
rect 15804 19700 15810 19712
rect 15856 19709 15884 19808
rect 19889 19805 19901 19839
rect 19935 19836 19947 19839
rect 20898 19836 20904 19848
rect 19935 19808 20904 19836
rect 19935 19805 19947 19808
rect 19889 19799 19947 19805
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 16393 19771 16451 19777
rect 16393 19737 16405 19771
rect 16439 19768 16451 19771
rect 16482 19768 16488 19780
rect 16439 19740 16488 19768
rect 16439 19737 16451 19740
rect 16393 19731 16451 19737
rect 16482 19728 16488 19740
rect 16540 19728 16546 19780
rect 15841 19703 15899 19709
rect 15841 19700 15853 19703
rect 15804 19672 15853 19700
rect 15804 19660 15810 19672
rect 15841 19669 15853 19672
rect 15887 19669 15899 19703
rect 15841 19663 15899 19669
rect 1104 19610 21804 19632
rect 1104 19558 4432 19610
rect 4484 19558 4496 19610
rect 4548 19558 4560 19610
rect 4612 19558 4624 19610
rect 4676 19558 11332 19610
rect 11384 19558 11396 19610
rect 11448 19558 11460 19610
rect 11512 19558 11524 19610
rect 11576 19558 18232 19610
rect 18284 19558 18296 19610
rect 18348 19558 18360 19610
rect 18412 19558 18424 19610
rect 18476 19558 21804 19610
rect 1104 19536 21804 19558
rect 5169 19499 5227 19505
rect 5169 19465 5181 19499
rect 5215 19496 5227 19499
rect 5442 19496 5448 19508
rect 5215 19468 5448 19496
rect 5215 19465 5227 19468
rect 5169 19459 5227 19465
rect 5442 19456 5448 19468
rect 5500 19456 5506 19508
rect 5629 19499 5687 19505
rect 5629 19465 5641 19499
rect 5675 19496 5687 19499
rect 5675 19468 6040 19496
rect 5675 19465 5687 19468
rect 5629 19459 5687 19465
rect 4890 19388 4896 19440
rect 4948 19428 4954 19440
rect 5350 19428 5356 19440
rect 4948 19400 5356 19428
rect 4948 19388 4954 19400
rect 5350 19388 5356 19400
rect 5408 19428 5414 19440
rect 6012 19437 6040 19468
rect 7742 19456 7748 19508
rect 7800 19496 7806 19508
rect 7929 19499 7987 19505
rect 7929 19496 7941 19499
rect 7800 19468 7941 19496
rect 7800 19456 7806 19468
rect 7929 19465 7941 19468
rect 7975 19465 7987 19499
rect 7929 19459 7987 19465
rect 14550 19456 14556 19508
rect 14608 19496 14614 19508
rect 15010 19496 15016 19508
rect 14608 19468 15016 19496
rect 14608 19456 14614 19468
rect 15010 19456 15016 19468
rect 15068 19456 15074 19508
rect 20622 19496 20628 19508
rect 20583 19468 20628 19496
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 5997 19431 6055 19437
rect 5408 19400 5856 19428
rect 5408 19388 5414 19400
rect 5828 19369 5856 19400
rect 5997 19397 6009 19431
rect 6043 19428 6055 19431
rect 6454 19428 6460 19440
rect 6043 19400 6460 19428
rect 6043 19397 6055 19400
rect 5997 19391 6055 19397
rect 6454 19388 6460 19400
rect 6512 19388 6518 19440
rect 7392 19400 8248 19428
rect 5813 19363 5871 19369
rect 5813 19329 5825 19363
rect 5859 19329 5871 19363
rect 5813 19323 5871 19329
rect 5166 19252 5172 19304
rect 5224 19292 5230 19304
rect 5353 19295 5411 19301
rect 5353 19292 5365 19295
rect 5224 19264 5365 19292
rect 5224 19252 5230 19264
rect 5353 19261 5365 19264
rect 5399 19261 5411 19295
rect 5353 19255 5411 19261
rect 5445 19295 5503 19301
rect 5445 19261 5457 19295
rect 5491 19292 5503 19295
rect 5626 19292 5632 19304
rect 5491 19264 5632 19292
rect 5491 19261 5503 19264
rect 5445 19255 5503 19261
rect 5626 19252 5632 19264
rect 5684 19252 5690 19304
rect 5718 19252 5724 19304
rect 5776 19292 5782 19304
rect 6089 19295 6147 19301
rect 5776 19264 5821 19292
rect 5776 19252 5782 19264
rect 6089 19261 6101 19295
rect 6135 19261 6147 19295
rect 6089 19255 6147 19261
rect 5736 19224 5764 19252
rect 6104 19224 6132 19255
rect 6454 19252 6460 19304
rect 6512 19292 6518 19304
rect 7392 19301 7420 19400
rect 7466 19320 7472 19372
rect 7524 19360 7530 19372
rect 8220 19369 8248 19400
rect 8021 19363 8079 19369
rect 8021 19360 8033 19363
rect 7524 19332 8033 19360
rect 7524 19320 7530 19332
rect 8021 19329 8033 19332
rect 8067 19329 8079 19363
rect 8021 19323 8079 19329
rect 8205 19363 8263 19369
rect 8205 19329 8217 19363
rect 8251 19360 8263 19363
rect 8754 19360 8760 19372
rect 8251 19332 8760 19360
rect 8251 19329 8263 19332
rect 8205 19323 8263 19329
rect 8754 19320 8760 19332
rect 8812 19320 8818 19372
rect 14642 19360 14648 19372
rect 14016 19332 14648 19360
rect 7377 19295 7435 19301
rect 7377 19292 7389 19295
rect 6512 19264 7389 19292
rect 6512 19252 6518 19264
rect 7377 19261 7389 19264
rect 7423 19261 7435 19295
rect 7558 19292 7564 19304
rect 7519 19264 7564 19292
rect 7377 19255 7435 19261
rect 7558 19252 7564 19264
rect 7616 19252 7622 19304
rect 7745 19295 7803 19301
rect 7745 19261 7757 19295
rect 7791 19261 7803 19295
rect 8294 19292 8300 19304
rect 8255 19264 8300 19292
rect 7745 19255 7803 19261
rect 7650 19224 7656 19236
rect 5736 19196 6132 19224
rect 7611 19196 7656 19224
rect 7650 19184 7656 19196
rect 7708 19184 7714 19236
rect 5810 19156 5816 19168
rect 5771 19128 5816 19156
rect 5810 19116 5816 19128
rect 5868 19116 5874 19168
rect 7558 19116 7564 19168
rect 7616 19156 7622 19168
rect 7760 19156 7788 19255
rect 8294 19252 8300 19264
rect 8352 19252 8358 19304
rect 8573 19295 8631 19301
rect 8573 19261 8585 19295
rect 8619 19292 8631 19295
rect 9582 19292 9588 19304
rect 8619 19264 9588 19292
rect 8619 19261 8631 19264
rect 8573 19255 8631 19261
rect 8021 19227 8079 19233
rect 8021 19193 8033 19227
rect 8067 19224 8079 19227
rect 8588 19224 8616 19255
rect 9582 19252 9588 19264
rect 9640 19252 9646 19304
rect 12710 19292 12716 19304
rect 12623 19264 12716 19292
rect 12710 19252 12716 19264
rect 12768 19292 12774 19304
rect 13817 19295 13875 19301
rect 12768 19264 13216 19292
rect 12768 19252 12774 19264
rect 8067 19196 8616 19224
rect 13188 19224 13216 19264
rect 13817 19261 13829 19295
rect 13863 19292 13875 19295
rect 13906 19292 13912 19304
rect 13863 19264 13912 19292
rect 13863 19261 13875 19264
rect 13817 19255 13875 19261
rect 13906 19252 13912 19264
rect 13964 19252 13970 19304
rect 14016 19301 14044 19332
rect 14642 19320 14648 19332
rect 14700 19320 14706 19372
rect 14001 19295 14059 19301
rect 14001 19261 14013 19295
rect 14047 19261 14059 19295
rect 14001 19255 14059 19261
rect 14369 19295 14427 19301
rect 14369 19261 14381 19295
rect 14415 19261 14427 19295
rect 14369 19255 14427 19261
rect 14185 19227 14243 19233
rect 14185 19224 14197 19227
rect 13188 19196 14197 19224
rect 8067 19193 8079 19196
rect 8021 19187 8079 19193
rect 14185 19193 14197 19196
rect 14231 19193 14243 19227
rect 14384 19224 14412 19255
rect 14458 19252 14464 19304
rect 14516 19292 14522 19304
rect 14553 19295 14611 19301
rect 14553 19292 14565 19295
rect 14516 19264 14565 19292
rect 14516 19252 14522 19264
rect 14553 19261 14565 19264
rect 14599 19261 14611 19295
rect 14734 19292 14740 19304
rect 14695 19264 14740 19292
rect 14553 19255 14611 19261
rect 14734 19252 14740 19264
rect 14792 19252 14798 19304
rect 14918 19292 14924 19304
rect 14879 19264 14924 19292
rect 14918 19252 14924 19264
rect 14976 19292 14982 19304
rect 15381 19295 15439 19301
rect 15381 19292 15393 19295
rect 14976 19264 15393 19292
rect 14976 19252 14982 19264
rect 15381 19261 15393 19264
rect 15427 19261 15439 19295
rect 15381 19255 15439 19261
rect 17126 19252 17132 19304
rect 17184 19292 17190 19304
rect 17589 19295 17647 19301
rect 17589 19292 17601 19295
rect 17184 19264 17601 19292
rect 17184 19252 17190 19264
rect 17589 19261 17601 19264
rect 17635 19292 17647 19295
rect 20438 19292 20444 19304
rect 17635 19264 20444 19292
rect 17635 19261 17647 19264
rect 17589 19255 17647 19261
rect 20438 19252 20444 19264
rect 20496 19252 20502 19304
rect 14384 19196 14964 19224
rect 14185 19187 14243 19193
rect 7616 19128 7788 19156
rect 8665 19159 8723 19165
rect 7616 19116 7622 19128
rect 8665 19125 8677 19159
rect 8711 19156 8723 19159
rect 9214 19156 9220 19168
rect 8711 19128 9220 19156
rect 8711 19125 8723 19128
rect 8665 19119 8723 19125
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 12618 19156 12624 19168
rect 12579 19128 12624 19156
rect 12618 19116 12624 19128
rect 12676 19116 12682 19168
rect 12986 19116 12992 19168
rect 13044 19156 13050 19168
rect 13817 19159 13875 19165
rect 13817 19156 13829 19159
rect 13044 19128 13829 19156
rect 13044 19116 13050 19128
rect 13817 19125 13829 19128
rect 13863 19125 13875 19159
rect 13817 19119 13875 19125
rect 13906 19116 13912 19168
rect 13964 19156 13970 19168
rect 14642 19156 14648 19168
rect 13964 19128 14648 19156
rect 13964 19116 13970 19128
rect 14642 19116 14648 19128
rect 14700 19116 14706 19168
rect 14936 19156 14964 19196
rect 15010 19184 15016 19236
rect 15068 19224 15074 19236
rect 15194 19224 15200 19236
rect 15068 19196 15113 19224
rect 15155 19196 15200 19224
rect 15068 19184 15074 19196
rect 15194 19184 15200 19196
rect 15252 19184 15258 19236
rect 15746 19156 15752 19168
rect 14936 19128 15752 19156
rect 15746 19116 15752 19128
rect 15804 19116 15810 19168
rect 17678 19116 17684 19168
rect 17736 19156 17742 19168
rect 17773 19159 17831 19165
rect 17773 19156 17785 19159
rect 17736 19128 17785 19156
rect 17736 19116 17742 19128
rect 17773 19125 17785 19128
rect 17819 19125 17831 19159
rect 17773 19119 17831 19125
rect 1104 19066 21804 19088
rect 1104 19014 7882 19066
rect 7934 19014 7946 19066
rect 7998 19014 8010 19066
rect 8062 19014 8074 19066
rect 8126 19014 14782 19066
rect 14834 19014 14846 19066
rect 14898 19014 14910 19066
rect 14962 19014 14974 19066
rect 15026 19014 21804 19066
rect 1104 18992 21804 19014
rect 19061 18955 19119 18961
rect 19061 18952 19073 18955
rect 15580 18924 19073 18952
rect 8757 18887 8815 18893
rect 8757 18853 8769 18887
rect 8803 18884 8815 18887
rect 9493 18887 9551 18893
rect 9493 18884 9505 18887
rect 8803 18856 9505 18884
rect 8803 18853 8815 18856
rect 8757 18847 8815 18853
rect 9493 18853 9505 18856
rect 9539 18853 9551 18887
rect 12986 18884 12992 18896
rect 12947 18856 12992 18884
rect 9493 18847 9551 18853
rect 12986 18844 12992 18856
rect 13044 18844 13050 18896
rect 15580 18884 15608 18924
rect 19061 18921 19073 18924
rect 19107 18921 19119 18955
rect 19061 18915 19119 18921
rect 13280 18856 15608 18884
rect 16577 18887 16635 18893
rect 6454 18776 6460 18828
rect 6512 18816 6518 18828
rect 6549 18819 6607 18825
rect 6549 18816 6561 18819
rect 6512 18788 6561 18816
rect 6512 18776 6518 18788
rect 6549 18785 6561 18788
rect 6595 18785 6607 18819
rect 6549 18779 6607 18785
rect 8665 18819 8723 18825
rect 8665 18785 8677 18819
rect 8711 18785 8723 18819
rect 8665 18779 8723 18785
rect 8478 18708 8484 18760
rect 8536 18748 8542 18760
rect 8680 18748 8708 18779
rect 8846 18776 8852 18828
rect 8904 18816 8910 18828
rect 9125 18819 9183 18825
rect 9125 18816 9137 18819
rect 8904 18788 9137 18816
rect 8904 18776 8910 18788
rect 9125 18785 9137 18788
rect 9171 18785 9183 18819
rect 9125 18779 9183 18785
rect 9214 18776 9220 18828
rect 9272 18816 9278 18828
rect 9401 18819 9459 18825
rect 9272 18788 9317 18816
rect 9272 18776 9278 18788
rect 9401 18785 9413 18819
rect 9447 18785 9459 18819
rect 9582 18816 9588 18828
rect 9640 18825 9646 18828
rect 9548 18788 9588 18816
rect 9401 18779 9459 18785
rect 9416 18748 9444 18779
rect 9582 18776 9588 18788
rect 9640 18779 9648 18825
rect 12526 18816 12532 18828
rect 12487 18788 12532 18816
rect 9640 18776 9646 18779
rect 12526 18776 12532 18788
rect 12584 18776 12590 18828
rect 12621 18819 12679 18825
rect 12621 18785 12633 18819
rect 12667 18816 12679 18819
rect 12710 18816 12716 18828
rect 12667 18788 12716 18816
rect 12667 18785 12679 18788
rect 12621 18779 12679 18785
rect 12710 18776 12716 18788
rect 12768 18776 12774 18828
rect 12897 18819 12955 18825
rect 12897 18785 12909 18819
rect 12943 18816 12955 18819
rect 13280 18816 13308 18856
rect 16577 18853 16589 18887
rect 16623 18884 16635 18887
rect 16945 18887 17003 18893
rect 16945 18884 16957 18887
rect 16623 18856 16957 18884
rect 16623 18853 16635 18856
rect 16577 18847 16635 18853
rect 16945 18853 16957 18856
rect 16991 18853 17003 18887
rect 16945 18847 17003 18853
rect 17678 18844 17684 18896
rect 17736 18844 17742 18896
rect 12943 18788 13308 18816
rect 12943 18785 12955 18788
rect 12897 18779 12955 18785
rect 13354 18776 13360 18828
rect 13412 18816 13418 18828
rect 15838 18816 15844 18828
rect 13412 18788 13457 18816
rect 15799 18788 15844 18816
rect 13412 18776 13418 18788
rect 15838 18776 15844 18788
rect 15896 18776 15902 18828
rect 16022 18816 16028 18828
rect 15983 18788 16028 18816
rect 16022 18776 16028 18788
rect 16080 18776 16086 18828
rect 16114 18776 16120 18828
rect 16172 18816 16178 18828
rect 16393 18819 16451 18825
rect 16172 18788 16217 18816
rect 16172 18776 16178 18788
rect 16393 18785 16405 18819
rect 16439 18816 16451 18819
rect 16482 18816 16488 18828
rect 16439 18788 16488 18816
rect 16439 18785 16451 18788
rect 16393 18779 16451 18785
rect 16482 18776 16488 18788
rect 16540 18776 16546 18828
rect 19150 18816 19156 18828
rect 19111 18788 19156 18816
rect 19150 18776 19156 18788
rect 19208 18776 19214 18828
rect 19245 18819 19303 18825
rect 19245 18785 19257 18819
rect 19291 18785 19303 18819
rect 19245 18779 19303 18785
rect 12802 18748 12808 18760
rect 8536 18720 9444 18748
rect 12763 18720 12808 18748
rect 8536 18708 8542 18720
rect 12802 18708 12808 18720
rect 12860 18748 12866 18760
rect 13081 18751 13139 18757
rect 13081 18748 13093 18751
rect 12860 18720 13093 18748
rect 12860 18708 12866 18720
rect 13081 18717 13093 18720
rect 13127 18717 13139 18751
rect 16206 18748 16212 18760
rect 16167 18720 16212 18748
rect 13081 18711 13139 18717
rect 16206 18708 16212 18720
rect 16264 18708 16270 18760
rect 16669 18751 16727 18757
rect 16669 18717 16681 18751
rect 16715 18748 16727 18751
rect 17678 18748 17684 18760
rect 16715 18720 17684 18748
rect 16715 18717 16727 18720
rect 16669 18711 16727 18717
rect 17678 18708 17684 18720
rect 17736 18708 17742 18760
rect 18414 18748 18420 18760
rect 18375 18720 18420 18748
rect 18414 18708 18420 18720
rect 18472 18708 18478 18760
rect 18782 18748 18788 18760
rect 18743 18720 18788 18748
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 19058 18708 19064 18760
rect 19116 18748 19122 18760
rect 19260 18748 19288 18779
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 19610 18816 19616 18828
rect 19392 18788 19616 18816
rect 19392 18776 19398 18788
rect 19610 18776 19616 18788
rect 19668 18776 19674 18828
rect 19797 18819 19855 18825
rect 19797 18785 19809 18819
rect 19843 18785 19855 18819
rect 19797 18779 19855 18785
rect 19116 18720 19288 18748
rect 19116 18708 19122 18720
rect 19426 18708 19432 18760
rect 19484 18748 19490 18760
rect 19812 18748 19840 18779
rect 19484 18720 19840 18748
rect 19484 18708 19490 18720
rect 8846 18640 8852 18692
rect 8904 18680 8910 18692
rect 12345 18683 12403 18689
rect 12345 18680 12357 18683
rect 8904 18652 12357 18680
rect 8904 18640 8910 18652
rect 12345 18649 12357 18652
rect 12391 18649 12403 18683
rect 12345 18643 12403 18649
rect 5626 18572 5632 18624
rect 5684 18612 5690 18624
rect 6641 18615 6699 18621
rect 6641 18612 6653 18615
rect 5684 18584 6653 18612
rect 5684 18572 5690 18584
rect 6641 18581 6653 18584
rect 6687 18612 6699 18615
rect 7558 18612 7564 18624
rect 6687 18584 7564 18612
rect 6687 18581 6699 18584
rect 6641 18575 6699 18581
rect 7558 18572 7564 18584
rect 7616 18612 7622 18624
rect 8938 18612 8944 18624
rect 7616 18584 8944 18612
rect 7616 18572 7622 18584
rect 8938 18572 8944 18584
rect 8996 18572 9002 18624
rect 9398 18572 9404 18624
rect 9456 18612 9462 18624
rect 9769 18615 9827 18621
rect 9769 18612 9781 18615
rect 9456 18584 9781 18612
rect 9456 18572 9462 18584
rect 9769 18581 9781 18584
rect 9815 18581 9827 18615
rect 13170 18612 13176 18624
rect 13131 18584 13176 18612
rect 9769 18575 9827 18581
rect 13170 18572 13176 18584
rect 13228 18572 13234 18624
rect 13265 18615 13323 18621
rect 13265 18581 13277 18615
rect 13311 18612 13323 18615
rect 16482 18612 16488 18624
rect 13311 18584 16488 18612
rect 13311 18581 13323 18584
rect 13265 18575 13323 18581
rect 16482 18572 16488 18584
rect 16540 18572 16546 18624
rect 19705 18615 19763 18621
rect 19705 18581 19717 18615
rect 19751 18612 19763 18615
rect 19794 18612 19800 18624
rect 19751 18584 19800 18612
rect 19751 18581 19763 18584
rect 19705 18575 19763 18581
rect 19794 18572 19800 18584
rect 19852 18572 19858 18624
rect 1104 18522 21804 18544
rect 1104 18470 4432 18522
rect 4484 18470 4496 18522
rect 4548 18470 4560 18522
rect 4612 18470 4624 18522
rect 4676 18470 11332 18522
rect 11384 18470 11396 18522
rect 11448 18470 11460 18522
rect 11512 18470 11524 18522
rect 11576 18470 18232 18522
rect 18284 18470 18296 18522
rect 18348 18470 18360 18522
rect 18412 18470 18424 18522
rect 18476 18470 21804 18522
rect 1104 18448 21804 18470
rect 8478 18408 8484 18420
rect 8439 18380 8484 18408
rect 8478 18368 8484 18380
rect 8536 18368 8542 18420
rect 8938 18408 8944 18420
rect 8899 18380 8944 18408
rect 8938 18368 8944 18380
rect 8996 18368 9002 18420
rect 16114 18368 16120 18420
rect 16172 18408 16178 18420
rect 16669 18411 16727 18417
rect 16669 18408 16681 18411
rect 16172 18380 16681 18408
rect 16172 18368 16178 18380
rect 16669 18377 16681 18380
rect 16715 18377 16727 18411
rect 16669 18371 16727 18377
rect 12986 18300 12992 18352
rect 13044 18300 13050 18352
rect 13354 18300 13360 18352
rect 13412 18340 13418 18352
rect 18693 18343 18751 18349
rect 18693 18340 18705 18343
rect 13412 18312 18705 18340
rect 13412 18300 13418 18312
rect 18693 18309 18705 18312
rect 18739 18309 18751 18343
rect 18693 18303 18751 18309
rect 19150 18300 19156 18352
rect 19208 18340 19214 18352
rect 19208 18312 19656 18340
rect 19208 18300 19214 18312
rect 2498 18232 2504 18284
rect 2556 18272 2562 18284
rect 2685 18275 2743 18281
rect 2685 18272 2697 18275
rect 2556 18244 2697 18272
rect 2556 18232 2562 18244
rect 2685 18241 2697 18244
rect 2731 18241 2743 18275
rect 2685 18235 2743 18241
rect 2961 18275 3019 18281
rect 2961 18241 2973 18275
rect 3007 18272 3019 18275
rect 4614 18272 4620 18284
rect 3007 18244 4620 18272
rect 3007 18241 3019 18244
rect 2961 18235 3019 18241
rect 4614 18232 4620 18244
rect 4672 18232 4678 18284
rect 9398 18272 9404 18284
rect 9359 18244 9404 18272
rect 9398 18232 9404 18244
rect 9456 18232 9462 18284
rect 13004 18272 13032 18300
rect 12820 18244 13032 18272
rect 8665 18207 8723 18213
rect 8665 18173 8677 18207
rect 8711 18173 8723 18207
rect 8787 18207 8845 18213
rect 8787 18204 8799 18207
rect 8665 18167 8723 18173
rect 8772 18173 8799 18204
rect 8833 18173 8845 18207
rect 8772 18167 8845 18173
rect 9033 18207 9091 18213
rect 9033 18173 9045 18207
rect 9079 18204 9091 18207
rect 9122 18204 9128 18216
rect 9079 18176 9128 18204
rect 9079 18173 9091 18176
rect 9033 18167 9091 18173
rect 3970 18096 3976 18148
rect 4028 18096 4034 18148
rect 8680 18136 8708 18167
rect 8589 18108 8708 18136
rect 8772 18136 8800 18167
rect 9122 18164 9128 18176
rect 9180 18164 9186 18216
rect 9217 18207 9275 18213
rect 9217 18173 9229 18207
rect 9263 18204 9275 18207
rect 9306 18204 9312 18216
rect 9263 18176 9312 18204
rect 9263 18173 9275 18176
rect 9217 18167 9275 18173
rect 9306 18164 9312 18176
rect 9364 18164 9370 18216
rect 10318 18204 10324 18216
rect 10231 18176 10324 18204
rect 10318 18164 10324 18176
rect 10376 18204 10382 18216
rect 10962 18204 10968 18216
rect 10376 18176 10968 18204
rect 10376 18164 10382 18176
rect 10962 18164 10968 18176
rect 11020 18164 11026 18216
rect 12618 18204 12624 18216
rect 12579 18176 12624 18204
rect 12618 18164 12624 18176
rect 12676 18164 12682 18216
rect 12820 18213 12848 18244
rect 13170 18232 13176 18284
rect 13228 18272 13234 18284
rect 13228 18244 13492 18272
rect 13228 18232 13234 18244
rect 12805 18207 12863 18213
rect 12805 18173 12817 18207
rect 12851 18173 12863 18207
rect 12986 18204 12992 18216
rect 12947 18176 12992 18204
rect 12805 18167 12863 18173
rect 12986 18164 12992 18176
rect 13044 18164 13050 18216
rect 13262 18204 13268 18216
rect 13223 18176 13268 18204
rect 13262 18164 13268 18176
rect 13320 18164 13326 18216
rect 13464 18213 13492 18244
rect 19058 18232 19064 18284
rect 19116 18272 19122 18284
rect 19521 18275 19579 18281
rect 19521 18272 19533 18275
rect 19116 18244 19533 18272
rect 19116 18232 19122 18244
rect 19521 18241 19533 18244
rect 19567 18241 19579 18275
rect 19521 18235 19579 18241
rect 19628 18272 19656 18312
rect 21266 18272 21272 18284
rect 19628 18244 21272 18272
rect 13449 18207 13507 18213
rect 13449 18173 13461 18207
rect 13495 18173 13507 18207
rect 16574 18204 16580 18216
rect 16535 18176 16580 18204
rect 13449 18167 13507 18173
rect 16574 18164 16580 18176
rect 16632 18164 16638 18216
rect 16761 18207 16819 18213
rect 16761 18173 16773 18207
rect 16807 18173 16819 18207
rect 16761 18167 16819 18173
rect 18785 18207 18843 18213
rect 18785 18173 18797 18207
rect 18831 18173 18843 18207
rect 18785 18167 18843 18173
rect 19245 18207 19303 18213
rect 19245 18173 19257 18207
rect 19291 18204 19303 18207
rect 19334 18204 19340 18216
rect 19291 18176 19340 18204
rect 19291 18173 19303 18176
rect 19245 18167 19303 18173
rect 12161 18139 12219 18145
rect 12161 18136 12173 18139
rect 8772 18108 12173 18136
rect 4433 18071 4491 18077
rect 4433 18037 4445 18071
rect 4479 18068 4491 18071
rect 5166 18068 5172 18080
rect 4479 18040 5172 18068
rect 4479 18037 4491 18040
rect 4433 18031 4491 18037
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 8589 18068 8617 18108
rect 8772 18080 8800 18108
rect 12161 18105 12173 18108
rect 12207 18105 12219 18139
rect 12161 18099 12219 18105
rect 16206 18096 16212 18148
rect 16264 18136 16270 18148
rect 16776 18136 16804 18167
rect 16850 18136 16856 18148
rect 16264 18108 16856 18136
rect 16264 18096 16270 18108
rect 16850 18096 16856 18108
rect 16908 18096 16914 18148
rect 18800 18136 18828 18167
rect 19334 18164 19340 18176
rect 19392 18164 19398 18216
rect 19426 18164 19432 18216
rect 19484 18204 19490 18216
rect 19628 18213 19656 18244
rect 21266 18232 21272 18244
rect 21324 18232 21330 18284
rect 19613 18207 19671 18213
rect 19484 18176 19529 18204
rect 19484 18164 19490 18176
rect 19613 18173 19625 18207
rect 19659 18173 19671 18207
rect 19794 18204 19800 18216
rect 19755 18176 19800 18204
rect 19613 18167 19671 18173
rect 19794 18164 19800 18176
rect 19852 18164 19858 18216
rect 19812 18136 19840 18164
rect 18800 18108 19840 18136
rect 8662 18068 8668 18080
rect 8589 18040 8668 18068
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 8754 18028 8760 18080
rect 8812 18028 8818 18080
rect 9401 18071 9459 18077
rect 9401 18037 9413 18071
rect 9447 18068 9459 18071
rect 9582 18068 9588 18080
rect 9447 18040 9588 18068
rect 9447 18037 9459 18040
rect 9401 18031 9459 18037
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 10505 18071 10563 18077
rect 10505 18037 10517 18071
rect 10551 18068 10563 18071
rect 10594 18068 10600 18080
rect 10551 18040 10600 18068
rect 10551 18037 10563 18040
rect 10505 18031 10563 18037
rect 10594 18028 10600 18040
rect 10652 18028 10658 18080
rect 16482 18028 16488 18080
rect 16540 18068 16546 18080
rect 18782 18068 18788 18080
rect 16540 18040 18788 18068
rect 16540 18028 16546 18040
rect 18782 18028 18788 18040
rect 18840 18068 18846 18080
rect 19061 18071 19119 18077
rect 19061 18068 19073 18071
rect 18840 18040 19073 18068
rect 18840 18028 18846 18040
rect 19061 18037 19073 18040
rect 19107 18037 19119 18071
rect 19061 18031 19119 18037
rect 1104 17978 21804 18000
rect 1104 17926 7882 17978
rect 7934 17926 7946 17978
rect 7998 17926 8010 17978
rect 8062 17926 8074 17978
rect 8126 17926 14782 17978
rect 14834 17926 14846 17978
rect 14898 17926 14910 17978
rect 14962 17926 14974 17978
rect 15026 17926 21804 17978
rect 1104 17904 21804 17926
rect 3881 17867 3939 17873
rect 3881 17833 3893 17867
rect 3927 17864 3939 17867
rect 3970 17864 3976 17876
rect 3927 17836 3976 17864
rect 3927 17833 3939 17836
rect 3881 17827 3939 17833
rect 3970 17824 3976 17836
rect 4028 17824 4034 17876
rect 4614 17864 4620 17876
rect 4575 17836 4620 17864
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 5994 17864 6000 17876
rect 4908 17836 6000 17864
rect 4908 17805 4936 17836
rect 5994 17824 6000 17836
rect 6052 17824 6058 17876
rect 15838 17864 15844 17876
rect 14752 17836 15844 17864
rect 4893 17799 4951 17805
rect 4893 17765 4905 17799
rect 4939 17765 4951 17799
rect 4893 17759 4951 17765
rect 4982 17756 4988 17808
rect 5040 17796 5046 17808
rect 5537 17799 5595 17805
rect 5040 17768 5488 17796
rect 5040 17756 5046 17768
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 3694 17688 3700 17740
rect 3752 17728 3758 17740
rect 5166 17737 5172 17740
rect 4065 17731 4123 17737
rect 4065 17728 4077 17731
rect 3752 17700 4077 17728
rect 3752 17688 3758 17700
rect 4065 17697 4077 17700
rect 4111 17697 4123 17731
rect 4065 17691 4123 17697
rect 4801 17731 4859 17737
rect 4801 17697 4813 17731
rect 4847 17697 4859 17731
rect 4801 17691 4859 17697
rect 5123 17731 5172 17737
rect 5123 17697 5135 17731
rect 5169 17697 5172 17731
rect 5123 17691 5172 17697
rect 1578 17524 1584 17536
rect 1539 17496 1584 17524
rect 1578 17484 1584 17496
rect 1636 17484 1642 17536
rect 4816 17524 4844 17691
rect 5166 17688 5172 17691
rect 5224 17688 5230 17740
rect 5258 17688 5264 17740
rect 5316 17728 5322 17740
rect 5460 17728 5488 17768
rect 5537 17765 5549 17799
rect 5583 17796 5595 17799
rect 5810 17796 5816 17808
rect 5583 17768 5816 17796
rect 5583 17765 5595 17768
rect 5537 17759 5595 17765
rect 5810 17756 5816 17768
rect 5868 17796 5874 17808
rect 9582 17796 9588 17808
rect 5868 17768 6500 17796
rect 9543 17768 9588 17796
rect 5868 17756 5874 17768
rect 5718 17728 5724 17740
rect 5316 17700 5361 17728
rect 5460 17700 5580 17728
rect 5679 17700 5724 17728
rect 5316 17688 5322 17700
rect 5552 17592 5580 17700
rect 5718 17688 5724 17700
rect 5776 17688 5782 17740
rect 6181 17731 6239 17737
rect 6181 17697 6193 17731
rect 6227 17697 6239 17731
rect 6181 17691 6239 17697
rect 6196 17660 6224 17691
rect 6270 17688 6276 17740
rect 6328 17728 6334 17740
rect 6472 17737 6500 17768
rect 9582 17756 9588 17768
rect 9640 17756 9646 17808
rect 10594 17756 10600 17808
rect 10652 17756 10658 17808
rect 6365 17731 6423 17737
rect 6365 17728 6377 17731
rect 6328 17700 6377 17728
rect 6328 17688 6334 17700
rect 6365 17697 6377 17700
rect 6411 17697 6423 17731
rect 6365 17691 6423 17697
rect 6457 17731 6515 17737
rect 6457 17697 6469 17731
rect 6503 17697 6515 17731
rect 6457 17691 6515 17697
rect 7742 17688 7748 17740
rect 7800 17728 7806 17740
rect 8021 17731 8079 17737
rect 8021 17728 8033 17731
rect 7800 17700 8033 17728
rect 7800 17688 7806 17700
rect 8021 17697 8033 17700
rect 8067 17697 8079 17731
rect 8021 17691 8079 17697
rect 8481 17731 8539 17737
rect 8481 17697 8493 17731
rect 8527 17728 8539 17731
rect 8754 17728 8760 17740
rect 8527 17700 8760 17728
rect 8527 17697 8539 17700
rect 8481 17691 8539 17697
rect 8754 17688 8760 17700
rect 8812 17688 8818 17740
rect 9030 17688 9036 17740
rect 9088 17728 9094 17740
rect 9309 17731 9367 17737
rect 9309 17728 9321 17731
rect 9088 17700 9321 17728
rect 9088 17688 9094 17700
rect 9309 17697 9321 17700
rect 9355 17697 9367 17731
rect 9309 17691 9367 17697
rect 11790 17688 11796 17740
rect 11848 17728 11854 17740
rect 12161 17731 12219 17737
rect 12161 17728 12173 17731
rect 11848 17700 12173 17728
rect 11848 17688 11854 17700
rect 12161 17697 12173 17700
rect 12207 17728 12219 17731
rect 12342 17728 12348 17740
rect 12207 17700 12348 17728
rect 12207 17697 12219 17700
rect 12161 17691 12219 17697
rect 12342 17688 12348 17700
rect 12400 17688 12406 17740
rect 12434 17688 12440 17740
rect 12492 17728 12498 17740
rect 12529 17731 12587 17737
rect 12529 17728 12541 17731
rect 12492 17700 12541 17728
rect 12492 17688 12498 17700
rect 12529 17697 12541 17700
rect 12575 17697 12587 17731
rect 12529 17691 12587 17697
rect 13906 17688 13912 17740
rect 13964 17728 13970 17740
rect 14752 17737 14780 17836
rect 15838 17824 15844 17836
rect 15896 17864 15902 17876
rect 17310 17864 17316 17876
rect 15896 17836 17316 17864
rect 15896 17824 15902 17836
rect 17310 17824 17316 17836
rect 17368 17824 17374 17876
rect 14829 17799 14887 17805
rect 14829 17765 14841 17799
rect 14875 17796 14887 17799
rect 16206 17796 16212 17808
rect 14875 17768 16212 17796
rect 14875 17765 14887 17768
rect 14829 17759 14887 17765
rect 16206 17756 16212 17768
rect 16264 17756 16270 17808
rect 14737 17731 14795 17737
rect 14737 17728 14749 17731
rect 13964 17700 14749 17728
rect 13964 17688 13970 17700
rect 14737 17697 14749 17700
rect 14783 17697 14795 17731
rect 14737 17691 14795 17697
rect 14921 17731 14979 17737
rect 14921 17697 14933 17731
rect 14967 17697 14979 17731
rect 14921 17691 14979 17697
rect 15105 17731 15163 17737
rect 15105 17697 15117 17731
rect 15151 17728 15163 17731
rect 15194 17728 15200 17740
rect 15151 17700 15200 17728
rect 15151 17697 15163 17700
rect 15105 17691 15163 17697
rect 6549 17663 6607 17669
rect 6549 17660 6561 17663
rect 6196 17632 6561 17660
rect 6549 17629 6561 17632
rect 6595 17660 6607 17663
rect 6730 17660 6736 17672
rect 6595 17632 6736 17660
rect 6595 17629 6607 17632
rect 6549 17623 6607 17629
rect 6730 17620 6736 17632
rect 6788 17620 6794 17672
rect 8202 17660 8208 17672
rect 8163 17632 8208 17660
rect 8202 17620 8208 17632
rect 8260 17620 8266 17672
rect 8294 17620 8300 17672
rect 8352 17660 8358 17672
rect 14936 17660 14964 17691
rect 15194 17688 15200 17700
rect 15252 17728 15258 17740
rect 16390 17728 16396 17740
rect 15252 17700 16396 17728
rect 15252 17688 15258 17700
rect 16390 17688 16396 17700
rect 16448 17688 16454 17740
rect 20438 17688 20444 17740
rect 20496 17728 20502 17740
rect 20717 17731 20775 17737
rect 20717 17728 20729 17731
rect 20496 17700 20729 17728
rect 20496 17688 20502 17700
rect 20717 17697 20729 17700
rect 20763 17697 20775 17731
rect 21450 17728 21456 17740
rect 21411 17700 21456 17728
rect 20717 17691 20775 17697
rect 21450 17688 21456 17700
rect 21508 17688 21514 17740
rect 16574 17660 16580 17672
rect 8352 17632 8397 17660
rect 14936 17632 16580 17660
rect 8352 17620 8358 17632
rect 16574 17620 16580 17632
rect 16632 17620 16638 17672
rect 6638 17592 6644 17604
rect 5552 17564 6644 17592
rect 6638 17552 6644 17564
rect 6696 17552 6702 17604
rect 8113 17595 8171 17601
rect 8113 17561 8125 17595
rect 8159 17592 8171 17595
rect 8478 17592 8484 17604
rect 8159 17564 8484 17592
rect 8159 17561 8171 17564
rect 8113 17555 8171 17561
rect 8478 17552 8484 17564
rect 8536 17552 8542 17604
rect 12253 17595 12311 17601
rect 12253 17561 12265 17595
rect 12299 17592 12311 17595
rect 12710 17592 12716 17604
rect 12299 17564 12716 17592
rect 12299 17561 12311 17564
rect 12253 17555 12311 17561
rect 12710 17552 12716 17564
rect 12768 17552 12774 17604
rect 5353 17527 5411 17533
rect 5353 17524 5365 17527
rect 4816 17496 5365 17524
rect 5353 17493 5365 17496
rect 5399 17493 5411 17527
rect 5353 17487 5411 17493
rect 7837 17527 7895 17533
rect 7837 17493 7849 17527
rect 7883 17524 7895 17527
rect 8386 17524 8392 17536
rect 7883 17496 8392 17524
rect 7883 17493 7895 17496
rect 7837 17487 7895 17493
rect 8386 17484 8392 17496
rect 8444 17484 8450 17536
rect 8662 17484 8668 17536
rect 8720 17524 8726 17536
rect 10134 17524 10140 17536
rect 8720 17496 10140 17524
rect 8720 17484 8726 17496
rect 10134 17484 10140 17496
rect 10192 17524 10198 17536
rect 11057 17527 11115 17533
rect 11057 17524 11069 17527
rect 10192 17496 11069 17524
rect 10192 17484 10198 17496
rect 11057 17493 11069 17496
rect 11103 17493 11115 17527
rect 12618 17524 12624 17536
rect 12579 17496 12624 17524
rect 11057 17487 11115 17493
rect 12618 17484 12624 17496
rect 12676 17484 12682 17536
rect 14553 17527 14611 17533
rect 14553 17493 14565 17527
rect 14599 17524 14611 17527
rect 14734 17524 14740 17536
rect 14599 17496 14740 17524
rect 14599 17493 14611 17496
rect 14553 17487 14611 17493
rect 14734 17484 14740 17496
rect 14792 17484 14798 17536
rect 20901 17527 20959 17533
rect 20901 17493 20913 17527
rect 20947 17524 20959 17527
rect 20990 17524 20996 17536
rect 20947 17496 20996 17524
rect 20947 17493 20959 17496
rect 20901 17487 20959 17493
rect 20990 17484 20996 17496
rect 21048 17484 21054 17536
rect 21174 17484 21180 17536
rect 21232 17524 21238 17536
rect 21269 17527 21327 17533
rect 21269 17524 21281 17527
rect 21232 17496 21281 17524
rect 21232 17484 21238 17496
rect 21269 17493 21281 17496
rect 21315 17493 21327 17527
rect 21269 17487 21327 17493
rect 1104 17434 21804 17456
rect 1104 17382 4432 17434
rect 4484 17382 4496 17434
rect 4548 17382 4560 17434
rect 4612 17382 4624 17434
rect 4676 17382 11332 17434
rect 11384 17382 11396 17434
rect 11448 17382 11460 17434
rect 11512 17382 11524 17434
rect 11576 17382 18232 17434
rect 18284 17382 18296 17434
rect 18348 17382 18360 17434
rect 18412 17382 18424 17434
rect 18476 17382 21804 17434
rect 1104 17360 21804 17382
rect 7101 17323 7159 17329
rect 7101 17289 7113 17323
rect 7147 17320 7159 17323
rect 8202 17320 8208 17332
rect 7147 17292 8208 17320
rect 7147 17289 7159 17292
rect 7101 17283 7159 17289
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 9122 17280 9128 17332
rect 9180 17320 9186 17332
rect 9490 17320 9496 17332
rect 9180 17292 9496 17320
rect 9180 17280 9186 17292
rect 9490 17280 9496 17292
rect 9548 17320 9554 17332
rect 10229 17323 10287 17329
rect 10229 17320 10241 17323
rect 9548 17292 10241 17320
rect 9548 17280 9554 17292
rect 10229 17289 10241 17292
rect 10275 17289 10287 17323
rect 10229 17283 10287 17289
rect 12618 17280 12624 17332
rect 12676 17320 12682 17332
rect 12989 17323 13047 17329
rect 12989 17320 13001 17323
rect 12676 17292 13001 17320
rect 12676 17280 12682 17292
rect 12989 17289 13001 17292
rect 13035 17289 13047 17323
rect 12989 17283 13047 17289
rect 13262 17280 13268 17332
rect 13320 17320 13326 17332
rect 13357 17323 13415 17329
rect 13357 17320 13369 17323
rect 13320 17292 13369 17320
rect 13320 17280 13326 17292
rect 13357 17289 13369 17292
rect 13403 17289 13415 17323
rect 16206 17320 16212 17332
rect 13357 17283 13415 17289
rect 14476 17292 15792 17320
rect 16167 17292 16212 17320
rect 5813 17255 5871 17261
rect 5813 17221 5825 17255
rect 5859 17252 5871 17255
rect 5902 17252 5908 17264
rect 5859 17224 5908 17252
rect 5859 17221 5871 17224
rect 5813 17215 5871 17221
rect 5902 17212 5908 17224
rect 5960 17212 5966 17264
rect 7374 17252 7380 17264
rect 6564 17224 7380 17252
rect 5920 17184 5948 17212
rect 5920 17156 6408 17184
rect 5166 17076 5172 17128
rect 5224 17116 5230 17128
rect 5537 17119 5595 17125
rect 5537 17116 5549 17119
rect 5224 17088 5549 17116
rect 5224 17076 5230 17088
rect 5537 17085 5549 17088
rect 5583 17085 5595 17119
rect 5537 17079 5595 17085
rect 5626 17076 5632 17128
rect 5684 17116 5690 17128
rect 5684 17088 5729 17116
rect 5684 17076 5690 17088
rect 5810 17076 5816 17128
rect 5868 17116 5874 17128
rect 5905 17119 5963 17125
rect 5905 17116 5917 17119
rect 5868 17088 5917 17116
rect 5868 17076 5874 17088
rect 5905 17085 5917 17088
rect 5951 17085 5963 17119
rect 5905 17079 5963 17085
rect 5997 17119 6055 17125
rect 5997 17085 6009 17119
rect 6043 17085 6055 17119
rect 6380 17116 6408 17156
rect 6454 17116 6460 17128
rect 6367 17088 6460 17116
rect 5997 17079 6055 17085
rect 5353 17051 5411 17057
rect 5353 17017 5365 17051
rect 5399 17048 5411 17051
rect 5718 17048 5724 17060
rect 5399 17020 5724 17048
rect 5399 17017 5411 17020
rect 5353 17011 5411 17017
rect 5718 17008 5724 17020
rect 5776 17048 5782 17060
rect 6012 17048 6040 17079
rect 6454 17076 6460 17088
rect 6512 17076 6518 17128
rect 6564 17116 6592 17224
rect 7374 17212 7380 17224
rect 7432 17212 7438 17264
rect 11977 17255 12035 17261
rect 11977 17221 11989 17255
rect 12023 17252 12035 17255
rect 12802 17252 12808 17264
rect 12023 17224 12808 17252
rect 12023 17221 12035 17224
rect 11977 17215 12035 17221
rect 12802 17212 12808 17224
rect 12860 17212 12866 17264
rect 6730 17184 6736 17196
rect 6691 17156 6736 17184
rect 6730 17144 6736 17156
rect 6788 17144 6794 17196
rect 12434 17144 12440 17196
rect 12492 17184 12498 17196
rect 12618 17184 12624 17196
rect 12492 17156 12537 17184
rect 12579 17156 12624 17184
rect 12492 17144 12498 17156
rect 12618 17144 12624 17156
rect 12676 17144 12682 17196
rect 14476 17193 14504 17292
rect 15764 17252 15792 17292
rect 16206 17280 16212 17292
rect 16264 17280 16270 17332
rect 15764 17224 17724 17252
rect 17696 17196 17724 17224
rect 13081 17187 13139 17193
rect 13081 17184 13093 17187
rect 12728 17156 13093 17184
rect 12728 17128 12756 17156
rect 13081 17153 13093 17156
rect 13127 17153 13139 17187
rect 13081 17147 13139 17153
rect 14461 17187 14519 17193
rect 14461 17153 14473 17187
rect 14507 17153 14519 17187
rect 14734 17184 14740 17196
rect 14695 17156 14740 17184
rect 14461 17147 14519 17153
rect 14734 17144 14740 17156
rect 14792 17144 14798 17196
rect 17678 17144 17684 17196
rect 17736 17184 17742 17196
rect 19705 17187 19763 17193
rect 19705 17184 19717 17187
rect 17736 17156 19717 17184
rect 17736 17144 17742 17156
rect 19705 17153 19717 17156
rect 19751 17153 19763 17187
rect 19705 17147 19763 17153
rect 6641 17119 6699 17125
rect 6641 17116 6653 17119
rect 6564 17088 6653 17116
rect 6641 17085 6653 17088
rect 6687 17085 6699 17119
rect 6822 17116 6828 17128
rect 6783 17088 6828 17116
rect 6641 17079 6699 17085
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 6917 17119 6975 17125
rect 6917 17085 6929 17119
rect 6963 17085 6975 17119
rect 10134 17116 10140 17128
rect 10095 17088 10140 17116
rect 6917 17079 6975 17085
rect 5776 17020 6040 17048
rect 6089 17051 6147 17057
rect 5776 17008 5782 17020
rect 6089 17017 6101 17051
rect 6135 17048 6147 17051
rect 6270 17048 6276 17060
rect 6135 17020 6276 17048
rect 6135 17017 6147 17020
rect 6089 17011 6147 17017
rect 6270 17008 6276 17020
rect 6328 17048 6334 17060
rect 6932 17048 6960 17079
rect 10134 17076 10140 17088
rect 10192 17076 10198 17128
rect 11885 17119 11943 17125
rect 11885 17085 11897 17119
rect 11931 17116 11943 17119
rect 12158 17116 12164 17128
rect 11931 17088 12164 17116
rect 11931 17085 11943 17088
rect 11885 17079 11943 17085
rect 12158 17076 12164 17088
rect 12216 17076 12222 17128
rect 12342 17116 12348 17128
rect 12303 17088 12348 17116
rect 12342 17076 12348 17088
rect 12400 17076 12406 17128
rect 12710 17116 12716 17128
rect 12671 17088 12716 17116
rect 12710 17076 12716 17088
rect 12768 17076 12774 17128
rect 12989 17119 13047 17125
rect 12989 17085 13001 17119
rect 13035 17085 13047 17119
rect 12989 17079 13047 17085
rect 6328 17020 6960 17048
rect 12176 17048 12204 17076
rect 13004 17048 13032 17079
rect 17126 17048 17132 17060
rect 12176 17020 13032 17048
rect 15962 17020 17132 17048
rect 6328 17008 6334 17020
rect 17126 17008 17132 17020
rect 17184 17048 17190 17060
rect 17586 17048 17592 17060
rect 17184 17020 17592 17048
rect 17184 17008 17190 17020
rect 17586 17008 17592 17020
rect 17644 17008 17650 17060
rect 19978 17048 19984 17060
rect 19939 17020 19984 17048
rect 19978 17008 19984 17020
rect 20036 17008 20042 17060
rect 20990 17008 20996 17060
rect 21048 17008 21054 17060
rect 17310 16940 17316 16992
rect 17368 16980 17374 16992
rect 19702 16980 19708 16992
rect 17368 16952 19708 16980
rect 17368 16940 17374 16952
rect 19702 16940 19708 16952
rect 19760 16940 19766 16992
rect 21453 16983 21511 16989
rect 21453 16949 21465 16983
rect 21499 16980 21511 16983
rect 21499 16952 21864 16980
rect 21499 16949 21511 16952
rect 21453 16943 21511 16949
rect 1104 16890 21804 16912
rect 1104 16838 7882 16890
rect 7934 16838 7946 16890
rect 7998 16838 8010 16890
rect 8062 16838 8074 16890
rect 8126 16838 14782 16890
rect 14834 16838 14846 16890
rect 14898 16838 14910 16890
rect 14962 16838 14974 16890
rect 15026 16838 21804 16890
rect 1104 16816 21804 16838
rect 16574 16736 16580 16788
rect 16632 16776 16638 16788
rect 16942 16776 16948 16788
rect 16632 16748 16948 16776
rect 16632 16736 16638 16748
rect 16942 16736 16948 16748
rect 17000 16776 17006 16788
rect 17773 16779 17831 16785
rect 17000 16748 17264 16776
rect 17000 16736 17006 16748
rect 6089 16711 6147 16717
rect 6089 16677 6101 16711
rect 6135 16677 6147 16711
rect 8386 16708 8392 16720
rect 6089 16671 6147 16677
rect 8128 16680 8392 16708
rect 5810 16640 5816 16652
rect 5771 16612 5816 16640
rect 5810 16600 5816 16612
rect 5868 16600 5874 16652
rect 5994 16600 6000 16652
rect 6052 16600 6058 16652
rect 6104 16640 6132 16671
rect 6273 16643 6331 16649
rect 6273 16640 6285 16643
rect 6104 16612 6285 16640
rect 6273 16609 6285 16612
rect 6319 16640 6331 16643
rect 6914 16640 6920 16652
rect 6319 16612 6920 16640
rect 6319 16609 6331 16612
rect 6273 16603 6331 16609
rect 6914 16600 6920 16612
rect 6972 16600 6978 16652
rect 8128 16649 8156 16680
rect 8386 16668 8392 16680
rect 8444 16668 8450 16720
rect 16850 16668 16856 16720
rect 16908 16708 16914 16720
rect 17126 16708 17132 16720
rect 16908 16680 17132 16708
rect 16908 16668 16914 16680
rect 17126 16668 17132 16680
rect 17184 16668 17190 16720
rect 17236 16717 17264 16748
rect 17773 16745 17785 16779
rect 17819 16776 17831 16779
rect 17954 16776 17960 16788
rect 17819 16748 17960 16776
rect 17819 16745 17831 16748
rect 17773 16739 17831 16745
rect 17954 16736 17960 16748
rect 18012 16736 18018 16788
rect 19978 16736 19984 16788
rect 20036 16776 20042 16788
rect 20165 16779 20223 16785
rect 20165 16776 20177 16779
rect 20036 16748 20177 16776
rect 20036 16736 20042 16748
rect 20165 16745 20177 16748
rect 20211 16745 20223 16779
rect 20165 16739 20223 16745
rect 17221 16711 17279 16717
rect 17221 16677 17233 16711
rect 17267 16677 17279 16711
rect 18598 16708 18604 16720
rect 17221 16671 17279 16677
rect 17420 16680 18604 16708
rect 8113 16643 8171 16649
rect 8113 16609 8125 16643
rect 8159 16609 8171 16643
rect 8113 16603 8171 16609
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16640 8263 16643
rect 8846 16640 8852 16652
rect 8251 16612 8852 16640
rect 8251 16609 8263 16612
rect 8205 16603 8263 16609
rect 8846 16600 8852 16612
rect 8904 16600 8910 16652
rect 15010 16600 15016 16652
rect 15068 16640 15074 16652
rect 15194 16640 15200 16652
rect 15068 16612 15200 16640
rect 15068 16600 15074 16612
rect 15194 16600 15200 16612
rect 15252 16640 15258 16652
rect 15252 16612 15976 16640
rect 15252 16600 15258 16612
rect 6012 16572 6040 16600
rect 6089 16575 6147 16581
rect 6089 16572 6101 16575
rect 6012 16544 6101 16572
rect 6089 16541 6101 16544
rect 6135 16541 6147 16575
rect 15948 16572 15976 16612
rect 16022 16600 16028 16652
rect 16080 16640 16086 16652
rect 17034 16640 17040 16652
rect 16080 16612 17040 16640
rect 16080 16600 16086 16612
rect 17034 16600 17040 16612
rect 17092 16600 17098 16652
rect 17420 16649 17448 16680
rect 18598 16668 18604 16680
rect 18656 16668 18662 16720
rect 18690 16668 18696 16720
rect 18748 16708 18754 16720
rect 19797 16711 19855 16717
rect 19797 16708 19809 16711
rect 18748 16680 19809 16708
rect 18748 16668 18754 16680
rect 19797 16677 19809 16680
rect 19843 16677 19855 16711
rect 19797 16671 19855 16677
rect 19889 16711 19947 16717
rect 19889 16677 19901 16711
rect 19935 16708 19947 16711
rect 19935 16680 20484 16708
rect 19935 16677 19947 16680
rect 19889 16671 19947 16677
rect 17405 16643 17463 16649
rect 17405 16609 17417 16643
rect 17451 16609 17463 16643
rect 17405 16603 17463 16609
rect 17497 16643 17555 16649
rect 17497 16609 17509 16643
rect 17543 16609 17555 16643
rect 17497 16603 17555 16609
rect 17512 16572 17540 16603
rect 17586 16600 17592 16652
rect 17644 16640 17650 16652
rect 19610 16640 19616 16652
rect 17644 16612 17689 16640
rect 17788 16612 19616 16640
rect 17644 16600 17650 16612
rect 17788 16572 17816 16612
rect 19610 16600 19616 16612
rect 19668 16600 19674 16652
rect 19702 16600 19708 16652
rect 19760 16640 19766 16652
rect 20456 16649 20484 16680
rect 19981 16643 20039 16649
rect 19981 16640 19993 16643
rect 19760 16612 19993 16640
rect 19760 16600 19766 16612
rect 19981 16609 19993 16612
rect 20027 16609 20039 16643
rect 19981 16603 20039 16609
rect 20441 16643 20499 16649
rect 20441 16609 20453 16643
rect 20487 16640 20499 16643
rect 21836 16640 21864 16952
rect 20487 16612 21864 16640
rect 20487 16609 20499 16612
rect 20441 16603 20499 16609
rect 15948 16544 17816 16572
rect 6089 16535 6147 16541
rect 5902 16504 5908 16516
rect 5863 16476 5908 16504
rect 5902 16464 5908 16476
rect 5960 16464 5966 16516
rect 6365 16439 6423 16445
rect 6365 16405 6377 16439
rect 6411 16436 6423 16439
rect 6546 16436 6552 16448
rect 6411 16408 6552 16436
rect 6411 16405 6423 16408
rect 6365 16399 6423 16405
rect 6546 16396 6552 16408
rect 6604 16396 6610 16448
rect 16853 16439 16911 16445
rect 16853 16405 16865 16439
rect 16899 16436 16911 16439
rect 17218 16436 17224 16448
rect 16899 16408 17224 16436
rect 16899 16405 16911 16408
rect 16853 16399 16911 16405
rect 17218 16396 17224 16408
rect 17276 16396 17282 16448
rect 19518 16396 19524 16448
rect 19576 16436 19582 16448
rect 19886 16436 19892 16448
rect 19576 16408 19892 16436
rect 19576 16396 19582 16408
rect 19886 16396 19892 16408
rect 19944 16436 19950 16448
rect 20349 16439 20407 16445
rect 20349 16436 20361 16439
rect 19944 16408 20361 16436
rect 19944 16396 19950 16408
rect 20349 16405 20361 16408
rect 20395 16405 20407 16439
rect 20349 16399 20407 16405
rect 1104 16346 21804 16368
rect 1104 16294 4432 16346
rect 4484 16294 4496 16346
rect 4548 16294 4560 16346
rect 4612 16294 4624 16346
rect 4676 16294 11332 16346
rect 11384 16294 11396 16346
rect 11448 16294 11460 16346
rect 11512 16294 11524 16346
rect 11576 16294 18232 16346
rect 18284 16294 18296 16346
rect 18348 16294 18360 16346
rect 18412 16294 18424 16346
rect 18476 16294 21804 16346
rect 1104 16272 21804 16294
rect 8389 16235 8447 16241
rect 8389 16232 8401 16235
rect 6472 16204 8401 16232
rect 1581 16031 1639 16037
rect 1581 15997 1593 16031
rect 1627 16028 1639 16031
rect 1946 16028 1952 16040
rect 1627 16000 1952 16028
rect 1627 15997 1639 16000
rect 1581 15991 1639 15997
rect 1946 15988 1952 16000
rect 2004 15988 2010 16040
rect 2133 16031 2191 16037
rect 2133 15997 2145 16031
rect 2179 16028 2191 16031
rect 2866 16028 2872 16040
rect 2179 16000 2872 16028
rect 2179 15997 2191 16000
rect 2133 15991 2191 15997
rect 2866 15988 2872 16000
rect 2924 15988 2930 16040
rect 5258 15988 5264 16040
rect 5316 16028 5322 16040
rect 6472 16037 6500 16204
rect 8389 16201 8401 16204
rect 8435 16201 8447 16235
rect 8389 16195 8447 16201
rect 14461 16235 14519 16241
rect 14461 16201 14473 16235
rect 14507 16232 14519 16235
rect 15102 16232 15108 16244
rect 14507 16204 15108 16232
rect 14507 16201 14519 16204
rect 14461 16195 14519 16201
rect 15102 16192 15108 16204
rect 15160 16192 15166 16244
rect 17586 16232 17592 16244
rect 16960 16204 17592 16232
rect 6638 16124 6644 16176
rect 6696 16164 6702 16176
rect 9306 16164 9312 16176
rect 6696 16136 9312 16164
rect 6696 16124 6702 16136
rect 9306 16124 9312 16136
rect 9364 16124 9370 16176
rect 14550 16124 14556 16176
rect 14608 16164 14614 16176
rect 15013 16167 15071 16173
rect 15013 16164 15025 16167
rect 14608 16136 15025 16164
rect 14608 16124 14614 16136
rect 15013 16133 15025 16136
rect 15059 16133 15071 16167
rect 15013 16127 15071 16133
rect 6822 16096 6828 16108
rect 6748 16068 6828 16096
rect 6457 16031 6515 16037
rect 6457 16028 6469 16031
rect 5316 16000 6469 16028
rect 5316 15988 5322 16000
rect 6457 15997 6469 16000
rect 6503 15997 6515 16031
rect 6457 15991 6515 15997
rect 6546 15988 6552 16040
rect 6604 16028 6610 16040
rect 6748 16037 6776 16068
rect 6822 16056 6828 16068
rect 6880 16096 6886 16108
rect 16206 16096 16212 16108
rect 6880 16068 7236 16096
rect 6880 16056 6886 16068
rect 6733 16031 6791 16037
rect 6604 16000 6649 16028
rect 6604 15988 6610 16000
rect 6733 15997 6745 16031
rect 6779 15997 6791 16031
rect 6914 16028 6920 16040
rect 6972 16037 6978 16040
rect 7208 16037 7236 16068
rect 8312 16068 8984 16096
rect 8312 16037 8340 16068
rect 8956 16040 8984 16068
rect 14568 16068 16212 16096
rect 6880 16000 6920 16028
rect 6733 15991 6791 15997
rect 6914 15988 6920 16000
rect 6972 15991 6980 16037
rect 7193 16031 7251 16037
rect 7193 15997 7205 16031
rect 7239 15997 7251 16031
rect 7193 15991 7251 15997
rect 8297 16031 8355 16037
rect 8297 15997 8309 16031
rect 8343 15997 8355 16031
rect 8297 15991 8355 15997
rect 8389 16031 8447 16037
rect 8389 15997 8401 16031
rect 8435 16028 8447 16031
rect 8481 16031 8539 16037
rect 8481 16028 8493 16031
rect 8435 16000 8493 16028
rect 8435 15997 8447 16000
rect 8389 15991 8447 15997
rect 8481 15997 8493 16000
rect 8527 15997 8539 16031
rect 8481 15991 8539 15997
rect 8574 16031 8632 16037
rect 8574 15997 8586 16031
rect 8620 15997 8632 16031
rect 8846 16028 8852 16040
rect 8807 16000 8852 16028
rect 8574 15991 8632 15997
rect 6972 15988 6978 15991
rect 2041 15963 2099 15969
rect 2041 15929 2053 15963
rect 2087 15960 2099 15963
rect 2682 15960 2688 15972
rect 2087 15932 2688 15960
rect 2087 15929 2099 15932
rect 2041 15923 2099 15929
rect 2682 15920 2688 15932
rect 2740 15920 2746 15972
rect 6825 15963 6883 15969
rect 6825 15929 6837 15963
rect 6871 15960 6883 15963
rect 7285 15963 7343 15969
rect 7285 15960 7297 15963
rect 6871 15932 7297 15960
rect 6871 15929 6883 15932
rect 6825 15923 6883 15929
rect 7285 15929 7297 15932
rect 7331 15929 7343 15963
rect 7285 15923 7343 15929
rect 8205 15963 8263 15969
rect 8205 15929 8217 15963
rect 8251 15960 8263 15963
rect 8588 15960 8616 15991
rect 8846 15988 8852 16000
rect 8904 15988 8910 16040
rect 8938 15988 8944 16040
rect 8996 16037 9002 16040
rect 8996 16028 9004 16037
rect 10962 16028 10968 16040
rect 8996 16000 9089 16028
rect 10923 16000 10968 16028
rect 8996 15991 9004 16000
rect 8996 15988 9002 15991
rect 10962 15988 10968 16000
rect 11020 15988 11026 16040
rect 8251 15932 8616 15960
rect 8757 15963 8815 15969
rect 8251 15929 8263 15932
rect 8205 15923 8263 15929
rect 8757 15929 8769 15963
rect 8803 15929 8815 15963
rect 8757 15923 8815 15929
rect 6914 15852 6920 15904
rect 6972 15892 6978 15904
rect 7101 15895 7159 15901
rect 7101 15892 7113 15895
rect 6972 15864 7113 15892
rect 6972 15852 6978 15864
rect 7101 15861 7113 15864
rect 7147 15861 7159 15895
rect 7101 15855 7159 15861
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 8772 15892 8800 15923
rect 9122 15892 9128 15904
rect 8444 15864 8800 15892
rect 9083 15864 9128 15892
rect 8444 15852 8450 15864
rect 9122 15852 9128 15864
rect 9180 15852 9186 15904
rect 11149 15895 11207 15901
rect 11149 15861 11161 15895
rect 11195 15892 11207 15895
rect 11238 15892 11244 15904
rect 11195 15864 11244 15892
rect 11195 15861 11207 15864
rect 11149 15855 11207 15861
rect 11238 15852 11244 15864
rect 11296 15852 11302 15904
rect 14568 15892 14596 16068
rect 15764 16037 15792 16068
rect 16206 16056 16212 16068
rect 16264 16056 16270 16108
rect 16960 16105 16988 16204
rect 17586 16192 17592 16204
rect 17644 16192 17650 16244
rect 18690 16232 18696 16244
rect 18651 16204 18696 16232
rect 18690 16192 18696 16204
rect 18748 16192 18754 16244
rect 19058 16232 19064 16244
rect 19019 16204 19064 16232
rect 19058 16192 19064 16204
rect 19116 16192 19122 16244
rect 16945 16099 17003 16105
rect 16945 16065 16957 16099
rect 16991 16065 17003 16099
rect 17218 16096 17224 16108
rect 17179 16068 17224 16096
rect 16945 16059 17003 16065
rect 17218 16056 17224 16068
rect 17276 16056 17282 16108
rect 19260 16068 20024 16096
rect 14642 16031 14700 16037
rect 14642 15997 14654 16031
rect 14688 15997 14700 16031
rect 14642 15991 14700 15997
rect 15105 16031 15163 16037
rect 15105 15997 15117 16031
rect 15151 16028 15163 16031
rect 15381 16031 15439 16037
rect 15381 16028 15393 16031
rect 15151 16000 15393 16028
rect 15151 15997 15163 16000
rect 15105 15991 15163 15997
rect 15381 15997 15393 16000
rect 15427 15997 15439 16031
rect 15381 15991 15439 15997
rect 15657 16031 15715 16037
rect 15657 15997 15669 16031
rect 15703 16028 15715 16031
rect 15749 16031 15807 16037
rect 15749 16028 15761 16031
rect 15703 16000 15761 16028
rect 15703 15997 15715 16000
rect 15657 15991 15715 15997
rect 15749 15997 15761 16000
rect 15795 15997 15807 16031
rect 15749 15991 15807 15997
rect 15933 16031 15991 16037
rect 15933 15997 15945 16031
rect 15979 16028 15991 16031
rect 16850 16028 16856 16040
rect 15979 16000 16856 16028
rect 15979 15997 15991 16000
rect 15933 15991 15991 15997
rect 14657 15960 14685 15991
rect 15396 15960 15424 15991
rect 15841 15963 15899 15969
rect 15841 15960 15853 15963
rect 14657 15932 15332 15960
rect 15396 15932 15853 15960
rect 14645 15895 14703 15901
rect 14645 15892 14657 15895
rect 14568 15864 14657 15892
rect 14645 15861 14657 15864
rect 14691 15861 14703 15895
rect 15194 15892 15200 15904
rect 15155 15864 15200 15892
rect 14645 15855 14703 15861
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 15304 15892 15332 15932
rect 15841 15929 15853 15932
rect 15887 15929 15899 15963
rect 15841 15923 15899 15929
rect 15565 15895 15623 15901
rect 15565 15892 15577 15895
rect 15304 15864 15577 15892
rect 15565 15861 15577 15864
rect 15611 15892 15623 15895
rect 15948 15892 15976 15991
rect 16850 15988 16856 16000
rect 16908 15988 16914 16040
rect 19260 16037 19288 16068
rect 19245 16031 19303 16037
rect 19245 15997 19257 16031
rect 19291 15997 19303 16031
rect 19245 15991 19303 15997
rect 19518 15988 19524 16040
rect 19576 16028 19582 16040
rect 19705 16031 19763 16037
rect 19576 16000 19621 16028
rect 19576 15988 19582 16000
rect 19705 15997 19717 16031
rect 19751 15997 19763 16031
rect 19886 16028 19892 16040
rect 19847 16000 19892 16028
rect 19705 15991 19763 15997
rect 17954 15920 17960 15972
rect 18012 15920 18018 15972
rect 18598 15920 18604 15972
rect 18656 15960 18662 15972
rect 18966 15960 18972 15972
rect 18656 15932 18972 15960
rect 18656 15920 18662 15932
rect 18966 15920 18972 15932
rect 19024 15960 19030 15972
rect 19429 15963 19487 15969
rect 19429 15960 19441 15963
rect 19024 15932 19441 15960
rect 19024 15920 19030 15932
rect 19429 15929 19441 15932
rect 19475 15960 19487 15963
rect 19720 15960 19748 15991
rect 19886 15988 19892 16000
rect 19944 15988 19950 16040
rect 19996 15972 20024 16068
rect 19475 15932 19748 15960
rect 19475 15929 19487 15932
rect 19429 15923 19487 15929
rect 19978 15920 19984 15972
rect 20036 15960 20042 15972
rect 20036 15932 20081 15960
rect 20036 15920 20042 15932
rect 15611 15864 15976 15892
rect 15611 15861 15623 15864
rect 15565 15855 15623 15861
rect 1104 15802 21804 15824
rect 1104 15750 7882 15802
rect 7934 15750 7946 15802
rect 7998 15750 8010 15802
rect 8062 15750 8074 15802
rect 8126 15750 14782 15802
rect 14834 15750 14846 15802
rect 14898 15750 14910 15802
rect 14962 15750 14974 15802
rect 15026 15750 21804 15802
rect 1104 15728 21804 15750
rect 8849 15691 8907 15697
rect 8849 15657 8861 15691
rect 8895 15688 8907 15691
rect 8938 15688 8944 15700
rect 8895 15660 8944 15688
rect 8895 15657 8907 15660
rect 8849 15651 8907 15657
rect 8938 15648 8944 15660
rect 8996 15648 9002 15700
rect 9030 15648 9036 15700
rect 9088 15688 9094 15700
rect 9861 15691 9919 15697
rect 9861 15688 9873 15691
rect 9088 15660 9873 15688
rect 9088 15648 9094 15660
rect 9861 15657 9873 15660
rect 9907 15657 9919 15691
rect 12158 15688 12164 15700
rect 12119 15660 12164 15688
rect 9861 15651 9919 15657
rect 12158 15648 12164 15660
rect 12216 15648 12222 15700
rect 12805 15691 12863 15697
rect 12805 15657 12817 15691
rect 12851 15688 12863 15691
rect 12897 15691 12955 15697
rect 12897 15688 12909 15691
rect 12851 15660 12909 15688
rect 12851 15657 12863 15660
rect 12805 15651 12863 15657
rect 12897 15657 12909 15660
rect 12943 15688 12955 15691
rect 12986 15688 12992 15700
rect 12943 15660 12992 15688
rect 12943 15657 12955 15660
rect 12897 15651 12955 15657
rect 12986 15648 12992 15660
rect 13044 15648 13050 15700
rect 14369 15691 14427 15697
rect 14369 15688 14381 15691
rect 13280 15660 14381 15688
rect 8754 15620 8760 15632
rect 8588 15592 8760 15620
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 2593 15555 2651 15561
rect 2593 15521 2605 15555
rect 2639 15552 2651 15555
rect 3053 15555 3111 15561
rect 3053 15552 3065 15555
rect 2639 15524 3065 15552
rect 2639 15521 2651 15524
rect 2593 15515 2651 15521
rect 3053 15521 3065 15524
rect 3099 15521 3111 15555
rect 3234 15552 3240 15564
rect 3195 15524 3240 15552
rect 3053 15515 3111 15521
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 8297 15555 8355 15561
rect 8297 15521 8309 15555
rect 8343 15521 8355 15555
rect 8297 15515 8355 15521
rect 1946 15444 1952 15496
rect 2004 15484 2010 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 2004 15456 2053 15484
rect 2004 15444 2010 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 2041 15447 2099 15453
rect 2501 15419 2559 15425
rect 2501 15385 2513 15419
rect 2547 15416 2559 15419
rect 2682 15416 2688 15428
rect 2547 15388 2688 15416
rect 2547 15385 2559 15388
rect 2501 15379 2559 15385
rect 2682 15376 2688 15388
rect 2740 15376 2746 15428
rect 8312 15416 8340 15515
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 8588 15561 8616 15592
rect 8754 15580 8760 15592
rect 8812 15580 8818 15632
rect 9125 15623 9183 15629
rect 9125 15589 9137 15623
rect 9171 15620 9183 15623
rect 10229 15623 10287 15629
rect 10229 15620 10241 15623
rect 9171 15592 10241 15620
rect 9171 15589 9183 15592
rect 9125 15583 9183 15589
rect 10229 15589 10241 15592
rect 10275 15589 10287 15623
rect 10229 15583 10287 15589
rect 11238 15580 11244 15632
rect 11296 15580 11302 15632
rect 13280 15629 13308 15660
rect 14369 15657 14381 15660
rect 14415 15657 14427 15691
rect 14369 15651 14427 15657
rect 14553 15691 14611 15697
rect 14553 15657 14565 15691
rect 14599 15688 14611 15691
rect 17126 15688 17132 15700
rect 14599 15660 14964 15688
rect 17087 15660 17132 15688
rect 14599 15657 14611 15660
rect 14553 15651 14611 15657
rect 13265 15623 13323 15629
rect 13265 15620 13277 15623
rect 12360 15592 13277 15620
rect 8573 15555 8631 15561
rect 8573 15552 8585 15555
rect 8536 15524 8585 15552
rect 8536 15512 8542 15524
rect 8573 15521 8585 15524
rect 8619 15521 8631 15555
rect 8573 15515 8631 15521
rect 8665 15555 8723 15561
rect 8665 15521 8677 15555
rect 8711 15552 8723 15555
rect 9401 15555 9459 15561
rect 9401 15552 9413 15555
rect 8711 15524 9413 15552
rect 8711 15521 8723 15524
rect 8665 15515 8723 15521
rect 9401 15521 9413 15524
rect 9447 15552 9459 15555
rect 9582 15552 9588 15564
rect 9447 15524 9588 15552
rect 9447 15521 9459 15524
rect 9401 15515 9459 15521
rect 9582 15512 9588 15524
rect 9640 15512 9646 15564
rect 12360 15561 12388 15592
rect 13265 15589 13277 15592
rect 13311 15589 13323 15623
rect 13265 15583 13323 15589
rect 9861 15555 9919 15561
rect 9861 15521 9873 15555
rect 9907 15552 9919 15555
rect 9953 15555 10011 15561
rect 9953 15552 9965 15555
rect 9907 15524 9965 15552
rect 9907 15521 9919 15524
rect 9861 15515 9919 15521
rect 9953 15521 9965 15524
rect 9999 15521 10011 15555
rect 9953 15515 10011 15521
rect 12345 15555 12403 15561
rect 12345 15521 12357 15555
rect 12391 15521 12403 15555
rect 12345 15515 12403 15521
rect 13081 15555 13139 15561
rect 13081 15521 13093 15555
rect 13127 15521 13139 15555
rect 14550 15552 14556 15564
rect 14511 15524 14556 15552
rect 13081 15515 13139 15521
rect 9122 15484 9128 15496
rect 9083 15456 9128 15484
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 9306 15484 9312 15496
rect 9267 15456 9312 15484
rect 9306 15444 9312 15456
rect 9364 15444 9370 15496
rect 12437 15487 12495 15493
rect 12437 15453 12449 15487
rect 12483 15484 12495 15487
rect 12526 15484 12532 15496
rect 12483 15456 12532 15484
rect 12483 15453 12495 15456
rect 12437 15447 12495 15453
rect 12526 15444 12532 15456
rect 12584 15484 12590 15496
rect 13096 15484 13124 15515
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 14936 15561 14964 15660
rect 17126 15648 17132 15660
rect 17184 15648 17190 15700
rect 17310 15688 17316 15700
rect 17271 15660 17316 15688
rect 17310 15648 17316 15660
rect 17368 15688 17374 15700
rect 17678 15688 17684 15700
rect 17368 15660 17684 15688
rect 17368 15648 17374 15660
rect 17678 15648 17684 15660
rect 17736 15648 17742 15700
rect 19426 15648 19432 15700
rect 19484 15688 19490 15700
rect 19889 15691 19947 15697
rect 19889 15688 19901 15691
rect 19484 15660 19901 15688
rect 19484 15648 19490 15660
rect 19889 15657 19901 15660
rect 19935 15657 19947 15691
rect 19889 15651 19947 15657
rect 20073 15691 20131 15697
rect 20073 15657 20085 15691
rect 20119 15688 20131 15691
rect 20162 15688 20168 15700
rect 20119 15660 20168 15688
rect 20119 15657 20131 15660
rect 20073 15651 20131 15657
rect 16942 15620 16948 15632
rect 16903 15592 16948 15620
rect 16942 15580 16948 15592
rect 17000 15580 17006 15632
rect 17034 15580 17040 15632
rect 17092 15620 17098 15632
rect 17221 15623 17279 15629
rect 17221 15620 17233 15623
rect 17092 15592 17233 15620
rect 17092 15580 17098 15592
rect 17221 15589 17233 15592
rect 17267 15589 17279 15623
rect 17221 15583 17279 15589
rect 14921 15555 14979 15561
rect 14921 15521 14933 15555
rect 14967 15552 14979 15555
rect 15194 15552 15200 15564
rect 14967 15524 15200 15552
rect 14967 15521 14979 15524
rect 14921 15515 14979 15521
rect 15194 15512 15200 15524
rect 15252 15512 15258 15564
rect 19613 15555 19671 15561
rect 19613 15521 19625 15555
rect 19659 15521 19671 15555
rect 19613 15515 19671 15521
rect 19797 15555 19855 15561
rect 19797 15521 19809 15555
rect 19843 15552 19855 15555
rect 20088 15552 20116 15651
rect 20162 15648 20168 15660
rect 20220 15648 20226 15700
rect 21266 15688 21272 15700
rect 21227 15660 21272 15688
rect 21266 15648 21272 15660
rect 21324 15648 21330 15700
rect 19843 15524 20116 15552
rect 20165 15555 20223 15561
rect 19843 15521 19855 15524
rect 19797 15515 19855 15521
rect 20165 15521 20177 15555
rect 20211 15521 20223 15555
rect 21450 15552 21456 15564
rect 21411 15524 21456 15552
rect 20165 15515 20223 15521
rect 12584 15456 13124 15484
rect 14568 15484 14596 15512
rect 15013 15487 15071 15493
rect 15013 15484 15025 15487
rect 14568 15456 15025 15484
rect 12584 15444 12590 15456
rect 15013 15453 15025 15456
rect 15059 15453 15071 15487
rect 19628 15484 19656 15515
rect 19978 15484 19984 15496
rect 19628 15456 19984 15484
rect 15013 15447 15071 15453
rect 19978 15444 19984 15456
rect 20036 15484 20042 15496
rect 20180 15484 20208 15515
rect 21450 15512 21456 15524
rect 21508 15512 21514 15564
rect 20036 15456 20208 15484
rect 20036 15444 20042 15456
rect 9858 15416 9864 15428
rect 8312 15388 9864 15416
rect 9858 15376 9864 15388
rect 9916 15376 9922 15428
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15348 1639 15351
rect 1854 15348 1860 15360
rect 1627 15320 1860 15348
rect 1627 15317 1639 15320
rect 1581 15311 1639 15317
rect 1854 15308 1860 15320
rect 1912 15308 1918 15360
rect 5626 15308 5632 15360
rect 5684 15348 5690 15360
rect 7282 15348 7288 15360
rect 5684 15320 7288 15348
rect 5684 15308 5690 15320
rect 7282 15308 7288 15320
rect 7340 15348 7346 15360
rect 8389 15351 8447 15357
rect 8389 15348 8401 15351
rect 7340 15320 8401 15348
rect 7340 15308 7346 15320
rect 8389 15317 8401 15320
rect 8435 15317 8447 15351
rect 9876 15348 9904 15376
rect 10870 15348 10876 15360
rect 9876 15320 10876 15348
rect 8389 15311 8447 15317
rect 10870 15308 10876 15320
rect 10928 15348 10934 15360
rect 11701 15351 11759 15357
rect 11701 15348 11713 15351
rect 10928 15320 11713 15348
rect 10928 15308 10934 15320
rect 11701 15317 11713 15320
rect 11747 15317 11759 15351
rect 11701 15311 11759 15317
rect 17497 15351 17555 15357
rect 17497 15317 17509 15351
rect 17543 15348 17555 15351
rect 18598 15348 18604 15360
rect 17543 15320 18604 15348
rect 17543 15317 17555 15320
rect 17497 15311 17555 15317
rect 18598 15308 18604 15320
rect 18656 15308 18662 15360
rect 1104 15258 21804 15280
rect 1104 15206 4432 15258
rect 4484 15206 4496 15258
rect 4548 15206 4560 15258
rect 4612 15206 4624 15258
rect 4676 15206 11332 15258
rect 11384 15206 11396 15258
rect 11448 15206 11460 15258
rect 11512 15206 11524 15258
rect 11576 15206 18232 15258
rect 18284 15206 18296 15258
rect 18348 15206 18360 15258
rect 18412 15206 18424 15258
rect 18476 15206 21804 15258
rect 1104 15184 21804 15206
rect 1581 15147 1639 15153
rect 1581 15113 1593 15147
rect 1627 15144 1639 15147
rect 1946 15144 1952 15156
rect 1627 15116 1952 15144
rect 1627 15113 1639 15116
rect 1581 15107 1639 15113
rect 1946 15104 1952 15116
rect 2004 15104 2010 15156
rect 6638 15144 6644 15156
rect 6599 15116 6644 15144
rect 6638 15104 6644 15116
rect 6696 15104 6702 15156
rect 6822 15144 6828 15156
rect 6783 15116 6828 15144
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 7282 15144 7288 15156
rect 7243 15116 7288 15144
rect 7282 15104 7288 15116
rect 7340 15104 7346 15156
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 13081 15147 13139 15153
rect 13081 15144 13093 15147
rect 12492 15116 13093 15144
rect 12492 15104 12498 15116
rect 13081 15113 13093 15116
rect 13127 15113 13139 15147
rect 13081 15107 13139 15113
rect 3881 15079 3939 15085
rect 3881 15045 3893 15079
rect 3927 15076 3939 15079
rect 3973 15079 4031 15085
rect 3973 15076 3985 15079
rect 3927 15048 3985 15076
rect 3927 15045 3939 15048
rect 3881 15039 3939 15045
rect 3973 15045 3985 15048
rect 4019 15045 4031 15079
rect 9493 15079 9551 15085
rect 9493 15076 9505 15079
rect 3973 15039 4031 15045
rect 5460 15048 9505 15076
rect 2038 15008 2044 15020
rect 1999 14980 2044 15008
rect 2038 14968 2044 14980
rect 2096 14968 2102 15020
rect 2133 15011 2191 15017
rect 2133 14977 2145 15011
rect 2179 14977 2191 15011
rect 3513 15011 3571 15017
rect 3513 15008 3525 15011
rect 2133 14971 2191 14977
rect 3436 14980 3525 15008
rect 1762 14900 1768 14952
rect 1820 14940 1826 14952
rect 2148 14940 2176 14971
rect 2866 14940 2872 14952
rect 1820 14912 2176 14940
rect 2827 14912 2872 14940
rect 1820 14900 1826 14912
rect 2866 14900 2872 14912
rect 2924 14940 2930 14952
rect 3436 14949 3464 14980
rect 3513 14977 3525 14980
rect 3559 15008 3571 15011
rect 5460 15008 5488 15048
rect 9493 15045 9505 15048
rect 9539 15045 9551 15079
rect 9493 15039 9551 15045
rect 9582 15036 9588 15088
rect 9640 15076 9646 15088
rect 10321 15079 10379 15085
rect 10321 15076 10333 15079
rect 9640 15048 10333 15076
rect 9640 15036 9646 15048
rect 10321 15045 10333 15048
rect 10367 15045 10379 15079
rect 14277 15079 14335 15085
rect 14277 15076 14289 15079
rect 10321 15039 10379 15045
rect 13648 15048 14289 15076
rect 3559 14980 5488 15008
rect 6457 15011 6515 15017
rect 3559 14977 3571 14980
rect 3513 14971 3571 14977
rect 6457 14977 6469 15011
rect 6503 15008 6515 15011
rect 6914 15008 6920 15020
rect 6503 14980 6920 15008
rect 6503 14977 6515 14980
rect 6457 14971 6515 14977
rect 6914 14968 6920 14980
rect 6972 14968 6978 15020
rect 8478 15008 8484 15020
rect 7116 14980 8484 15008
rect 3421 14943 3479 14949
rect 2924 14912 3372 14940
rect 2924 14900 2930 14912
rect 3344 14884 3372 14912
rect 3421 14909 3433 14943
rect 3467 14909 3479 14943
rect 3421 14903 3479 14909
rect 4157 14943 4215 14949
rect 4157 14909 4169 14943
rect 4203 14909 4215 14943
rect 4157 14903 4215 14909
rect 5077 14943 5135 14949
rect 5077 14909 5089 14943
rect 5123 14940 5135 14943
rect 5258 14940 5264 14952
rect 5123 14912 5264 14940
rect 5123 14909 5135 14912
rect 5077 14903 5135 14909
rect 2961 14875 3019 14881
rect 2961 14841 2973 14875
rect 3007 14841 3019 14875
rect 3326 14872 3332 14884
rect 3239 14844 3332 14872
rect 2961 14835 3019 14841
rect 1946 14804 1952 14816
rect 1907 14776 1952 14804
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 2976 14804 3004 14835
rect 3326 14832 3332 14844
rect 3384 14872 3390 14884
rect 4172 14872 4200 14903
rect 5258 14900 5264 14912
rect 5316 14900 5322 14952
rect 6733 14943 6791 14949
rect 6733 14909 6745 14943
rect 6779 14909 6791 14943
rect 7006 14940 7012 14952
rect 6967 14912 7012 14940
rect 6733 14903 6791 14909
rect 3384 14844 4200 14872
rect 6748 14872 6776 14903
rect 7006 14900 7012 14912
rect 7064 14900 7070 14952
rect 7116 14949 7144 14980
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 15008 10103 15011
rect 12066 15008 12072 15020
rect 10091 14980 12072 15008
rect 10091 14977 10103 14980
rect 10045 14971 10103 14977
rect 12066 14968 12072 14980
rect 12124 14968 12130 15020
rect 13648 15017 13676 15048
rect 14277 15045 14289 15048
rect 14323 15045 14335 15079
rect 14277 15039 14335 15045
rect 13633 15011 13691 15017
rect 13633 15008 13645 15011
rect 13372 14980 13645 15008
rect 7101 14943 7159 14949
rect 7101 14909 7113 14943
rect 7147 14909 7159 14943
rect 7101 14903 7159 14909
rect 7377 14943 7435 14949
rect 7377 14909 7389 14943
rect 7423 14940 7435 14943
rect 7558 14940 7564 14952
rect 7423 14912 7564 14940
rect 7423 14909 7435 14912
rect 7377 14903 7435 14909
rect 7392 14872 7420 14903
rect 7558 14900 7564 14912
rect 7616 14900 7622 14952
rect 9858 14900 9864 14952
rect 9916 14940 9922 14952
rect 13372 14949 13400 14980
rect 13633 14977 13645 14980
rect 13679 14977 13691 15011
rect 13633 14971 13691 14977
rect 13725 15011 13783 15017
rect 13725 14977 13737 15011
rect 13771 15008 13783 15011
rect 13771 14980 15792 15008
rect 13771 14977 13783 14980
rect 13725 14971 13783 14977
rect 10229 14943 10287 14949
rect 10229 14940 10241 14943
rect 9916 14912 10241 14940
rect 9916 14900 9922 14912
rect 10229 14909 10241 14912
rect 10275 14909 10287 14943
rect 10229 14903 10287 14909
rect 13265 14943 13323 14949
rect 13265 14909 13277 14943
rect 13311 14909 13323 14943
rect 13265 14903 13323 14909
rect 13357 14943 13415 14949
rect 13357 14909 13369 14943
rect 13403 14909 13415 14943
rect 13357 14903 13415 14909
rect 9766 14872 9772 14884
rect 6748 14844 7420 14872
rect 9727 14844 9772 14872
rect 3384 14832 3390 14844
rect 9766 14832 9772 14844
rect 9824 14832 9830 14884
rect 11146 14872 11152 14884
rect 10244 14844 11152 14872
rect 3234 14804 3240 14816
rect 2976 14776 3240 14804
rect 3234 14764 3240 14776
rect 3292 14804 3298 14816
rect 3881 14807 3939 14813
rect 3881 14804 3893 14807
rect 3292 14776 3893 14804
rect 3292 14764 3298 14776
rect 3881 14773 3893 14776
rect 3927 14773 3939 14807
rect 4890 14804 4896 14816
rect 4851 14776 4896 14804
rect 3881 14767 3939 14773
rect 4890 14764 4896 14776
rect 4948 14764 4954 14816
rect 5626 14764 5632 14816
rect 5684 14804 5690 14816
rect 6457 14807 6515 14813
rect 6457 14804 6469 14807
rect 5684 14776 6469 14804
rect 5684 14764 5690 14776
rect 6457 14773 6469 14776
rect 6503 14773 6515 14807
rect 6457 14767 6515 14773
rect 9953 14807 10011 14813
rect 9953 14773 9965 14807
rect 9999 14804 10011 14807
rect 10244 14804 10272 14844
rect 11146 14832 11152 14844
rect 11204 14832 11210 14884
rect 13280 14872 13308 14903
rect 13740 14872 13768 14971
rect 14553 14943 14611 14949
rect 14553 14909 14565 14943
rect 14599 14940 14611 14943
rect 14642 14940 14648 14952
rect 14599 14912 14648 14940
rect 14599 14909 14611 14912
rect 14553 14903 14611 14909
rect 14642 14900 14648 14912
rect 14700 14900 14706 14952
rect 13280 14844 13768 14872
rect 14277 14875 14335 14881
rect 14277 14841 14289 14875
rect 14323 14872 14335 14875
rect 15194 14872 15200 14884
rect 14323 14844 15200 14872
rect 14323 14841 14335 14844
rect 14277 14835 14335 14841
rect 15194 14832 15200 14844
rect 15252 14832 15258 14884
rect 15764 14816 15792 14980
rect 19797 14943 19855 14949
rect 19797 14909 19809 14943
rect 19843 14909 19855 14943
rect 19978 14940 19984 14952
rect 19939 14912 19984 14940
rect 19797 14903 19855 14909
rect 9999 14776 10272 14804
rect 14461 14807 14519 14813
rect 9999 14773 10011 14776
rect 9953 14767 10011 14773
rect 14461 14773 14473 14807
rect 14507 14804 14519 14807
rect 15562 14804 15568 14816
rect 14507 14776 15568 14804
rect 14507 14773 14519 14776
rect 14461 14767 14519 14773
rect 15562 14764 15568 14776
rect 15620 14764 15626 14816
rect 15746 14764 15752 14816
rect 15804 14804 15810 14816
rect 19613 14807 19671 14813
rect 19613 14804 19625 14807
rect 15804 14776 19625 14804
rect 15804 14764 15810 14776
rect 19613 14773 19625 14776
rect 19659 14773 19671 14807
rect 19812 14804 19840 14903
rect 19978 14900 19984 14912
rect 20036 14900 20042 14952
rect 20162 14940 20168 14952
rect 20123 14912 20168 14940
rect 20162 14900 20168 14912
rect 20220 14900 20226 14952
rect 19886 14832 19892 14884
rect 19944 14872 19950 14884
rect 19944 14844 19989 14872
rect 19944 14832 19950 14844
rect 20346 14804 20352 14816
rect 19812 14776 20352 14804
rect 19613 14767 19671 14773
rect 20346 14764 20352 14776
rect 20404 14764 20410 14816
rect 1104 14714 21804 14736
rect 1104 14662 7882 14714
rect 7934 14662 7946 14714
rect 7998 14662 8010 14714
rect 8062 14662 8074 14714
rect 8126 14662 14782 14714
rect 14834 14662 14846 14714
rect 14898 14662 14910 14714
rect 14962 14662 14974 14714
rect 15026 14662 21804 14714
rect 1104 14640 21804 14662
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 7282 14600 7288 14612
rect 5316 14572 7288 14600
rect 5316 14560 5322 14572
rect 7282 14560 7288 14572
rect 7340 14600 7346 14612
rect 10962 14600 10968 14612
rect 7340 14572 10968 14600
rect 7340 14560 7346 14572
rect 10962 14560 10968 14572
rect 11020 14560 11026 14612
rect 14550 14600 14556 14612
rect 14511 14572 14556 14600
rect 14550 14560 14556 14572
rect 14608 14560 14614 14612
rect 14642 14560 14648 14612
rect 14700 14600 14706 14612
rect 14737 14603 14795 14609
rect 14737 14600 14749 14603
rect 14700 14572 14749 14600
rect 14700 14560 14706 14572
rect 14737 14569 14749 14572
rect 14783 14569 14795 14603
rect 14737 14563 14795 14569
rect 4890 14492 4896 14544
rect 4948 14492 4954 14544
rect 5626 14532 5632 14544
rect 5587 14504 5632 14532
rect 5626 14492 5632 14504
rect 5684 14492 5690 14544
rect 14752 14532 14780 14563
rect 17126 14560 17132 14612
rect 17184 14600 17190 14612
rect 17313 14603 17371 14609
rect 17313 14600 17325 14603
rect 17184 14572 17325 14600
rect 17184 14560 17190 14572
rect 17313 14569 17325 14572
rect 17359 14569 17371 14603
rect 18966 14600 18972 14612
rect 18927 14572 18972 14600
rect 17313 14563 17371 14569
rect 18966 14560 18972 14572
rect 19024 14560 19030 14612
rect 20162 14600 20168 14612
rect 20123 14572 20168 14600
rect 20162 14560 20168 14572
rect 20220 14560 20226 14612
rect 20346 14600 20352 14612
rect 20307 14572 20352 14600
rect 20346 14560 20352 14572
rect 20404 14560 20410 14612
rect 15381 14535 15439 14541
rect 15381 14532 15393 14535
rect 14752 14504 14872 14532
rect 5905 14467 5963 14473
rect 5905 14433 5917 14467
rect 5951 14464 5963 14467
rect 8478 14464 8484 14476
rect 5951 14436 8484 14464
rect 5951 14433 5963 14436
rect 5905 14427 5963 14433
rect 8478 14424 8484 14436
rect 8536 14464 8542 14476
rect 9030 14464 9036 14476
rect 8536 14436 9036 14464
rect 8536 14424 8542 14436
rect 9030 14424 9036 14436
rect 9088 14424 9094 14476
rect 12805 14467 12863 14473
rect 12805 14433 12817 14467
rect 12851 14464 12863 14467
rect 13906 14464 13912 14476
rect 12851 14436 13912 14464
rect 12851 14433 12863 14436
rect 12805 14427 12863 14433
rect 13906 14424 13912 14436
rect 13964 14424 13970 14476
rect 14734 14467 14792 14473
rect 14734 14433 14746 14467
rect 14780 14433 14792 14467
rect 14734 14427 14792 14433
rect 12897 14399 12955 14405
rect 12897 14365 12909 14399
rect 12943 14396 12955 14399
rect 13814 14396 13820 14408
rect 12943 14368 13820 14396
rect 12943 14365 12955 14368
rect 12897 14359 12955 14365
rect 13814 14356 13820 14368
rect 13872 14356 13878 14408
rect 4157 14263 4215 14269
rect 4157 14229 4169 14263
rect 4203 14260 4215 14263
rect 5258 14260 5264 14272
rect 4203 14232 5264 14260
rect 4203 14229 4215 14232
rect 4157 14223 4215 14229
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 6822 14220 6828 14272
rect 6880 14260 6886 14272
rect 7742 14260 7748 14272
rect 6880 14232 7748 14260
rect 6880 14220 6886 14232
rect 7742 14220 7748 14232
rect 7800 14260 7806 14272
rect 8662 14260 8668 14272
rect 7800 14232 8668 14260
rect 7800 14220 7806 14232
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 14752 14260 14780 14427
rect 14844 14396 14872 14504
rect 15212 14504 15393 14532
rect 15212 14476 15240 14504
rect 15381 14501 15393 14504
rect 15427 14501 15439 14535
rect 15381 14495 15439 14501
rect 15194 14464 15200 14476
rect 15155 14436 15200 14464
rect 15194 14424 15200 14436
rect 15252 14424 15258 14476
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 15473 14467 15531 14473
rect 15473 14433 15485 14467
rect 15519 14464 15531 14467
rect 15562 14464 15568 14476
rect 15519 14436 15568 14464
rect 15519 14433 15531 14436
rect 15473 14427 15531 14433
rect 15304 14396 15332 14427
rect 15562 14424 15568 14436
rect 15620 14424 15626 14476
rect 15746 14464 15752 14476
rect 15707 14436 15752 14464
rect 15746 14424 15752 14436
rect 15804 14424 15810 14476
rect 17405 14467 17463 14473
rect 17405 14433 17417 14467
rect 17451 14464 17463 14467
rect 18046 14464 18052 14476
rect 17451 14436 18052 14464
rect 17451 14433 17463 14436
rect 17405 14427 17463 14433
rect 18046 14424 18052 14436
rect 18104 14424 18110 14476
rect 18690 14424 18696 14476
rect 18748 14464 18754 14476
rect 18877 14467 18935 14473
rect 18877 14464 18889 14467
rect 18748 14436 18889 14464
rect 18748 14424 18754 14436
rect 18877 14433 18889 14436
rect 18923 14464 18935 14467
rect 19150 14464 19156 14476
rect 18923 14436 19156 14464
rect 18923 14433 18935 14436
rect 18877 14427 18935 14433
rect 19150 14424 19156 14436
rect 19208 14424 19214 14476
rect 19334 14424 19340 14476
rect 19392 14464 19398 14476
rect 19886 14464 19892 14476
rect 19392 14436 19892 14464
rect 19392 14424 19398 14436
rect 19886 14424 19892 14436
rect 19944 14464 19950 14476
rect 20290 14467 20348 14473
rect 20290 14464 20302 14467
rect 19944 14436 20302 14464
rect 19944 14424 19950 14436
rect 20290 14433 20302 14436
rect 20336 14464 20348 14467
rect 20809 14467 20867 14473
rect 20809 14464 20821 14467
rect 20336 14436 20821 14464
rect 20336 14433 20348 14436
rect 20290 14427 20348 14433
rect 20809 14433 20821 14436
rect 20855 14433 20867 14467
rect 20809 14427 20867 14433
rect 14844 14368 15332 14396
rect 15105 14331 15163 14337
rect 15105 14297 15117 14331
rect 15151 14328 15163 14331
rect 15657 14331 15715 14337
rect 15657 14328 15669 14331
rect 15151 14300 15669 14328
rect 15151 14297 15163 14300
rect 15105 14291 15163 14297
rect 15657 14297 15669 14300
rect 15703 14297 15715 14331
rect 15657 14291 15715 14297
rect 15562 14260 15568 14272
rect 14752 14232 15568 14260
rect 15562 14220 15568 14232
rect 15620 14220 15626 14272
rect 20070 14220 20076 14272
rect 20128 14260 20134 14272
rect 20346 14260 20352 14272
rect 20128 14232 20352 14260
rect 20128 14220 20134 14232
rect 20346 14220 20352 14232
rect 20404 14260 20410 14272
rect 20717 14263 20775 14269
rect 20717 14260 20729 14263
rect 20404 14232 20729 14260
rect 20404 14220 20410 14232
rect 20717 14229 20729 14232
rect 20763 14229 20775 14263
rect 20717 14223 20775 14229
rect 1104 14170 21804 14192
rect 1104 14118 4432 14170
rect 4484 14118 4496 14170
rect 4548 14118 4560 14170
rect 4612 14118 4624 14170
rect 4676 14118 11332 14170
rect 11384 14118 11396 14170
rect 11448 14118 11460 14170
rect 11512 14118 11524 14170
rect 11576 14118 18232 14170
rect 18284 14118 18296 14170
rect 18348 14118 18360 14170
rect 18412 14118 18424 14170
rect 18476 14118 21804 14170
rect 1104 14096 21804 14118
rect 1946 14016 1952 14068
rect 2004 14056 2010 14068
rect 6457 14059 6515 14065
rect 6457 14056 6469 14059
rect 2004 14028 6469 14056
rect 2004 14016 2010 14028
rect 6457 14025 6469 14028
rect 6503 14025 6515 14059
rect 6457 14019 6515 14025
rect 7101 14059 7159 14065
rect 7101 14025 7113 14059
rect 7147 14056 7159 14059
rect 7466 14056 7472 14068
rect 7147 14028 7472 14056
rect 7147 14025 7159 14028
rect 7101 14019 7159 14025
rect 7466 14016 7472 14028
rect 7524 14056 7530 14068
rect 8018 14056 8024 14068
rect 7524 14028 8024 14056
rect 7524 14016 7530 14028
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 8113 14059 8171 14065
rect 8113 14025 8125 14059
rect 8159 14056 8171 14059
rect 8570 14056 8576 14068
rect 8159 14028 8576 14056
rect 8159 14025 8171 14028
rect 8113 14019 8171 14025
rect 8570 14016 8576 14028
rect 8628 14016 8634 14068
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 10229 14059 10287 14065
rect 10229 14056 10241 14059
rect 9824 14028 10241 14056
rect 9824 14016 9830 14028
rect 10229 14025 10241 14028
rect 10275 14025 10287 14059
rect 10229 14019 10287 14025
rect 13814 14016 13820 14068
rect 13872 14056 13878 14068
rect 15102 14056 15108 14068
rect 13872 14028 15108 14056
rect 13872 14016 13878 14028
rect 15102 14016 15108 14028
rect 15160 14016 15166 14068
rect 17865 14059 17923 14065
rect 17865 14025 17877 14059
rect 17911 14056 17923 14059
rect 18141 14059 18199 14065
rect 18141 14056 18153 14059
rect 17911 14028 18153 14056
rect 17911 14025 17923 14028
rect 17865 14019 17923 14025
rect 18141 14025 18153 14028
rect 18187 14056 18199 14059
rect 18966 14056 18972 14068
rect 18187 14028 18972 14056
rect 18187 14025 18199 14028
rect 18141 14019 18199 14025
rect 18966 14016 18972 14028
rect 19024 14016 19030 14068
rect 5810 13948 5816 14000
rect 5868 13988 5874 14000
rect 6181 13991 6239 13997
rect 6181 13988 6193 13991
rect 5868 13960 6193 13988
rect 5868 13948 5874 13960
rect 6181 13957 6193 13960
rect 6227 13988 6239 13991
rect 7837 13991 7895 13997
rect 7837 13988 7849 13991
rect 6227 13960 7328 13988
rect 6227 13957 6239 13960
rect 6181 13951 6239 13957
rect 6733 13923 6791 13929
rect 6733 13889 6745 13923
rect 6779 13920 6791 13923
rect 7101 13923 7159 13929
rect 7101 13920 7113 13923
rect 6779 13892 7113 13920
rect 6779 13889 6791 13892
rect 6733 13883 6791 13889
rect 7101 13889 7113 13892
rect 7147 13889 7159 13923
rect 7101 13883 7159 13889
rect 5166 13812 5172 13864
rect 5224 13852 5230 13864
rect 6089 13855 6147 13861
rect 6089 13852 6101 13855
rect 5224 13824 6101 13852
rect 5224 13812 5230 13824
rect 6089 13821 6101 13824
rect 6135 13852 6147 13855
rect 6454 13852 6460 13864
rect 6135 13824 6460 13852
rect 6135 13821 6147 13824
rect 6089 13815 6147 13821
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 6638 13852 6644 13864
rect 6599 13824 6644 13852
rect 6638 13812 6644 13824
rect 6696 13812 6702 13864
rect 6822 13852 6828 13864
rect 6783 13824 6828 13852
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7300 13861 7328 13960
rect 7576 13960 7849 13988
rect 7576 13864 7604 13960
rect 7837 13957 7849 13960
rect 7883 13957 7895 13991
rect 9861 13991 9919 13997
rect 9861 13988 9873 13991
rect 7837 13951 7895 13957
rect 7944 13960 9873 13988
rect 7944 13920 7972 13960
rect 9861 13957 9873 13960
rect 9907 13957 9919 13991
rect 9861 13951 9919 13957
rect 17497 13991 17555 13997
rect 17497 13957 17509 13991
rect 17543 13988 17555 13991
rect 18046 13988 18052 14000
rect 17543 13960 18052 13988
rect 17543 13957 17555 13960
rect 17497 13951 17555 13957
rect 18046 13948 18052 13960
rect 18104 13948 18110 14000
rect 7760 13892 7972 13920
rect 6917 13855 6975 13861
rect 6917 13821 6929 13855
rect 6963 13821 6975 13855
rect 6917 13815 6975 13821
rect 7285 13855 7343 13861
rect 7285 13821 7297 13855
rect 7331 13821 7343 13855
rect 7285 13815 7343 13821
rect 7469 13855 7527 13861
rect 7469 13821 7481 13855
rect 7515 13852 7527 13855
rect 7558 13852 7564 13864
rect 7515 13824 7564 13852
rect 7515 13821 7527 13824
rect 7469 13815 7527 13821
rect 6730 13676 6736 13728
rect 6788 13716 6794 13728
rect 6932 13716 6960 13815
rect 7558 13812 7564 13824
rect 7616 13812 7622 13864
rect 7760 13861 7788 13892
rect 9582 13880 9588 13932
rect 9640 13920 9646 13932
rect 9769 13923 9827 13929
rect 9769 13920 9781 13923
rect 9640 13892 9781 13920
rect 9640 13880 9646 13892
rect 9769 13889 9781 13892
rect 9815 13889 9827 13923
rect 9769 13883 9827 13889
rect 17957 13923 18015 13929
rect 17957 13889 17969 13923
rect 18003 13889 18015 13923
rect 17957 13883 18015 13889
rect 7745 13855 7803 13861
rect 7745 13821 7757 13855
rect 7791 13821 7803 13855
rect 7745 13815 7803 13821
rect 7190 13744 7196 13796
rect 7248 13784 7254 13796
rect 7760 13784 7788 13815
rect 8018 13812 8024 13864
rect 8076 13852 8082 13864
rect 9490 13852 9496 13864
rect 8076 13824 8121 13852
rect 9451 13824 9496 13852
rect 8076 13812 8082 13824
rect 9490 13812 9496 13824
rect 9548 13812 9554 13864
rect 9677 13855 9735 13861
rect 9677 13821 9689 13855
rect 9723 13821 9735 13855
rect 9677 13815 9735 13821
rect 9953 13855 10011 13861
rect 9953 13821 9965 13855
rect 9999 13852 10011 13855
rect 10134 13852 10140 13864
rect 9999 13824 10140 13852
rect 9999 13821 10011 13824
rect 9953 13815 10011 13821
rect 7248 13756 7788 13784
rect 7248 13744 7254 13756
rect 7650 13716 7656 13728
rect 6788 13688 6960 13716
rect 7611 13688 7656 13716
rect 6788 13676 6794 13688
rect 7650 13676 7656 13688
rect 7708 13676 7714 13728
rect 8202 13676 8208 13728
rect 8260 13716 8266 13728
rect 9692 13716 9720 13815
rect 10134 13812 10140 13824
rect 10192 13812 10198 13864
rect 17773 13855 17831 13861
rect 17773 13821 17785 13855
rect 17819 13821 17831 13855
rect 17773 13815 17831 13821
rect 17788 13784 17816 13815
rect 17862 13812 17868 13864
rect 17920 13852 17926 13864
rect 17972 13852 18000 13883
rect 17920 13824 18000 13852
rect 18233 13855 18291 13861
rect 17920 13812 17926 13824
rect 18233 13821 18245 13855
rect 18279 13821 18291 13855
rect 18233 13815 18291 13821
rect 18785 13855 18843 13861
rect 18785 13821 18797 13855
rect 18831 13852 18843 13855
rect 19334 13852 19340 13864
rect 18831 13824 19340 13852
rect 18831 13821 18843 13824
rect 18785 13815 18843 13821
rect 18248 13784 18276 13815
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 18690 13784 18696 13796
rect 17788 13756 18696 13784
rect 18690 13744 18696 13756
rect 18748 13784 18754 13796
rect 18877 13787 18935 13793
rect 18877 13784 18889 13787
rect 18748 13756 18889 13784
rect 18748 13744 18754 13756
rect 18877 13753 18889 13756
rect 18923 13753 18935 13787
rect 18877 13747 18935 13753
rect 9858 13716 9864 13728
rect 8260 13688 9864 13716
rect 8260 13676 8266 13688
rect 9858 13676 9864 13688
rect 9916 13676 9922 13728
rect 17954 13716 17960 13728
rect 17915 13688 17960 13716
rect 17954 13676 17960 13688
rect 18012 13676 18018 13728
rect 1104 13626 21804 13648
rect 1104 13574 7882 13626
rect 7934 13574 7946 13626
rect 7998 13574 8010 13626
rect 8062 13574 8074 13626
rect 8126 13574 14782 13626
rect 14834 13574 14846 13626
rect 14898 13574 14910 13626
rect 14962 13574 14974 13626
rect 15026 13574 21804 13626
rect 1104 13552 21804 13574
rect 1578 13472 1584 13524
rect 1636 13512 1642 13524
rect 1857 13515 1915 13521
rect 1857 13512 1869 13515
rect 1636 13484 1869 13512
rect 1636 13472 1642 13484
rect 1857 13481 1869 13484
rect 1903 13481 1915 13515
rect 3326 13512 3332 13524
rect 3287 13484 3332 13512
rect 1857 13475 1915 13481
rect 3326 13472 3332 13484
rect 3384 13472 3390 13524
rect 7374 13512 7380 13524
rect 7335 13484 7380 13512
rect 7374 13472 7380 13484
rect 7432 13472 7438 13524
rect 8294 13512 8300 13524
rect 8255 13484 8300 13512
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 17773 13515 17831 13521
rect 17773 13512 17785 13515
rect 8404 13484 16160 13512
rect 5534 13404 5540 13456
rect 5592 13444 5598 13456
rect 8404 13444 8432 13484
rect 12066 13444 12072 13456
rect 5592 13416 8432 13444
rect 12027 13416 12072 13444
rect 5592 13404 5598 13416
rect 12066 13404 12072 13416
rect 12124 13404 12130 13456
rect 12161 13447 12219 13453
rect 12161 13413 12173 13447
rect 12207 13413 12219 13447
rect 12161 13407 12219 13413
rect 1949 13379 2007 13385
rect 1949 13345 1961 13379
rect 1995 13345 2007 13379
rect 1949 13339 2007 13345
rect 1762 13308 1768 13320
rect 1723 13280 1768 13308
rect 1762 13268 1768 13280
rect 1820 13268 1826 13320
rect 1964 13308 1992 13339
rect 3142 13336 3148 13388
rect 3200 13376 3206 13388
rect 3237 13379 3295 13385
rect 3237 13376 3249 13379
rect 3200 13348 3249 13376
rect 3200 13336 3206 13348
rect 3237 13345 3249 13348
rect 3283 13345 3295 13379
rect 3237 13339 3295 13345
rect 6638 13336 6644 13388
rect 6696 13376 6702 13388
rect 7285 13379 7343 13385
rect 7285 13376 7297 13379
rect 6696 13348 7297 13376
rect 6696 13336 6702 13348
rect 7285 13345 7297 13348
rect 7331 13345 7343 13379
rect 7285 13339 7343 13345
rect 4890 13308 4896 13320
rect 1964 13280 4896 13308
rect 4890 13268 4896 13280
rect 4948 13268 4954 13320
rect 7300 13308 7328 13339
rect 8110 13336 8116 13388
rect 8168 13376 8174 13388
rect 8205 13379 8263 13385
rect 8205 13376 8217 13379
rect 8168 13348 8217 13376
rect 8168 13336 8174 13348
rect 8205 13345 8217 13348
rect 8251 13376 8263 13379
rect 10962 13376 10968 13388
rect 8251 13348 10968 13376
rect 8251 13345 8263 13348
rect 8205 13339 8263 13345
rect 10962 13336 10968 13348
rect 11020 13336 11026 13388
rect 12176 13376 12204 13407
rect 14366 13404 14372 13456
rect 14424 13444 14430 13456
rect 14642 13444 14648 13456
rect 14424 13416 14648 13444
rect 14424 13404 14430 13416
rect 14642 13404 14648 13416
rect 14700 13404 14706 13456
rect 12802 13376 12808 13388
rect 11072 13348 12204 13376
rect 12763 13348 12808 13376
rect 10042 13308 10048 13320
rect 7300 13280 10048 13308
rect 10042 13268 10048 13280
rect 10100 13268 10106 13320
rect 11072 13308 11100 13348
rect 12802 13336 12808 13348
rect 12860 13336 12866 13388
rect 12989 13379 13047 13385
rect 12989 13345 13001 13379
rect 13035 13345 13047 13379
rect 12989 13339 13047 13345
rect 10152 13280 11100 13308
rect 4798 13200 4804 13252
rect 4856 13240 4862 13252
rect 10152 13240 10180 13280
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 13004 13308 13032 13339
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 14553 13379 14611 13385
rect 14553 13376 14565 13379
rect 13964 13348 14565 13376
rect 13964 13336 13970 13348
rect 14553 13345 14565 13348
rect 14599 13345 14611 13379
rect 14553 13339 14611 13345
rect 14737 13379 14795 13385
rect 14737 13345 14749 13379
rect 14783 13345 14795 13379
rect 14737 13339 14795 13345
rect 14921 13379 14979 13385
rect 14921 13345 14933 13379
rect 14967 13376 14979 13379
rect 15102 13376 15108 13388
rect 14967 13348 15108 13376
rect 14967 13345 14979 13348
rect 14921 13339 14979 13345
rect 12216 13280 12261 13308
rect 12406 13280 13032 13308
rect 14752 13308 14780 13339
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 15562 13308 15568 13320
rect 14752 13280 15568 13308
rect 12216 13268 12222 13280
rect 4856 13212 10180 13240
rect 4856 13200 4862 13212
rect 10410 13200 10416 13252
rect 10468 13240 10474 13252
rect 10870 13240 10876 13252
rect 10468 13212 10876 13240
rect 10468 13200 10474 13212
rect 10870 13200 10876 13212
rect 10928 13240 10934 13252
rect 12250 13240 12256 13252
rect 10928 13212 12256 13240
rect 10928 13200 10934 13212
rect 12250 13200 12256 13212
rect 12308 13240 12314 13252
rect 12406 13240 12434 13280
rect 15562 13268 15568 13280
rect 15620 13308 15626 13320
rect 15657 13311 15715 13317
rect 15657 13308 15669 13311
rect 15620 13280 15669 13308
rect 15620 13268 15626 13280
rect 15657 13277 15669 13280
rect 15703 13308 15715 13311
rect 16132 13308 16160 13484
rect 17420 13484 17785 13512
rect 16666 13404 16672 13456
rect 16724 13404 16730 13456
rect 17420 13453 17448 13484
rect 17773 13481 17785 13484
rect 17819 13481 17831 13515
rect 19429 13515 19487 13521
rect 19429 13512 19441 13515
rect 17773 13475 17831 13481
rect 18156 13484 19441 13512
rect 17405 13447 17463 13453
rect 17405 13413 17417 13447
rect 17451 13413 17463 13447
rect 17405 13407 17463 13413
rect 17678 13404 17684 13456
rect 17736 13444 17742 13456
rect 18156 13444 18184 13484
rect 19429 13481 19441 13484
rect 19475 13481 19487 13515
rect 19429 13475 19487 13481
rect 18966 13444 18972 13456
rect 17736 13416 18184 13444
rect 17736 13404 17742 13416
rect 18046 13376 18052 13388
rect 18007 13348 18052 13376
rect 18046 13336 18052 13348
rect 18104 13336 18110 13388
rect 18156 13385 18184 13416
rect 18892 13416 18972 13444
rect 18141 13379 18199 13385
rect 18141 13345 18153 13379
rect 18187 13345 18199 13379
rect 18690 13376 18696 13388
rect 18651 13348 18696 13376
rect 18141 13339 18199 13345
rect 18690 13336 18696 13348
rect 18748 13336 18754 13388
rect 18892 13385 18920 13416
rect 18966 13404 18972 13416
rect 19024 13404 19030 13456
rect 19334 13444 19340 13456
rect 19076 13416 19340 13444
rect 19076 13385 19104 13416
rect 19334 13404 19340 13416
rect 19392 13444 19398 13456
rect 19889 13447 19947 13453
rect 19392 13416 19840 13444
rect 19392 13404 19398 13416
rect 19812 13388 19840 13416
rect 19889 13413 19901 13447
rect 19935 13444 19947 13447
rect 20070 13444 20076 13456
rect 19935 13416 20076 13444
rect 19935 13413 19947 13416
rect 19889 13407 19947 13413
rect 20070 13404 20076 13416
rect 20128 13404 20134 13456
rect 18877 13379 18935 13385
rect 18877 13345 18889 13379
rect 18923 13345 18935 13379
rect 18877 13339 18935 13345
rect 19061 13379 19119 13385
rect 19061 13345 19073 13379
rect 19107 13345 19119 13379
rect 19061 13339 19119 13345
rect 19245 13379 19303 13385
rect 19245 13345 19257 13379
rect 19291 13376 19303 13379
rect 19429 13379 19487 13385
rect 19429 13376 19441 13379
rect 19291 13348 19441 13376
rect 19291 13345 19303 13348
rect 19245 13339 19303 13345
rect 19429 13345 19441 13348
rect 19475 13345 19487 13379
rect 19610 13376 19616 13388
rect 19571 13348 19616 13376
rect 19429 13339 19487 13345
rect 15703 13280 15976 13308
rect 16132 13280 17632 13308
rect 15703 13277 15715 13280
rect 15657 13271 15715 13277
rect 12308 13212 12434 13240
rect 12621 13243 12679 13249
rect 12308 13200 12314 13212
rect 12621 13209 12633 13243
rect 12667 13240 12679 13243
rect 13722 13240 13728 13252
rect 12667 13212 13728 13240
rect 12667 13209 12679 13212
rect 12621 13203 12679 13209
rect 13722 13200 13728 13212
rect 13780 13200 13786 13252
rect 2130 13132 2136 13184
rect 2188 13172 2194 13184
rect 2317 13175 2375 13181
rect 2317 13172 2329 13175
rect 2188 13144 2329 13172
rect 2188 13132 2194 13144
rect 2317 13141 2329 13144
rect 2363 13141 2375 13175
rect 2317 13135 2375 13141
rect 13173 13175 13231 13181
rect 13173 13141 13185 13175
rect 13219 13172 13231 13175
rect 13262 13172 13268 13184
rect 13219 13144 13268 13172
rect 13219 13141 13231 13144
rect 13173 13135 13231 13141
rect 13262 13132 13268 13144
rect 13320 13132 13326 13184
rect 14369 13175 14427 13181
rect 14369 13141 14381 13175
rect 14415 13172 14427 13175
rect 15838 13172 15844 13184
rect 14415 13144 15844 13172
rect 14415 13141 14427 13144
rect 14369 13135 14427 13141
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 15948 13172 15976 13280
rect 17604 13240 17632 13280
rect 17678 13268 17684 13320
rect 17736 13308 17742 13320
rect 17954 13308 17960 13320
rect 17736 13280 17781 13308
rect 17915 13280 17960 13308
rect 17736 13268 17742 13280
rect 17954 13268 17960 13280
rect 18012 13268 18018 13320
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13308 18291 13311
rect 18598 13308 18604 13320
rect 18279 13280 18604 13308
rect 18279 13277 18291 13280
rect 18233 13271 18291 13277
rect 18598 13268 18604 13280
rect 18656 13268 18662 13320
rect 18969 13311 19027 13317
rect 18969 13277 18981 13311
rect 19015 13308 19027 13311
rect 19150 13308 19156 13320
rect 19015 13280 19156 13308
rect 19015 13277 19027 13280
rect 18969 13271 19027 13277
rect 19150 13268 19156 13280
rect 19208 13268 19214 13320
rect 19444 13308 19472 13339
rect 19610 13336 19616 13348
rect 19668 13336 19674 13388
rect 19794 13376 19800 13388
rect 19755 13348 19800 13376
rect 19794 13336 19800 13348
rect 19852 13336 19858 13388
rect 19981 13379 20039 13385
rect 19981 13345 19993 13379
rect 20027 13345 20039 13379
rect 19981 13339 20039 13345
rect 19996 13308 20024 13339
rect 20438 13336 20444 13388
rect 20496 13376 20502 13388
rect 20625 13379 20683 13385
rect 20625 13376 20637 13379
rect 20496 13348 20637 13376
rect 20496 13336 20502 13348
rect 20625 13345 20637 13348
rect 20671 13345 20683 13379
rect 21450 13376 21456 13388
rect 21411 13348 21456 13376
rect 20625 13339 20683 13345
rect 21450 13336 21456 13348
rect 21508 13336 21514 13388
rect 19444 13280 20024 13308
rect 21269 13243 21327 13249
rect 21269 13240 21281 13243
rect 17604 13212 21281 13240
rect 21269 13209 21281 13212
rect 21315 13209 21327 13243
rect 21269 13203 21327 13209
rect 17310 13172 17316 13184
rect 15948 13144 17316 13172
rect 17310 13132 17316 13144
rect 17368 13132 17374 13184
rect 18509 13175 18567 13181
rect 18509 13141 18521 13175
rect 18555 13172 18567 13175
rect 18874 13172 18880 13184
rect 18555 13144 18880 13172
rect 18555 13141 18567 13144
rect 18509 13135 18567 13141
rect 18874 13132 18880 13144
rect 18932 13132 18938 13184
rect 19978 13132 19984 13184
rect 20036 13172 20042 13184
rect 20165 13175 20223 13181
rect 20165 13172 20177 13175
rect 20036 13144 20177 13172
rect 20036 13132 20042 13144
rect 20165 13141 20177 13144
rect 20211 13141 20223 13175
rect 20165 13135 20223 13141
rect 20714 13132 20720 13184
rect 20772 13172 20778 13184
rect 20809 13175 20867 13181
rect 20809 13172 20821 13175
rect 20772 13144 20821 13172
rect 20772 13132 20778 13144
rect 20809 13141 20821 13144
rect 20855 13141 20867 13175
rect 20809 13135 20867 13141
rect 1104 13082 21804 13104
rect 1104 13030 4432 13082
rect 4484 13030 4496 13082
rect 4548 13030 4560 13082
rect 4612 13030 4624 13082
rect 4676 13030 11332 13082
rect 11384 13030 11396 13082
rect 11448 13030 11460 13082
rect 11512 13030 11524 13082
rect 11576 13030 18232 13082
rect 18284 13030 18296 13082
rect 18348 13030 18360 13082
rect 18412 13030 18424 13082
rect 18476 13030 21804 13082
rect 1104 13008 21804 13030
rect 1486 12968 1492 12980
rect 1447 12940 1492 12968
rect 1486 12928 1492 12940
rect 1544 12928 1550 12980
rect 2685 12971 2743 12977
rect 2685 12937 2697 12971
rect 2731 12968 2743 12971
rect 3142 12968 3148 12980
rect 2731 12940 3148 12968
rect 2731 12937 2743 12940
rect 2685 12931 2743 12937
rect 3142 12928 3148 12940
rect 3200 12928 3206 12980
rect 4890 12968 4896 12980
rect 4851 12940 4896 12968
rect 4890 12928 4896 12940
rect 4948 12928 4954 12980
rect 5258 12968 5264 12980
rect 5171 12940 5264 12968
rect 5258 12928 5264 12940
rect 5316 12968 5322 12980
rect 6178 12968 6184 12980
rect 5316 12940 6184 12968
rect 5316 12928 5322 12940
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 6638 12928 6644 12980
rect 6696 12968 6702 12980
rect 6733 12971 6791 12977
rect 6733 12968 6745 12971
rect 6696 12940 6745 12968
rect 6696 12928 6702 12940
rect 6733 12937 6745 12940
rect 6779 12937 6791 12971
rect 6733 12931 6791 12937
rect 8662 12928 8668 12980
rect 8720 12968 8726 12980
rect 9217 12971 9275 12977
rect 9217 12968 9229 12971
rect 8720 12940 9229 12968
rect 8720 12928 8726 12940
rect 9217 12937 9229 12940
rect 9263 12937 9275 12971
rect 9858 12968 9864 12980
rect 9819 12940 9864 12968
rect 9217 12931 9275 12937
rect 9858 12928 9864 12940
rect 9916 12928 9922 12980
rect 10042 12968 10048 12980
rect 10003 12940 10048 12968
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 12066 12928 12072 12980
rect 12124 12968 12130 12980
rect 16577 12971 16635 12977
rect 12124 12940 13492 12968
rect 12124 12928 12130 12940
rect 9582 12900 9588 12912
rect 8496 12872 9588 12900
rect 2777 12835 2835 12841
rect 2777 12832 2789 12835
rect 2148 12804 2789 12832
rect 2148 12776 2176 12804
rect 2777 12801 2789 12804
rect 2823 12801 2835 12835
rect 5350 12832 5356 12844
rect 2777 12795 2835 12801
rect 5276 12804 5356 12832
rect 2130 12764 2136 12776
rect 2091 12736 2136 12764
rect 2130 12724 2136 12736
rect 2188 12724 2194 12776
rect 2685 12767 2743 12773
rect 2685 12733 2697 12767
rect 2731 12764 2743 12767
rect 2958 12764 2964 12776
rect 2731 12736 2964 12764
rect 2731 12733 2743 12736
rect 2685 12727 2743 12733
rect 2958 12724 2964 12736
rect 3016 12724 3022 12776
rect 3145 12767 3203 12773
rect 3145 12733 3157 12767
rect 3191 12764 3203 12767
rect 3326 12764 3332 12776
rect 3191 12736 3332 12764
rect 3191 12733 3203 12736
rect 3145 12727 3203 12733
rect 3326 12724 3332 12736
rect 3384 12724 3390 12776
rect 5166 12764 5172 12776
rect 5127 12736 5172 12764
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 5276 12773 5304 12804
rect 5350 12792 5356 12804
rect 5408 12832 5414 12844
rect 8110 12832 8116 12844
rect 5408 12804 8116 12832
rect 5408 12792 5414 12804
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 8496 12776 8524 12872
rect 9582 12860 9588 12872
rect 9640 12900 9646 12912
rect 9953 12903 10011 12909
rect 9953 12900 9965 12903
rect 9640 12872 9965 12900
rect 9640 12860 9646 12872
rect 9953 12869 9965 12872
rect 9999 12869 10011 12903
rect 10060 12900 10088 12928
rect 11238 12900 11244 12912
rect 10060 12872 11244 12900
rect 9953 12863 10011 12869
rect 9309 12835 9367 12841
rect 9309 12801 9321 12835
rect 9355 12832 9367 12835
rect 9490 12832 9496 12844
rect 9355 12804 9496 12832
rect 9355 12801 9367 12804
rect 9309 12795 9367 12801
rect 9490 12792 9496 12804
rect 9548 12832 9554 12844
rect 9968 12832 9996 12863
rect 11238 12860 11244 12872
rect 11296 12860 11302 12912
rect 11425 12903 11483 12909
rect 11425 12869 11437 12903
rect 11471 12900 11483 12903
rect 12802 12900 12808 12912
rect 11471 12872 12808 12900
rect 11471 12869 11483 12872
rect 11425 12863 11483 12869
rect 12176 12841 12204 12872
rect 12802 12860 12808 12872
rect 12860 12860 12866 12912
rect 10413 12835 10471 12841
rect 9548 12804 9720 12832
rect 9968 12804 10272 12832
rect 9548 12792 9554 12804
rect 5261 12767 5319 12773
rect 5261 12733 5273 12767
rect 5307 12733 5319 12767
rect 6454 12764 6460 12776
rect 6415 12736 6460 12764
rect 5261 12727 5319 12733
rect 6454 12724 6460 12736
rect 6512 12724 6518 12776
rect 7742 12764 7748 12776
rect 7703 12736 7748 12764
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 8294 12764 8300 12776
rect 8255 12736 8300 12764
rect 8294 12724 8300 12736
rect 8352 12724 8358 12776
rect 8478 12764 8484 12776
rect 8439 12736 8484 12764
rect 8478 12724 8484 12736
rect 8536 12724 8542 12776
rect 9692 12773 9720 12804
rect 9217 12767 9275 12773
rect 9217 12733 9229 12767
rect 9263 12733 9275 12767
rect 9217 12727 9275 12733
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12733 9735 12767
rect 10134 12764 10140 12776
rect 10095 12736 10140 12764
rect 9677 12727 9735 12733
rect 1581 12699 1639 12705
rect 1581 12665 1593 12699
rect 1627 12696 1639 12699
rect 3234 12696 3240 12708
rect 1627 12668 3240 12696
rect 1627 12665 1639 12668
rect 1581 12659 1639 12665
rect 3234 12656 3240 12668
rect 3292 12656 3298 12708
rect 6178 12656 6184 12708
rect 6236 12696 6242 12708
rect 6641 12699 6699 12705
rect 6641 12696 6653 12699
rect 6236 12668 6653 12696
rect 6236 12656 6242 12668
rect 6641 12665 6653 12668
rect 6687 12696 6699 12699
rect 7190 12696 7196 12708
rect 6687 12668 7196 12696
rect 6687 12665 6699 12668
rect 6641 12659 6699 12665
rect 7190 12656 7196 12668
rect 7248 12656 7254 12708
rect 7466 12656 7472 12708
rect 7524 12696 7530 12708
rect 7561 12699 7619 12705
rect 7561 12696 7573 12699
rect 7524 12668 7573 12696
rect 7524 12656 7530 12668
rect 7561 12665 7573 12668
rect 7607 12665 7619 12699
rect 7561 12659 7619 12665
rect 7650 12656 7656 12708
rect 7708 12696 7714 12708
rect 9232 12696 9260 12727
rect 10134 12724 10140 12736
rect 10192 12724 10198 12776
rect 10244 12764 10272 12804
rect 10413 12801 10425 12835
rect 10459 12832 10471 12835
rect 12161 12835 12219 12841
rect 10459 12804 12112 12832
rect 10459 12801 10471 12804
rect 10413 12795 10471 12801
rect 10781 12767 10839 12773
rect 10781 12764 10793 12767
rect 10244 12736 10793 12764
rect 10781 12733 10793 12736
rect 10827 12733 10839 12767
rect 10781 12727 10839 12733
rect 10965 12767 11023 12773
rect 10965 12733 10977 12767
rect 11011 12764 11023 12767
rect 12084 12764 12112 12804
rect 12161 12801 12173 12835
rect 12207 12801 12219 12835
rect 12161 12795 12219 12801
rect 12250 12792 12256 12844
rect 12308 12832 12314 12844
rect 13464 12841 13492 12940
rect 16577 12937 16589 12971
rect 16623 12968 16635 12971
rect 16666 12968 16672 12980
rect 16623 12940 16672 12968
rect 16623 12937 16635 12940
rect 16577 12931 16635 12937
rect 16666 12928 16672 12940
rect 16724 12928 16730 12980
rect 17405 12971 17463 12977
rect 17405 12937 17417 12971
rect 17451 12968 17463 12971
rect 17862 12968 17868 12980
rect 17451 12940 17868 12968
rect 17451 12937 17463 12940
rect 17405 12931 17463 12937
rect 17862 12928 17868 12940
rect 17920 12928 17926 12980
rect 20070 12928 20076 12980
rect 20128 12968 20134 12980
rect 21453 12971 21511 12977
rect 21453 12968 21465 12971
rect 20128 12940 21465 12968
rect 20128 12928 20134 12940
rect 21453 12937 21465 12940
rect 21499 12937 21511 12971
rect 21453 12931 21511 12937
rect 16758 12900 16764 12912
rect 13556 12872 16764 12900
rect 13449 12835 13507 12841
rect 12308 12804 12353 12832
rect 12308 12792 12314 12804
rect 13449 12801 13461 12835
rect 13495 12801 13507 12835
rect 13449 12795 13507 12801
rect 13262 12764 13268 12776
rect 11011 12736 11836 12764
rect 12084 12736 12434 12764
rect 13223 12736 13268 12764
rect 11011 12733 11023 12736
rect 10965 12727 11023 12733
rect 9490 12696 9496 12708
rect 7708 12668 9496 12696
rect 7708 12656 7714 12668
rect 9490 12656 9496 12668
rect 9548 12656 9554 12708
rect 10980 12696 11008 12727
rect 9600 12668 11008 12696
rect 8481 12631 8539 12637
rect 8481 12597 8493 12631
rect 8527 12628 8539 12631
rect 9122 12628 9128 12640
rect 8527 12600 9128 12628
rect 8527 12597 8539 12600
rect 8481 12591 8539 12597
rect 9122 12588 9128 12600
rect 9180 12588 9186 12640
rect 9600 12637 9628 12668
rect 11054 12656 11060 12708
rect 11112 12696 11118 12708
rect 11238 12696 11244 12708
rect 11112 12668 11157 12696
rect 11199 12668 11244 12696
rect 11112 12656 11118 12668
rect 11238 12656 11244 12668
rect 11296 12656 11302 12708
rect 9585 12631 9643 12637
rect 9585 12597 9597 12631
rect 9631 12597 9643 12631
rect 9585 12591 9643 12597
rect 10873 12631 10931 12637
rect 10873 12597 10885 12631
rect 10919 12628 10931 12631
rect 11330 12628 11336 12640
rect 10919 12600 11336 12628
rect 10919 12597 10931 12600
rect 10873 12591 10931 12597
rect 11330 12588 11336 12600
rect 11388 12588 11394 12640
rect 11698 12628 11704 12640
rect 11659 12600 11704 12628
rect 11698 12588 11704 12600
rect 11756 12588 11762 12640
rect 11808 12628 11836 12736
rect 12406 12696 12434 12736
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 13357 12767 13415 12773
rect 13357 12733 13369 12767
rect 13403 12764 13415 12767
rect 13556 12764 13584 12872
rect 16758 12860 16764 12872
rect 16816 12860 16822 12912
rect 19334 12900 19340 12912
rect 16868 12872 19340 12900
rect 13403 12736 13584 12764
rect 14737 12767 14795 12773
rect 13403 12733 13415 12736
rect 13357 12727 13415 12733
rect 14737 12733 14749 12767
rect 14783 12764 14795 12767
rect 16761 12767 16819 12773
rect 16761 12764 16773 12767
rect 14783 12736 16773 12764
rect 14783 12733 14795 12736
rect 14737 12727 14795 12733
rect 16761 12733 16773 12736
rect 16807 12764 16819 12767
rect 16868 12764 16896 12872
rect 19334 12860 19340 12872
rect 19392 12860 19398 12912
rect 17678 12792 17684 12844
rect 17736 12832 17742 12844
rect 19150 12832 19156 12844
rect 17736 12804 19156 12832
rect 17736 12792 17742 12804
rect 19150 12792 19156 12804
rect 19208 12832 19214 12844
rect 19705 12835 19763 12841
rect 19705 12832 19717 12835
rect 19208 12804 19717 12832
rect 19208 12792 19214 12804
rect 19705 12801 19717 12804
rect 19751 12801 19763 12835
rect 19978 12832 19984 12844
rect 19939 12804 19984 12832
rect 19705 12795 19763 12801
rect 19978 12792 19984 12804
rect 20036 12792 20042 12844
rect 17310 12764 17316 12776
rect 16807 12736 16896 12764
rect 17271 12736 17316 12764
rect 16807 12733 16819 12736
rect 16761 12727 16819 12733
rect 17310 12724 17316 12736
rect 17368 12724 17374 12776
rect 18874 12764 18880 12776
rect 18835 12736 18880 12764
rect 18874 12724 18880 12736
rect 18932 12724 18938 12776
rect 17954 12696 17960 12708
rect 12406 12668 17960 12696
rect 17954 12656 17960 12668
rect 18012 12656 18018 12708
rect 18598 12656 18604 12708
rect 18656 12696 18662 12708
rect 19061 12699 19119 12705
rect 19061 12696 19073 12699
rect 18656 12668 19073 12696
rect 18656 12656 18662 12668
rect 19061 12665 19073 12668
rect 19107 12665 19119 12699
rect 19061 12659 19119 12665
rect 20714 12656 20720 12708
rect 20772 12656 20778 12708
rect 12069 12631 12127 12637
rect 12069 12628 12081 12631
rect 11808 12600 12081 12628
rect 12069 12597 12081 12600
rect 12115 12597 12127 12631
rect 12894 12628 12900 12640
rect 12855 12600 12900 12628
rect 12069 12591 12127 12597
rect 12894 12588 12900 12600
rect 12952 12588 12958 12640
rect 14921 12631 14979 12637
rect 14921 12597 14933 12631
rect 14967 12628 14979 12631
rect 15102 12628 15108 12640
rect 14967 12600 15108 12628
rect 14967 12597 14979 12600
rect 14921 12591 14979 12597
rect 15102 12588 15108 12600
rect 15160 12588 15166 12640
rect 19242 12628 19248 12640
rect 19203 12600 19248 12628
rect 19242 12588 19248 12600
rect 19300 12588 19306 12640
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 20346 12628 20352 12640
rect 19392 12600 20352 12628
rect 19392 12588 19398 12600
rect 20346 12588 20352 12600
rect 20404 12588 20410 12640
rect 1104 12538 21804 12560
rect 1104 12486 7882 12538
rect 7934 12486 7946 12538
rect 7998 12486 8010 12538
rect 8062 12486 8074 12538
rect 8126 12486 14782 12538
rect 14834 12486 14846 12538
rect 14898 12486 14910 12538
rect 14962 12486 14974 12538
rect 15026 12486 21804 12538
rect 1104 12464 21804 12486
rect 5166 12384 5172 12436
rect 5224 12384 5230 12436
rect 5534 12424 5540 12436
rect 5495 12396 5540 12424
rect 5534 12384 5540 12396
rect 5592 12384 5598 12436
rect 6730 12424 6736 12436
rect 5644 12396 6736 12424
rect 3326 12356 3332 12368
rect 3287 12328 3332 12356
rect 3326 12316 3332 12328
rect 3384 12316 3390 12368
rect 4798 12316 4804 12368
rect 4856 12356 4862 12368
rect 5184 12356 5212 12384
rect 5644 12356 5672 12396
rect 6730 12384 6736 12396
rect 6788 12424 6794 12436
rect 10318 12424 10324 12436
rect 6788 12396 10324 12424
rect 6788 12384 6794 12396
rect 10318 12384 10324 12396
rect 10376 12384 10382 12436
rect 11977 12427 12035 12433
rect 11977 12393 11989 12427
rect 12023 12424 12035 12427
rect 12158 12424 12164 12436
rect 12023 12396 12164 12424
rect 12023 12393 12035 12396
rect 11977 12387 12035 12393
rect 12158 12384 12164 12396
rect 12216 12384 12222 12436
rect 14366 12424 14372 12436
rect 14327 12396 14372 12424
rect 14366 12384 14372 12396
rect 14424 12384 14430 12436
rect 7466 12356 7472 12368
rect 4856 12328 5672 12356
rect 6012 12328 7472 12356
rect 4856 12316 4862 12328
rect 3510 12288 3516 12300
rect 3471 12260 3516 12288
rect 3510 12248 3516 12260
rect 3568 12248 3574 12300
rect 5166 12248 5172 12300
rect 5224 12288 5230 12300
rect 5629 12291 5687 12297
rect 5629 12288 5641 12291
rect 5224 12260 5641 12288
rect 5224 12248 5230 12260
rect 5629 12257 5641 12260
rect 5675 12257 5687 12291
rect 5629 12251 5687 12257
rect 5810 12248 5816 12300
rect 5868 12288 5874 12300
rect 6012 12297 6040 12328
rect 7466 12316 7472 12328
rect 7524 12316 7530 12368
rect 11330 12316 11336 12368
rect 11388 12356 11394 12368
rect 11388 12328 11836 12356
rect 11388 12316 11394 12328
rect 11808 12300 11836 12328
rect 15102 12316 15108 12368
rect 15160 12316 15166 12368
rect 15838 12356 15844 12368
rect 15799 12328 15844 12356
rect 15838 12316 15844 12328
rect 15896 12316 15902 12368
rect 5997 12291 6055 12297
rect 5997 12288 6009 12291
rect 5868 12260 6009 12288
rect 5868 12248 5874 12260
rect 5997 12257 6009 12260
rect 6043 12257 6055 12291
rect 5997 12251 6055 12257
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12288 6331 12291
rect 6638 12288 6644 12300
rect 6319 12260 6644 12288
rect 6319 12257 6331 12260
rect 6273 12251 6331 12257
rect 6638 12248 6644 12260
rect 6696 12248 6702 12300
rect 11698 12288 11704 12300
rect 11659 12260 11704 12288
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 11790 12248 11796 12300
rect 11848 12288 11854 12300
rect 16117 12291 16175 12297
rect 11848 12260 11893 12288
rect 11848 12248 11854 12260
rect 16117 12257 16129 12291
rect 16163 12288 16175 12291
rect 17678 12288 17684 12300
rect 16163 12260 17684 12288
rect 16163 12257 16175 12260
rect 16117 12251 16175 12257
rect 17678 12248 17684 12260
rect 17736 12248 17742 12300
rect 5537 12223 5595 12229
rect 5537 12189 5549 12223
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 6089 12223 6147 12229
rect 6089 12189 6101 12223
rect 6135 12189 6147 12223
rect 6089 12183 6147 12189
rect 5552 12152 5580 12183
rect 5813 12155 5871 12161
rect 5813 12152 5825 12155
rect 5552 12124 5825 12152
rect 5813 12121 5825 12124
rect 5859 12121 5871 12155
rect 6104 12152 6132 12183
rect 6178 12180 6184 12232
rect 6236 12220 6242 12232
rect 6236 12192 6281 12220
rect 6236 12180 6242 12192
rect 6454 12152 6460 12164
rect 6104 12124 6460 12152
rect 5813 12115 5871 12121
rect 6454 12112 6460 12124
rect 6512 12112 6518 12164
rect 5077 12087 5135 12093
rect 5077 12053 5089 12087
rect 5123 12084 5135 12087
rect 5258 12084 5264 12096
rect 5123 12056 5264 12084
rect 5123 12053 5135 12056
rect 5077 12047 5135 12053
rect 5258 12044 5264 12056
rect 5316 12044 5322 12096
rect 1104 11994 21804 12016
rect 1104 11942 4432 11994
rect 4484 11942 4496 11994
rect 4548 11942 4560 11994
rect 4612 11942 4624 11994
rect 4676 11942 11332 11994
rect 11384 11942 11396 11994
rect 11448 11942 11460 11994
rect 11512 11942 11524 11994
rect 11576 11942 18232 11994
rect 18284 11942 18296 11994
rect 18348 11942 18360 11994
rect 18412 11942 18424 11994
rect 18476 11942 21804 11994
rect 1104 11920 21804 11942
rect 10134 11840 10140 11892
rect 10192 11880 10198 11892
rect 10502 11880 10508 11892
rect 10192 11852 10508 11880
rect 10192 11840 10198 11852
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 6822 11812 6828 11824
rect 5920 11784 6828 11812
rect 5629 11747 5687 11753
rect 5629 11744 5641 11747
rect 5552 11716 5641 11744
rect 5552 11608 5580 11716
rect 5629 11713 5641 11716
rect 5675 11713 5687 11747
rect 5810 11744 5816 11756
rect 5771 11716 5816 11744
rect 5629 11707 5687 11713
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 5920 11753 5948 11784
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 7742 11772 7748 11824
rect 7800 11812 7806 11824
rect 9401 11815 9459 11821
rect 9401 11812 9413 11815
rect 7800 11784 9413 11812
rect 7800 11772 7806 11784
rect 5905 11747 5963 11753
rect 5905 11713 5917 11747
rect 5951 11713 5963 11747
rect 5905 11707 5963 11713
rect 6457 11747 6515 11753
rect 6457 11713 6469 11747
rect 6503 11744 6515 11747
rect 6638 11744 6644 11756
rect 6503 11716 6644 11744
rect 6503 11713 6515 11716
rect 6457 11707 6515 11713
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 7760 11744 7788 11772
rect 8036 11753 8064 11784
rect 9401 11781 9413 11784
rect 9447 11781 9459 11815
rect 9401 11775 9459 11781
rect 6840 11716 7788 11744
rect 8021 11747 8079 11753
rect 5718 11676 5724 11688
rect 5679 11648 5724 11676
rect 5718 11636 5724 11648
rect 5776 11676 5782 11688
rect 6178 11676 6184 11688
rect 5776 11648 6184 11676
rect 5776 11636 5782 11648
rect 6178 11636 6184 11648
rect 6236 11636 6242 11688
rect 6840 11685 6868 11716
rect 8021 11713 8033 11747
rect 8067 11744 8079 11747
rect 8205 11747 8263 11753
rect 8067 11716 8101 11744
rect 8067 11713 8079 11716
rect 8021 11707 8079 11713
rect 8205 11713 8217 11747
rect 8251 11744 8263 11747
rect 8478 11744 8484 11756
rect 8251 11716 8484 11744
rect 8251 11713 8263 11716
rect 8205 11707 8263 11713
rect 8478 11704 8484 11716
rect 8536 11744 8542 11756
rect 8536 11716 9628 11744
rect 8536 11704 8542 11716
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6288 11648 6837 11676
rect 6288 11608 6316 11648
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 7742 11636 7748 11688
rect 7800 11676 7806 11688
rect 7929 11679 7987 11685
rect 7929 11676 7941 11679
rect 7800 11648 7941 11676
rect 7800 11636 7806 11648
rect 7929 11645 7941 11648
rect 7975 11645 7987 11679
rect 7929 11639 7987 11645
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11676 8171 11679
rect 8662 11676 8668 11688
rect 8159 11648 8668 11676
rect 8159 11645 8171 11648
rect 8113 11639 8171 11645
rect 8662 11636 8668 11648
rect 8720 11676 8726 11688
rect 9600 11685 9628 11716
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 10137 11747 10195 11753
rect 10137 11744 10149 11747
rect 10100 11716 10149 11744
rect 10100 11704 10106 11716
rect 10137 11713 10149 11716
rect 10183 11713 10195 11747
rect 10137 11707 10195 11713
rect 9309 11679 9367 11685
rect 9309 11676 9321 11679
rect 8720 11648 9321 11676
rect 8720 11636 8726 11648
rect 9309 11645 9321 11648
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 10229 11679 10287 11685
rect 10229 11645 10241 11679
rect 10275 11645 10287 11679
rect 10229 11639 10287 11645
rect 10413 11679 10471 11685
rect 10413 11645 10425 11679
rect 10459 11645 10471 11679
rect 10413 11639 10471 11645
rect 5552 11580 6316 11608
rect 6641 11611 6699 11617
rect 6641 11577 6653 11611
rect 6687 11608 6699 11611
rect 10042 11608 10048 11620
rect 6687 11580 6868 11608
rect 10003 11580 10048 11608
rect 6687 11577 6699 11580
rect 6641 11571 6699 11577
rect 6840 11552 6868 11580
rect 10042 11568 10048 11580
rect 10100 11608 10106 11620
rect 10244 11608 10272 11639
rect 10100 11580 10272 11608
rect 10100 11568 10106 11580
rect 4982 11500 4988 11552
rect 5040 11540 5046 11552
rect 5445 11543 5503 11549
rect 5445 11540 5457 11543
rect 5040 11512 5457 11540
rect 5040 11500 5046 11512
rect 5445 11509 5457 11512
rect 5491 11509 5503 11543
rect 5445 11503 5503 11509
rect 6822 11500 6828 11552
rect 6880 11500 6886 11552
rect 8202 11500 8208 11552
rect 8260 11540 8266 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 8260 11512 8401 11540
rect 8260 11500 8266 11512
rect 8389 11509 8401 11512
rect 8435 11509 8447 11543
rect 8389 11503 8447 11509
rect 9122 11500 9128 11552
rect 9180 11540 9186 11552
rect 10428 11540 10456 11639
rect 9180 11512 10456 11540
rect 10597 11543 10655 11549
rect 9180 11500 9186 11512
rect 10597 11509 10609 11543
rect 10643 11540 10655 11543
rect 18414 11540 18420 11552
rect 10643 11512 18420 11540
rect 10643 11509 10655 11512
rect 10597 11503 10655 11509
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 1104 11450 21804 11472
rect 1104 11398 7882 11450
rect 7934 11398 7946 11450
rect 7998 11398 8010 11450
rect 8062 11398 8074 11450
rect 8126 11398 14782 11450
rect 14834 11398 14846 11450
rect 14898 11398 14910 11450
rect 14962 11398 14974 11450
rect 15026 11398 21804 11450
rect 1104 11376 21804 11398
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 3510 11336 3516 11348
rect 3068 11308 3516 11336
rect 3068 11277 3096 11308
rect 3510 11296 3516 11308
rect 3568 11336 3574 11348
rect 4249 11339 4307 11345
rect 4249 11336 4261 11339
rect 3568 11308 4261 11336
rect 3568 11296 3574 11308
rect 4249 11305 4261 11308
rect 4295 11305 4307 11339
rect 4249 11299 4307 11305
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 7558 11336 7564 11348
rect 7248 11308 7564 11336
rect 7248 11296 7254 11308
rect 7558 11296 7564 11308
rect 7616 11336 7622 11348
rect 10413 11339 10471 11345
rect 7616 11308 8432 11336
rect 7616 11296 7622 11308
rect 3053 11271 3111 11277
rect 3053 11237 3065 11271
rect 3099 11237 3111 11271
rect 7009 11271 7067 11277
rect 3053 11231 3111 11237
rect 3436 11240 4568 11268
rect 1949 11203 2007 11209
rect 1949 11169 1961 11203
rect 1995 11169 2007 11203
rect 2958 11200 2964 11212
rect 2919 11172 2964 11200
rect 1949 11163 2007 11169
rect 1762 11132 1768 11144
rect 1723 11104 1768 11132
rect 1762 11092 1768 11104
rect 1820 11092 1826 11144
rect 1964 11132 1992 11163
rect 2958 11160 2964 11172
rect 3016 11200 3022 11212
rect 3436 11200 3464 11240
rect 4540 11209 4568 11240
rect 7009 11237 7021 11271
rect 7055 11268 7067 11271
rect 8113 11271 8171 11277
rect 7055 11240 7788 11268
rect 7055 11237 7067 11240
rect 7009 11231 7067 11237
rect 3016 11172 3464 11200
rect 3513 11203 3571 11209
rect 3016 11160 3022 11172
rect 3513 11169 3525 11203
rect 3559 11200 3571 11203
rect 4525 11203 4583 11209
rect 3559 11172 3924 11200
rect 3559 11169 3571 11172
rect 3513 11163 3571 11169
rect 3896 11141 3924 11172
rect 4525 11169 4537 11203
rect 4571 11169 4583 11203
rect 4525 11163 4583 11169
rect 6638 11160 6644 11212
rect 6696 11200 6702 11212
rect 6917 11203 6975 11209
rect 6917 11200 6929 11203
rect 6696 11172 6929 11200
rect 6696 11160 6702 11172
rect 6917 11169 6929 11172
rect 6963 11169 6975 11203
rect 7190 11200 7196 11212
rect 7151 11172 7196 11200
rect 6917 11163 6975 11169
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7300 11209 7328 11240
rect 7760 11212 7788 11240
rect 8113 11237 8125 11271
rect 8159 11268 8171 11271
rect 8202 11268 8208 11280
rect 8159 11240 8208 11268
rect 8159 11237 8171 11240
rect 8113 11231 8171 11237
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 7374 11160 7380 11212
rect 7432 11200 7438 11212
rect 7561 11203 7619 11209
rect 7561 11200 7573 11203
rect 7432 11172 7573 11200
rect 7432 11160 7438 11172
rect 7561 11169 7573 11172
rect 7607 11169 7619 11203
rect 7742 11200 7748 11212
rect 7703 11172 7748 11200
rect 7561 11163 7619 11169
rect 7742 11160 7748 11172
rect 7800 11200 7806 11212
rect 8404 11209 8432 11308
rect 10413 11305 10425 11339
rect 10459 11336 10471 11339
rect 10502 11336 10508 11348
rect 10459 11308 10508 11336
rect 10459 11305 10471 11308
rect 10413 11299 10471 11305
rect 10502 11296 10508 11308
rect 10560 11296 10566 11348
rect 11793 11339 11851 11345
rect 11793 11305 11805 11339
rect 11839 11336 11851 11339
rect 18414 11336 18420 11348
rect 11839 11308 18276 11336
rect 18375 11308 18420 11336
rect 11839 11305 11851 11308
rect 11793 11299 11851 11305
rect 10045 11271 10103 11277
rect 10045 11237 10057 11271
rect 10091 11237 10103 11271
rect 10045 11231 10103 11237
rect 8389 11203 8447 11209
rect 7800 11172 8248 11200
rect 7800 11160 7806 11172
rect 3881 11135 3939 11141
rect 1964 11104 2774 11132
rect 2317 11067 2375 11073
rect 2317 11033 2329 11067
rect 2363 11064 2375 11067
rect 2406 11064 2412 11076
rect 2363 11036 2412 11064
rect 2363 11033 2375 11036
rect 2317 11027 2375 11033
rect 2406 11024 2412 11036
rect 2464 11024 2470 11076
rect 2746 11064 2774 11104
rect 3881 11101 3893 11135
rect 3927 11132 3939 11135
rect 7469 11135 7527 11141
rect 3927 11104 7236 11132
rect 3927 11101 3939 11104
rect 3881 11095 3939 11101
rect 4154 11064 4160 11076
rect 2746 11036 4160 11064
rect 4154 11024 4160 11036
rect 4212 11024 4218 11076
rect 4249 11067 4307 11073
rect 4249 11033 4261 11067
rect 4295 11064 4307 11067
rect 4341 11067 4399 11073
rect 4341 11064 4353 11067
rect 4295 11036 4353 11064
rect 4295 11033 4307 11036
rect 4249 11027 4307 11033
rect 4341 11033 4353 11036
rect 4387 11033 4399 11067
rect 4341 11027 4399 11033
rect 7208 10996 7236 11104
rect 7469 11101 7481 11135
rect 7515 11132 7527 11135
rect 8110 11132 8116 11144
rect 7515 11104 8116 11132
rect 7515 11101 7527 11104
rect 7469 11095 7527 11101
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 8220 11141 8248 11172
rect 8389 11169 8401 11203
rect 8435 11169 8447 11203
rect 8389 11163 8447 11169
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11200 8539 11203
rect 8662 11200 8668 11212
rect 8527 11172 8668 11200
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 8662 11160 8668 11172
rect 8720 11160 8726 11212
rect 10060 11200 10088 11231
rect 10134 11228 10140 11280
rect 10192 11268 10198 11280
rect 10250 11271 10308 11277
rect 10250 11268 10262 11271
rect 10192 11240 10262 11268
rect 10192 11228 10198 11240
rect 10250 11237 10262 11240
rect 10296 11237 10308 11271
rect 10250 11231 10308 11237
rect 11885 11271 11943 11277
rect 11885 11237 11897 11271
rect 11931 11268 11943 11271
rect 12066 11268 12072 11280
rect 11931 11240 12072 11268
rect 11931 11237 11943 11240
rect 11885 11231 11943 11237
rect 12066 11228 12072 11240
rect 12124 11228 12130 11280
rect 12897 11271 12955 11277
rect 12897 11237 12909 11271
rect 12943 11268 12955 11271
rect 13078 11268 13084 11280
rect 12943 11240 13084 11268
rect 12943 11237 12955 11240
rect 12897 11231 12955 11237
rect 13078 11228 13084 11240
rect 13136 11228 13142 11280
rect 17862 11268 17868 11280
rect 17236 11240 17868 11268
rect 10410 11200 10416 11212
rect 10060 11172 10416 11200
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 11054 11160 11060 11212
rect 11112 11200 11118 11212
rect 12989 11203 13047 11209
rect 12989 11200 13001 11203
rect 11112 11172 13001 11200
rect 11112 11160 11118 11172
rect 12989 11169 13001 11172
rect 13035 11169 13047 11203
rect 15010 11200 15016 11212
rect 14971 11172 15016 11200
rect 12989 11163 13047 11169
rect 15010 11160 15016 11172
rect 15068 11160 15074 11212
rect 17236 11209 17264 11240
rect 17862 11228 17868 11240
rect 17920 11228 17926 11280
rect 18248 11268 18276 11308
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 21266 11268 21272 11280
rect 18248 11240 21272 11268
rect 21266 11228 21272 11240
rect 21324 11228 21330 11280
rect 17129 11203 17187 11209
rect 17129 11169 17141 11203
rect 17175 11200 17187 11203
rect 17221 11203 17279 11209
rect 17221 11200 17233 11203
rect 17175 11172 17233 11200
rect 17175 11169 17187 11172
rect 17129 11163 17187 11169
rect 17221 11169 17233 11172
rect 17267 11169 17279 11203
rect 17221 11163 17279 11169
rect 17678 11160 17684 11212
rect 17736 11200 17742 11212
rect 17773 11203 17831 11209
rect 17773 11200 17785 11203
rect 17736 11172 17785 11200
rect 17736 11160 17742 11172
rect 17773 11169 17785 11172
rect 17819 11169 17831 11203
rect 17773 11163 17831 11169
rect 19334 11160 19340 11212
rect 19392 11200 19398 11212
rect 20073 11203 20131 11209
rect 20073 11200 20085 11203
rect 19392 11172 20085 11200
rect 19392 11160 19398 11172
rect 20073 11169 20085 11172
rect 20119 11169 20131 11203
rect 20073 11163 20131 11169
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11101 8263 11135
rect 11790 11132 11796 11144
rect 11751 11104 11796 11132
rect 8205 11095 8263 11101
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 12066 11092 12072 11144
rect 12124 11132 12130 11144
rect 12713 11135 12771 11141
rect 12713 11132 12725 11135
rect 12124 11104 12725 11132
rect 12124 11092 12130 11104
rect 12713 11101 12725 11104
rect 12759 11132 12771 11135
rect 15286 11132 15292 11144
rect 12759 11104 15292 11132
rect 12759 11101 12771 11104
rect 12713 11095 12771 11101
rect 15286 11092 15292 11104
rect 15344 11132 15350 11144
rect 18046 11132 18052 11144
rect 15344 11104 18052 11132
rect 15344 11092 15350 11104
rect 18046 11092 18052 11104
rect 18104 11132 18110 11144
rect 18141 11135 18199 11141
rect 18141 11132 18153 11135
rect 18104 11104 18153 11132
rect 18104 11092 18110 11104
rect 18141 11101 18153 11104
rect 18187 11101 18199 11135
rect 18141 11095 18199 11101
rect 18325 11135 18383 11141
rect 18325 11101 18337 11135
rect 18371 11132 18383 11135
rect 21174 11132 21180 11144
rect 18371 11104 21180 11132
rect 18371 11101 18383 11104
rect 18325 11095 18383 11101
rect 21174 11092 21180 11104
rect 21232 11092 21238 11144
rect 7374 11064 7380 11076
rect 7335 11036 7380 11064
rect 7374 11024 7380 11036
rect 7432 11024 7438 11076
rect 7558 11024 7564 11076
rect 7616 11064 7622 11076
rect 7745 11067 7803 11073
rect 7745 11064 7757 11067
rect 7616 11036 7757 11064
rect 7616 11024 7622 11036
rect 7745 11033 7757 11036
rect 7791 11033 7803 11067
rect 11333 11067 11391 11073
rect 11333 11064 11345 11067
rect 7745 11027 7803 11033
rect 8220 11036 11345 11064
rect 8220 10996 8248 11036
rect 11333 11033 11345 11036
rect 11379 11033 11391 11067
rect 11333 11027 11391 11033
rect 13357 11067 13415 11073
rect 13357 11033 13369 11067
rect 13403 11064 13415 11067
rect 14826 11064 14832 11076
rect 13403 11036 14832 11064
rect 13403 11033 13415 11036
rect 13357 11027 13415 11033
rect 14826 11024 14832 11036
rect 14884 11024 14890 11076
rect 15197 11067 15255 11073
rect 15197 11033 15209 11067
rect 15243 11064 15255 11067
rect 15378 11064 15384 11076
rect 15243 11036 15384 11064
rect 15243 11033 15255 11036
rect 15197 11027 15255 11033
rect 15378 11024 15384 11036
rect 15436 11064 15442 11076
rect 17129 11067 17187 11073
rect 17129 11064 17141 11067
rect 15436 11036 17141 11064
rect 15436 11024 15442 11036
rect 17129 11033 17141 11036
rect 17175 11033 17187 11067
rect 18782 11064 18788 11076
rect 18743 11036 18788 11064
rect 17129 11027 17187 11033
rect 18782 11024 18788 11036
rect 18840 11024 18846 11076
rect 20162 11024 20168 11076
rect 20220 11064 20226 11076
rect 20257 11067 20315 11073
rect 20257 11064 20269 11067
rect 20220 11036 20269 11064
rect 20220 11024 20226 11036
rect 20257 11033 20269 11036
rect 20303 11033 20315 11067
rect 20257 11027 20315 11033
rect 7208 10968 8248 10996
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 10229 10999 10287 11005
rect 8352 10968 8397 10996
rect 8352 10956 8358 10968
rect 10229 10965 10241 10999
rect 10275 10996 10287 10999
rect 10962 10996 10968 11008
rect 10275 10968 10968 10996
rect 10275 10965 10287 10968
rect 10229 10959 10287 10965
rect 10962 10956 10968 10968
rect 11020 10956 11026 11008
rect 17218 10996 17224 11008
rect 17179 10968 17224 10996
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 1104 10906 21804 10928
rect 1104 10854 4432 10906
rect 4484 10854 4496 10906
rect 4548 10854 4560 10906
rect 4612 10854 4624 10906
rect 4676 10854 11332 10906
rect 11384 10854 11396 10906
rect 11448 10854 11460 10906
rect 11512 10854 11524 10906
rect 11576 10854 18232 10906
rect 18284 10854 18296 10906
rect 18348 10854 18360 10906
rect 18412 10854 18424 10906
rect 18476 10854 21804 10906
rect 1104 10832 21804 10854
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 4617 10795 4675 10801
rect 4617 10792 4629 10795
rect 4212 10764 4629 10792
rect 4212 10752 4218 10764
rect 4617 10761 4629 10764
rect 4663 10761 4675 10795
rect 4617 10755 4675 10761
rect 4985 10795 5043 10801
rect 4985 10761 4997 10795
rect 5031 10792 5043 10795
rect 5350 10792 5356 10804
rect 5031 10764 5356 10792
rect 5031 10761 5043 10764
rect 4985 10755 5043 10761
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 7929 10795 7987 10801
rect 7929 10761 7941 10795
rect 7975 10792 7987 10795
rect 11054 10792 11060 10804
rect 7975 10764 11060 10792
rect 7975 10761 7987 10764
rect 7929 10755 7987 10761
rect 6454 10684 6460 10736
rect 6512 10724 6518 10736
rect 6512 10696 6776 10724
rect 6512 10684 6518 10696
rect 6748 10668 6776 10696
rect 6730 10656 6736 10668
rect 6643 10628 6736 10656
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10656 6975 10659
rect 7944 10656 7972 10755
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 13449 10795 13507 10801
rect 13449 10761 13461 10795
rect 13495 10792 13507 10795
rect 13814 10792 13820 10804
rect 13495 10764 13820 10792
rect 13495 10761 13507 10764
rect 13449 10755 13507 10761
rect 13814 10752 13820 10764
rect 13872 10792 13878 10804
rect 15010 10792 15016 10804
rect 13872 10764 15016 10792
rect 13872 10752 13878 10764
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 15381 10795 15439 10801
rect 15381 10761 15393 10795
rect 15427 10792 15439 10795
rect 16117 10795 16175 10801
rect 16117 10792 16129 10795
rect 15427 10764 16129 10792
rect 15427 10761 15439 10764
rect 15381 10755 15439 10761
rect 6963 10628 7972 10656
rect 9309 10659 9367 10665
rect 6963 10625 6975 10628
rect 6917 10619 6975 10625
rect 9309 10625 9321 10659
rect 9355 10656 9367 10659
rect 10042 10656 10048 10668
rect 9355 10628 10048 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 12894 10616 12900 10668
rect 12952 10656 12958 10668
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 12952 10628 13093 10656
rect 12952 10616 12958 10628
rect 13081 10625 13093 10628
rect 13127 10625 13139 10659
rect 15749 10659 15807 10665
rect 15749 10656 15761 10659
rect 13081 10619 13139 10625
rect 14844 10628 15761 10656
rect 14844 10600 14872 10628
rect 15749 10625 15761 10628
rect 15795 10625 15807 10659
rect 15749 10619 15807 10625
rect 2682 10588 2688 10600
rect 2643 10560 2688 10588
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 4798 10588 4804 10600
rect 4759 10560 4804 10588
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 5077 10591 5135 10597
rect 5077 10557 5089 10591
rect 5123 10557 5135 10591
rect 6638 10588 6644 10600
rect 6599 10560 6644 10588
rect 5077 10551 5135 10557
rect 2866 10520 2872 10532
rect 2827 10492 2872 10520
rect 2866 10480 2872 10492
rect 2924 10480 2930 10532
rect 5092 10520 5120 10551
rect 6638 10548 6644 10560
rect 6696 10548 6702 10600
rect 6822 10588 6828 10600
rect 6783 10560 6828 10588
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10588 8079 10591
rect 8202 10588 8208 10600
rect 8067 10560 8208 10588
rect 8067 10557 8079 10560
rect 8021 10551 8079 10557
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 9122 10588 9128 10600
rect 9083 10560 9128 10588
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 9401 10591 9459 10597
rect 9401 10557 9413 10591
rect 9447 10557 9459 10591
rect 9401 10551 9459 10557
rect 5718 10520 5724 10532
rect 5092 10492 5724 10520
rect 5718 10480 5724 10492
rect 5776 10520 5782 10532
rect 6840 10520 6868 10548
rect 5776 10492 6868 10520
rect 9416 10520 9444 10551
rect 9490 10548 9496 10600
rect 9548 10588 9554 10600
rect 13449 10591 13507 10597
rect 9548 10560 9593 10588
rect 9548 10548 9554 10560
rect 13449 10557 13461 10591
rect 13495 10588 13507 10591
rect 13630 10588 13636 10600
rect 13495 10560 13636 10588
rect 13495 10557 13507 10560
rect 13449 10551 13507 10557
rect 13630 10548 13636 10560
rect 13688 10548 13694 10600
rect 14826 10588 14832 10600
rect 14787 10560 14832 10588
rect 14826 10548 14832 10560
rect 14884 10548 14890 10600
rect 15378 10588 15384 10600
rect 15339 10560 15384 10588
rect 15378 10548 15384 10560
rect 15436 10548 15442 10600
rect 9416 10492 9628 10520
rect 5776 10480 5782 10492
rect 9600 10464 9628 10492
rect 5442 10412 5448 10464
rect 5500 10452 5506 10464
rect 6457 10455 6515 10461
rect 6457 10452 6469 10455
rect 5500 10424 6469 10452
rect 5500 10412 5506 10424
rect 6457 10421 6469 10424
rect 6503 10421 6515 10455
rect 8938 10452 8944 10464
rect 8899 10424 8944 10452
rect 6457 10415 6515 10421
rect 8938 10412 8944 10424
rect 8996 10412 9002 10464
rect 9582 10452 9588 10464
rect 9543 10424 9588 10452
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 16040 10452 16068 10764
rect 16117 10761 16129 10764
rect 16163 10761 16175 10795
rect 17218 10792 17224 10804
rect 16117 10755 16175 10761
rect 17144 10764 17224 10792
rect 17144 10597 17172 10764
rect 17218 10752 17224 10764
rect 17276 10752 17282 10804
rect 17678 10792 17684 10804
rect 17639 10764 17684 10792
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 18509 10795 18567 10801
rect 18509 10792 18521 10795
rect 17788 10764 18521 10792
rect 17589 10659 17647 10665
rect 17589 10625 17601 10659
rect 17635 10656 17647 10659
rect 17696 10656 17724 10752
rect 17635 10628 17724 10656
rect 17635 10625 17647 10628
rect 17589 10619 17647 10625
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10588 16175 10591
rect 16945 10591 17003 10597
rect 16945 10588 16957 10591
rect 16163 10560 16957 10588
rect 16163 10557 16175 10560
rect 16117 10551 16175 10557
rect 16945 10557 16957 10560
rect 16991 10557 17003 10591
rect 16945 10551 17003 10557
rect 17129 10591 17187 10597
rect 17129 10557 17141 10591
rect 17175 10557 17187 10591
rect 17129 10551 17187 10557
rect 17221 10591 17279 10597
rect 17221 10557 17233 10591
rect 17267 10588 17279 10591
rect 17788 10588 17816 10764
rect 18509 10761 18521 10764
rect 18555 10761 18567 10795
rect 18509 10755 18567 10761
rect 19242 10752 19248 10804
rect 19300 10752 19306 10804
rect 19794 10752 19800 10804
rect 19852 10792 19858 10804
rect 20901 10795 20959 10801
rect 20901 10792 20913 10795
rect 19852 10764 20913 10792
rect 19852 10752 19858 10764
rect 20901 10761 20913 10764
rect 20947 10761 20959 10795
rect 20901 10755 20959 10761
rect 17862 10684 17868 10736
rect 17920 10724 17926 10736
rect 17920 10696 18736 10724
rect 17920 10684 17926 10696
rect 18046 10616 18052 10668
rect 18104 10656 18110 10668
rect 18233 10659 18291 10665
rect 18233 10656 18245 10659
rect 18104 10628 18245 10656
rect 18104 10616 18110 10628
rect 18233 10625 18245 10628
rect 18279 10625 18291 10659
rect 18233 10619 18291 10625
rect 18708 10597 18736 10696
rect 19150 10656 19156 10668
rect 19111 10628 19156 10656
rect 19150 10616 19156 10628
rect 19208 10616 19214 10668
rect 19260 10656 19288 10752
rect 19429 10659 19487 10665
rect 19429 10656 19441 10659
rect 19260 10628 19441 10656
rect 19429 10625 19441 10628
rect 19475 10625 19487 10659
rect 19429 10619 19487 10625
rect 17267 10560 17816 10588
rect 18693 10591 18751 10597
rect 17267 10557 17279 10560
rect 17221 10551 17279 10557
rect 18693 10557 18705 10591
rect 18739 10557 18751 10591
rect 18693 10551 18751 10557
rect 17954 10480 17960 10532
rect 18012 10520 18018 10532
rect 18049 10523 18107 10529
rect 18049 10520 18061 10523
rect 18012 10492 18061 10520
rect 18012 10480 18018 10492
rect 18049 10489 18061 10492
rect 18095 10489 18107 10523
rect 18049 10483 18107 10489
rect 20162 10480 20168 10532
rect 20220 10480 20226 10532
rect 16758 10452 16764 10464
rect 16040 10424 16764 10452
rect 16758 10412 16764 10424
rect 16816 10412 16822 10464
rect 18141 10455 18199 10461
rect 18141 10421 18153 10455
rect 18187 10452 18199 10455
rect 18874 10452 18880 10464
rect 18187 10424 18880 10452
rect 18187 10421 18199 10424
rect 18141 10415 18199 10421
rect 18874 10412 18880 10424
rect 18932 10412 18938 10464
rect 1104 10362 21804 10384
rect 1104 10310 7882 10362
rect 7934 10310 7946 10362
rect 7998 10310 8010 10362
rect 8062 10310 8074 10362
rect 8126 10310 14782 10362
rect 14834 10310 14846 10362
rect 14898 10310 14910 10362
rect 14962 10310 14974 10362
rect 15026 10310 21804 10362
rect 1104 10288 21804 10310
rect 1486 10248 1492 10260
rect 1447 10220 1492 10248
rect 1486 10208 1492 10220
rect 1544 10208 1550 10260
rect 5074 10208 5080 10260
rect 5132 10248 5138 10260
rect 5261 10251 5319 10257
rect 5261 10248 5273 10251
rect 5132 10220 5273 10248
rect 5132 10208 5138 10220
rect 5261 10217 5273 10220
rect 5307 10217 5319 10251
rect 6362 10248 6368 10260
rect 6323 10220 6368 10248
rect 5261 10211 5319 10217
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 9766 10208 9772 10260
rect 9824 10248 9830 10260
rect 12066 10248 12072 10260
rect 9824 10220 12072 10248
rect 9824 10208 9830 10220
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 13630 10248 13636 10260
rect 13591 10220 13636 10248
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 17218 10208 17224 10260
rect 17276 10248 17282 10260
rect 19150 10248 19156 10260
rect 17276 10220 19156 10248
rect 17276 10208 17282 10220
rect 19150 10208 19156 10220
rect 19208 10208 19214 10260
rect 21266 10248 21272 10260
rect 21227 10220 21272 10248
rect 21266 10208 21272 10220
rect 21324 10208 21330 10260
rect 5442 10180 5448 10192
rect 5403 10152 5448 10180
rect 5442 10140 5448 10152
rect 5500 10140 5506 10192
rect 6273 10183 6331 10189
rect 6273 10149 6285 10183
rect 6319 10180 6331 10183
rect 9122 10180 9128 10192
rect 6319 10152 9128 10180
rect 6319 10149 6331 10152
rect 6273 10143 6331 10149
rect 9122 10140 9128 10152
rect 9180 10180 9186 10192
rect 13357 10183 13415 10189
rect 9180 10152 10272 10180
rect 9180 10140 9186 10152
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10112 1639 10115
rect 1670 10112 1676 10124
rect 1627 10084 1676 10112
rect 1627 10081 1639 10084
rect 1581 10075 1639 10081
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 6822 10072 6828 10124
rect 6880 10112 6886 10124
rect 9766 10112 9772 10124
rect 6880 10084 9674 10112
rect 9727 10084 9772 10112
rect 6880 10072 6886 10084
rect 5166 10044 5172 10056
rect 5127 10016 5172 10044
rect 5166 10004 5172 10016
rect 5224 10044 5230 10056
rect 6457 10047 6515 10053
rect 6457 10044 6469 10047
rect 5224 10016 6469 10044
rect 5224 10004 5230 10016
rect 6457 10013 6469 10016
rect 6503 10013 6515 10047
rect 9214 10044 9220 10056
rect 9175 10016 9220 10044
rect 6457 10007 6515 10013
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9646 10044 9674 10084
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 10042 10112 10048 10124
rect 10003 10084 10048 10112
rect 10042 10072 10048 10084
rect 10100 10072 10106 10124
rect 10244 10121 10272 10152
rect 13357 10149 13369 10183
rect 13403 10180 13415 10183
rect 13814 10180 13820 10192
rect 13403 10152 13820 10180
rect 13403 10149 13415 10152
rect 13357 10143 13415 10149
rect 13814 10140 13820 10152
rect 13872 10140 13878 10192
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10081 10287 10115
rect 12894 10112 12900 10124
rect 12855 10084 12900 10112
rect 10229 10075 10287 10081
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 13446 10112 13452 10124
rect 13407 10084 13452 10112
rect 13446 10072 13452 10084
rect 13504 10072 13510 10124
rect 13538 10072 13544 10124
rect 13596 10112 13602 10124
rect 21450 10112 21456 10124
rect 13596 10084 13641 10112
rect 21411 10084 21456 10112
rect 13596 10072 13602 10084
rect 21450 10072 21456 10084
rect 21508 10072 21514 10124
rect 9953 10047 10011 10053
rect 9953 10044 9965 10047
rect 9646 10016 9965 10044
rect 9953 10013 9965 10016
rect 9999 10013 10011 10047
rect 9953 10007 10011 10013
rect 5721 9979 5779 9985
rect 5721 9945 5733 9979
rect 5767 9976 5779 9979
rect 10318 9976 10324 9988
rect 5767 9948 10324 9976
rect 5767 9945 5779 9948
rect 5721 9939 5779 9945
rect 10318 9936 10324 9948
rect 10376 9936 10382 9988
rect 5902 9908 5908 9920
rect 5863 9880 5908 9908
rect 5902 9868 5908 9880
rect 5960 9868 5966 9920
rect 10413 9911 10471 9917
rect 10413 9877 10425 9911
rect 10459 9908 10471 9911
rect 13354 9908 13360 9920
rect 10459 9880 13360 9908
rect 10459 9877 10471 9880
rect 10413 9871 10471 9877
rect 13354 9868 13360 9880
rect 13412 9868 13418 9920
rect 1104 9818 21804 9840
rect 1104 9766 4432 9818
rect 4484 9766 4496 9818
rect 4548 9766 4560 9818
rect 4612 9766 4624 9818
rect 4676 9766 11332 9818
rect 11384 9766 11396 9818
rect 11448 9766 11460 9818
rect 11512 9766 11524 9818
rect 11576 9766 18232 9818
rect 18284 9766 18296 9818
rect 18348 9766 18360 9818
rect 18412 9766 18424 9818
rect 18476 9766 21804 9818
rect 1104 9744 21804 9766
rect 2777 9639 2835 9645
rect 2777 9605 2789 9639
rect 2823 9636 2835 9639
rect 2869 9639 2927 9645
rect 2869 9636 2881 9639
rect 2823 9608 2881 9636
rect 2823 9605 2835 9608
rect 2777 9599 2835 9605
rect 2869 9605 2881 9608
rect 2915 9605 2927 9639
rect 2869 9599 2927 9605
rect 5261 9639 5319 9645
rect 5261 9605 5273 9639
rect 5307 9636 5319 9639
rect 12713 9639 12771 9645
rect 5307 9608 11744 9636
rect 5307 9605 5319 9608
rect 5261 9599 5319 9605
rect 2406 9568 2412 9580
rect 1780 9540 2412 9568
rect 1780 9509 1808 9540
rect 2406 9528 2412 9540
rect 2464 9528 2470 9580
rect 7282 9528 7288 9580
rect 7340 9568 7346 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 7340 9540 7389 9568
rect 7340 9528 7346 9540
rect 7377 9537 7389 9540
rect 7423 9537 7435 9571
rect 9214 9568 9220 9580
rect 7377 9531 7435 9537
rect 7944 9540 9220 9568
rect 1765 9503 1823 9509
rect 1765 9469 1777 9503
rect 1811 9469 1823 9503
rect 1765 9463 1823 9469
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9500 2375 9503
rect 2590 9500 2596 9512
rect 2363 9472 2596 9500
rect 2363 9469 2375 9472
rect 2317 9463 2375 9469
rect 2590 9460 2596 9472
rect 2648 9500 2654 9512
rect 2866 9500 2872 9512
rect 2648 9472 2872 9500
rect 2648 9460 2654 9472
rect 2866 9460 2872 9472
rect 2924 9500 2930 9512
rect 3053 9503 3111 9509
rect 3053 9500 3065 9503
rect 2924 9472 3065 9500
rect 2924 9460 2930 9472
rect 3053 9469 3065 9472
rect 3099 9469 3111 9503
rect 4982 9500 4988 9512
rect 4943 9472 4988 9500
rect 3053 9463 3111 9469
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 7944 9500 7972 9540
rect 8312 9509 8340 9540
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 9674 9568 9680 9580
rect 9635 9540 9680 9568
rect 9493 9531 9551 9537
rect 5184 9472 7972 9500
rect 8021 9503 8079 9509
rect 5184 9444 5212 9472
rect 8021 9469 8033 9503
rect 8067 9469 8079 9503
rect 8021 9463 8079 9469
rect 8297 9503 8355 9509
rect 8297 9469 8309 9503
rect 8343 9469 8355 9503
rect 8297 9463 8355 9469
rect 2222 9432 2228 9444
rect 2183 9404 2228 9432
rect 2222 9392 2228 9404
rect 2280 9392 2286 9444
rect 4614 9392 4620 9444
rect 4672 9432 4678 9444
rect 4709 9435 4767 9441
rect 4709 9432 4721 9435
rect 4672 9404 4721 9432
rect 4672 9392 4678 9404
rect 4709 9401 4721 9404
rect 4755 9432 4767 9435
rect 5166 9432 5172 9444
rect 4755 9404 5172 9432
rect 4755 9401 4767 9404
rect 4709 9395 4767 9401
rect 5166 9392 5172 9404
rect 5224 9392 5230 9444
rect 8036 9432 8064 9463
rect 8386 9432 8392 9444
rect 8036 9404 8392 9432
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 9508 9432 9536 9531
rect 9674 9528 9680 9540
rect 9732 9528 9738 9580
rect 10597 9571 10655 9577
rect 10597 9568 10609 9571
rect 9784 9540 10609 9568
rect 9582 9460 9588 9512
rect 9640 9500 9646 9512
rect 9784 9500 9812 9540
rect 10597 9537 10609 9540
rect 10643 9537 10655 9571
rect 10597 9531 10655 9537
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9568 10747 9571
rect 10962 9568 10968 9580
rect 10735 9540 10968 9568
rect 10735 9537 10747 9540
rect 10689 9531 10747 9537
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 11716 9568 11744 9608
rect 12713 9605 12725 9639
rect 12759 9636 12771 9639
rect 12805 9639 12863 9645
rect 12805 9636 12817 9639
rect 12759 9608 12817 9636
rect 12759 9605 12771 9608
rect 12713 9599 12771 9605
rect 12805 9605 12817 9608
rect 12851 9605 12863 9639
rect 12805 9599 12863 9605
rect 12345 9571 12403 9577
rect 12345 9568 12357 9571
rect 11716 9540 12357 9568
rect 10410 9500 10416 9512
rect 9640 9472 9812 9500
rect 10323 9472 10416 9500
rect 9640 9460 9646 9472
rect 10410 9460 10416 9472
rect 10468 9500 10474 9512
rect 11716 9509 11744 9540
rect 12345 9537 12357 9540
rect 12391 9537 12403 9571
rect 12345 9531 12403 9537
rect 11701 9503 11759 9509
rect 10468 9472 10548 9500
rect 10468 9460 10474 9472
rect 9674 9432 9680 9444
rect 9508 9404 9680 9432
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 9769 9435 9827 9441
rect 9769 9401 9781 9435
rect 9815 9432 9827 9435
rect 10229 9435 10287 9441
rect 10229 9432 10241 9435
rect 9815 9404 10241 9432
rect 9815 9401 9827 9404
rect 9769 9395 9827 9401
rect 10229 9401 10241 9404
rect 10275 9401 10287 9435
rect 10520 9432 10548 9472
rect 11701 9469 11713 9503
rect 11747 9469 11759 9503
rect 11701 9463 11759 9469
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 12434 9500 12440 9512
rect 12299 9472 12440 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 12434 9460 12440 9472
rect 12492 9500 12498 9512
rect 12989 9503 13047 9509
rect 12989 9500 13001 9503
rect 12492 9472 13001 9500
rect 12492 9460 12498 9472
rect 12989 9469 13001 9472
rect 13035 9500 13047 9503
rect 13446 9500 13452 9512
rect 13035 9472 13452 9500
rect 13035 9469 13047 9472
rect 12989 9463 13047 9469
rect 13446 9460 13452 9472
rect 13504 9460 13510 9512
rect 12066 9432 12072 9444
rect 10520 9404 12072 9432
rect 10229 9395 10287 9401
rect 12066 9392 12072 9404
rect 12124 9392 12130 9444
rect 12161 9435 12219 9441
rect 12161 9401 12173 9435
rect 12207 9432 12219 9435
rect 12207 9404 12434 9432
rect 12207 9401 12219 9404
rect 12161 9395 12219 9401
rect 2728 9364 2734 9376
rect 2689 9336 2734 9364
rect 2728 9324 2734 9336
rect 2786 9324 2792 9376
rect 4798 9364 4804 9376
rect 4759 9336 4804 9364
rect 4798 9324 4804 9336
rect 4856 9324 4862 9376
rect 10134 9364 10140 9376
rect 10095 9336 10140 9364
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 12406 9364 12434 9404
rect 12713 9367 12771 9373
rect 12713 9364 12725 9367
rect 12406 9336 12725 9364
rect 12713 9333 12725 9336
rect 12759 9364 12771 9367
rect 13538 9364 13544 9376
rect 12759 9336 13544 9364
rect 12759 9333 12771 9336
rect 12713 9327 12771 9333
rect 13538 9324 13544 9336
rect 13596 9324 13602 9376
rect 1104 9274 21804 9296
rect 1104 9222 7882 9274
rect 7934 9222 7946 9274
rect 7998 9222 8010 9274
rect 8062 9222 8074 9274
rect 8126 9222 14782 9274
rect 14834 9222 14846 9274
rect 14898 9222 14910 9274
rect 14962 9222 14974 9274
rect 15026 9222 21804 9274
rect 1104 9200 21804 9222
rect 2222 9120 2228 9172
rect 2280 9160 2286 9172
rect 2682 9160 2688 9172
rect 2280 9132 2688 9160
rect 2280 9120 2286 9132
rect 2682 9120 2688 9132
rect 2740 9120 2746 9172
rect 4893 9163 4951 9169
rect 4893 9129 4905 9163
rect 4939 9160 4951 9163
rect 6730 9160 6736 9172
rect 4939 9132 6736 9160
rect 4939 9129 4951 9132
rect 4893 9123 4951 9129
rect 6730 9120 6736 9132
rect 6788 9120 6794 9172
rect 10410 9160 10416 9172
rect 9508 9132 10416 9160
rect 1578 9052 1584 9104
rect 1636 9092 1642 9104
rect 1636 9064 6868 9092
rect 1636 9052 1642 9064
rect 4709 9027 4767 9033
rect 4709 8993 4721 9027
rect 4755 8993 4767 9027
rect 4709 8987 4767 8993
rect 4985 9027 5043 9033
rect 4985 8993 4997 9027
rect 5031 9024 5043 9027
rect 5350 9024 5356 9036
rect 5031 8996 5356 9024
rect 5031 8993 5043 8996
rect 4985 8987 5043 8993
rect 4614 8888 4620 8900
rect 2700 8860 4620 8888
rect 2700 8832 2728 8860
rect 4614 8848 4620 8860
rect 4672 8848 4678 8900
rect 4724 8888 4752 8987
rect 5350 8984 5356 8996
rect 5408 8984 5414 9036
rect 6641 9027 6699 9033
rect 6641 8993 6653 9027
rect 6687 9024 6699 9027
rect 6730 9024 6736 9036
rect 6687 8996 6736 9024
rect 6687 8993 6699 8996
rect 6641 8987 6699 8993
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 6840 9033 6868 9064
rect 9508 9033 9536 9132
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 14553 9163 14611 9169
rect 14553 9129 14565 9163
rect 14599 9160 14611 9163
rect 15197 9163 15255 9169
rect 15197 9160 15209 9163
rect 14599 9132 15209 9160
rect 14599 9129 14611 9132
rect 14553 9123 14611 9129
rect 15197 9129 15209 9132
rect 15243 9129 15255 9163
rect 15197 9123 15255 9129
rect 15289 9163 15347 9169
rect 15289 9129 15301 9163
rect 15335 9160 15347 9163
rect 15470 9160 15476 9172
rect 15335 9132 15476 9160
rect 15335 9129 15347 9132
rect 15289 9123 15347 9129
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 10962 9092 10968 9104
rect 9692 9064 10968 9092
rect 9692 9033 9720 9064
rect 10962 9052 10968 9064
rect 11020 9052 11026 9104
rect 11701 9095 11759 9101
rect 11701 9061 11713 9095
rect 11747 9092 11759 9095
rect 12434 9092 12440 9104
rect 11747 9064 12440 9092
rect 11747 9061 11759 9064
rect 11701 9055 11759 9061
rect 12434 9052 12440 9064
rect 12492 9052 12498 9104
rect 16758 9092 16764 9104
rect 16719 9064 16764 9092
rect 16758 9052 16764 9064
rect 16816 9052 16822 9104
rect 6825 9027 6883 9033
rect 6825 8993 6837 9027
rect 6871 8993 6883 9027
rect 6825 8987 6883 8993
rect 9493 9027 9551 9033
rect 9493 8993 9505 9027
rect 9539 8993 9551 9027
rect 9493 8987 9551 8993
rect 9677 9027 9735 9033
rect 9677 8993 9689 9027
rect 9723 8993 9735 9027
rect 9677 8987 9735 8993
rect 10410 8984 10416 9036
rect 10468 9024 10474 9036
rect 11517 9027 11575 9033
rect 11517 9024 11529 9027
rect 10468 8996 11529 9024
rect 10468 8984 10474 8996
rect 11517 8993 11529 8996
rect 11563 8993 11575 9027
rect 11517 8987 11575 8993
rect 12066 8984 12072 9036
rect 12124 9024 12130 9036
rect 14369 9027 14427 9033
rect 14369 9024 14381 9027
rect 12124 8996 14381 9024
rect 12124 8984 12130 8996
rect 14369 8993 14381 8996
rect 14415 8993 14427 9027
rect 14369 8987 14427 8993
rect 18417 9027 18475 9033
rect 18417 8993 18429 9027
rect 18463 9024 18475 9027
rect 18598 9024 18604 9036
rect 18463 8996 18604 9024
rect 18463 8993 18475 8996
rect 18417 8987 18475 8993
rect 18598 8984 18604 8996
rect 18656 8984 18662 9036
rect 7193 8959 7251 8965
rect 7193 8925 7205 8959
rect 7239 8956 7251 8959
rect 8386 8956 8392 8968
rect 7239 8928 8392 8956
rect 7239 8925 7251 8928
rect 7193 8919 7251 8925
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 15286 8916 15292 8968
rect 15344 8956 15350 8968
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 15344 8928 15393 8956
rect 15344 8916 15350 8928
rect 15381 8925 15393 8928
rect 15427 8925 15439 8959
rect 15381 8919 15439 8925
rect 8294 8888 8300 8900
rect 4724 8860 8300 8888
rect 8294 8848 8300 8860
rect 8352 8848 8358 8900
rect 1762 8780 1768 8832
rect 1820 8820 1826 8832
rect 2682 8820 2688 8832
rect 1820 8792 2688 8820
rect 1820 8780 1826 8792
rect 2682 8780 2688 8792
rect 2740 8780 2746 8832
rect 2777 8823 2835 8829
rect 2777 8789 2789 8823
rect 2823 8820 2835 8823
rect 3510 8820 3516 8832
rect 2823 8792 3516 8820
rect 2823 8789 2835 8792
rect 2777 8783 2835 8789
rect 3510 8780 3516 8792
rect 3568 8780 3574 8832
rect 3602 8780 3608 8832
rect 3660 8820 3666 8832
rect 4525 8823 4583 8829
rect 4525 8820 4537 8823
rect 3660 8792 4537 8820
rect 3660 8780 3666 8792
rect 4525 8789 4537 8792
rect 4571 8789 4583 8823
rect 9582 8820 9588 8832
rect 9543 8792 9588 8820
rect 4525 8783 4583 8789
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 9858 8820 9864 8832
rect 9819 8792 9864 8820
rect 9858 8780 9864 8792
rect 9916 8780 9922 8832
rect 14829 8823 14887 8829
rect 14829 8789 14841 8823
rect 14875 8820 14887 8823
rect 15102 8820 15108 8832
rect 14875 8792 15108 8820
rect 14875 8789 14887 8792
rect 14829 8783 14887 8789
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 16850 8820 16856 8832
rect 16811 8792 16856 8820
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 17310 8780 17316 8832
rect 17368 8820 17374 8832
rect 18325 8823 18383 8829
rect 18325 8820 18337 8823
rect 17368 8792 18337 8820
rect 17368 8780 17374 8792
rect 18325 8789 18337 8792
rect 18371 8789 18383 8823
rect 18325 8783 18383 8789
rect 1104 8730 21804 8752
rect 1104 8678 4432 8730
rect 4484 8678 4496 8730
rect 4548 8678 4560 8730
rect 4612 8678 4624 8730
rect 4676 8678 11332 8730
rect 11384 8678 11396 8730
rect 11448 8678 11460 8730
rect 11512 8678 11524 8730
rect 11576 8678 18232 8730
rect 18284 8678 18296 8730
rect 18348 8678 18360 8730
rect 18412 8678 18424 8730
rect 18476 8678 21804 8730
rect 1104 8656 21804 8678
rect 2130 8616 2136 8628
rect 2043 8588 2136 8616
rect 2130 8576 2136 8588
rect 2188 8616 2194 8628
rect 16758 8616 16764 8628
rect 2188 8588 2774 8616
rect 16671 8588 16764 8616
rect 2188 8576 2194 8588
rect 1581 8551 1639 8557
rect 1581 8517 1593 8551
rect 1627 8548 1639 8551
rect 2746 8548 2774 8588
rect 16758 8576 16764 8588
rect 16816 8616 16822 8628
rect 17313 8619 17371 8625
rect 17313 8616 17325 8619
rect 16816 8588 17325 8616
rect 16816 8576 16822 8588
rect 17313 8585 17325 8588
rect 17359 8585 17371 8619
rect 17313 8579 17371 8585
rect 7101 8551 7159 8557
rect 1627 8520 2636 8548
rect 2746 8520 3004 8548
rect 1627 8517 1639 8520
rect 1581 8511 1639 8517
rect 2608 8489 2636 8520
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8449 2651 8483
rect 2593 8443 2651 8449
rect 2682 8440 2688 8492
rect 2740 8480 2746 8492
rect 2976 8489 3004 8520
rect 7101 8517 7113 8551
rect 7147 8548 7159 8551
rect 19153 8551 19211 8557
rect 7147 8520 12434 8548
rect 7147 8517 7159 8520
rect 7101 8511 7159 8517
rect 2961 8483 3019 8489
rect 2740 8452 2785 8480
rect 2740 8440 2746 8452
rect 2961 8449 2973 8483
rect 3007 8449 3019 8483
rect 3510 8480 3516 8492
rect 3471 8452 3516 8480
rect 2961 8443 3019 8449
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 6638 8480 6644 8492
rect 6599 8452 6644 8480
rect 6638 8440 6644 8452
rect 6696 8440 6702 8492
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8480 8355 8483
rect 10410 8480 10416 8492
rect 8343 8452 10416 8480
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 12406 8480 12434 8520
rect 18156 8520 18920 8548
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 12406 8452 16957 8480
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8412 2559 8415
rect 3602 8412 3608 8424
rect 2547 8384 3608 8412
rect 2547 8381 2559 8384
rect 2501 8375 2559 8381
rect 3602 8372 3608 8384
rect 3660 8372 3666 8424
rect 5166 8372 5172 8424
rect 5224 8412 5230 8424
rect 6549 8415 6607 8421
rect 6549 8412 6561 8415
rect 5224 8384 6561 8412
rect 5224 8372 5230 8384
rect 6549 8381 6561 8384
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8412 7619 8415
rect 8386 8412 8392 8424
rect 7607 8384 8392 8412
rect 7607 8381 7619 8384
rect 7561 8375 7619 8381
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 8481 8415 8539 8421
rect 8481 8381 8493 8415
rect 8527 8412 8539 8415
rect 8573 8415 8631 8421
rect 8573 8412 8585 8415
rect 8527 8384 8585 8412
rect 8527 8381 8539 8384
rect 8481 8375 8539 8381
rect 8573 8381 8585 8384
rect 8619 8381 8631 8415
rect 8573 8375 8631 8381
rect 10962 8372 10968 8424
rect 11020 8412 11026 8424
rect 11885 8415 11943 8421
rect 11885 8412 11897 8415
rect 11020 8384 11897 8412
rect 11020 8372 11026 8384
rect 11885 8381 11897 8384
rect 11931 8381 11943 8415
rect 12066 8412 12072 8424
rect 12027 8384 12072 8412
rect 11885 8375 11943 8381
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 16224 8421 16252 8452
rect 16945 8449 16957 8452
rect 16991 8449 17003 8483
rect 17310 8480 17316 8492
rect 17271 8452 17316 8480
rect 16945 8443 17003 8449
rect 17310 8440 17316 8452
rect 17368 8440 17374 8492
rect 16209 8415 16267 8421
rect 16209 8381 16221 8415
rect 16255 8381 16267 8415
rect 16209 8375 16267 8381
rect 16761 8415 16819 8421
rect 16761 8381 16773 8415
rect 16807 8412 16819 8415
rect 16850 8412 16856 8424
rect 16807 8384 16856 8412
rect 16807 8381 16819 8384
rect 16761 8375 16819 8381
rect 16850 8372 16856 8384
rect 16908 8412 16914 8424
rect 18156 8421 18184 8520
rect 18782 8480 18788 8492
rect 18708 8452 18788 8480
rect 18708 8421 18736 8452
rect 18782 8440 18788 8452
rect 18840 8440 18846 8492
rect 18892 8480 18920 8520
rect 19153 8517 19165 8551
rect 19199 8548 19211 8551
rect 19245 8551 19303 8557
rect 19245 8548 19257 8551
rect 19199 8520 19257 8548
rect 19199 8517 19211 8520
rect 19153 8511 19211 8517
rect 19245 8517 19257 8520
rect 19291 8517 19303 8551
rect 19245 8511 19303 8517
rect 18892 8452 19472 8480
rect 19444 8421 19472 8452
rect 18141 8415 18199 8421
rect 18141 8412 18153 8415
rect 16908 8384 18153 8412
rect 16908 8372 16914 8384
rect 18141 8381 18153 8384
rect 18187 8381 18199 8415
rect 18141 8375 18199 8381
rect 18693 8415 18751 8421
rect 18693 8381 18705 8415
rect 18739 8381 18751 8415
rect 18693 8375 18751 8381
rect 19429 8415 19487 8421
rect 19429 8381 19441 8415
rect 19475 8381 19487 8415
rect 21450 8412 21456 8424
rect 21411 8384 21456 8412
rect 19429 8375 19487 8381
rect 21450 8372 21456 8384
rect 21508 8372 21514 8424
rect 3421 8347 3479 8353
rect 3421 8313 3433 8347
rect 3467 8344 3479 8347
rect 3970 8344 3976 8356
rect 3467 8316 3976 8344
rect 3467 8313 3479 8316
rect 3421 8307 3479 8313
rect 3970 8304 3976 8316
rect 4028 8304 4034 8356
rect 6638 8344 6644 8356
rect 6599 8316 6644 8344
rect 6638 8304 6644 8316
rect 6696 8304 6702 8356
rect 12253 8347 12311 8353
rect 12253 8313 12265 8347
rect 12299 8344 12311 8347
rect 12802 8344 12808 8356
rect 12299 8316 12808 8344
rect 12299 8313 12311 8316
rect 12253 8307 12311 8313
rect 12802 8304 12808 8316
rect 12860 8304 12866 8356
rect 18233 8347 18291 8353
rect 18233 8313 18245 8347
rect 18279 8344 18291 8347
rect 18598 8344 18604 8356
rect 18279 8316 18604 8344
rect 18279 8313 18291 8316
rect 18233 8307 18291 8313
rect 18598 8304 18604 8316
rect 18656 8344 18662 8356
rect 18656 8316 19196 8344
rect 18656 8304 18662 8316
rect 19168 8285 19196 8316
rect 19153 8279 19211 8285
rect 19153 8245 19165 8279
rect 19199 8245 19211 8279
rect 21266 8276 21272 8288
rect 21227 8248 21272 8276
rect 19153 8239 19211 8245
rect 21266 8236 21272 8248
rect 21324 8236 21330 8288
rect 1104 8186 21804 8208
rect 1104 8134 7882 8186
rect 7934 8134 7946 8186
rect 7998 8134 8010 8186
rect 8062 8134 8074 8186
rect 8126 8134 14782 8186
rect 14834 8134 14846 8186
rect 14898 8134 14910 8186
rect 14962 8134 14974 8186
rect 15026 8134 21804 8186
rect 1104 8112 21804 8134
rect 8570 8072 8576 8084
rect 8036 8044 8576 8072
rect 8036 8013 8064 8044
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 12802 8072 12808 8084
rect 12763 8044 12808 8072
rect 12802 8032 12808 8044
rect 12860 8032 12866 8084
rect 15381 8075 15439 8081
rect 15381 8041 15393 8075
rect 15427 8041 15439 8075
rect 15381 8035 15439 8041
rect 8021 8007 8079 8013
rect 8021 7973 8033 8007
rect 8067 7973 8079 8007
rect 8386 8004 8392 8016
rect 8347 7976 8392 8004
rect 8021 7967 8079 7973
rect 8386 7964 8392 7976
rect 8444 7964 8450 8016
rect 12897 8007 12955 8013
rect 12897 7973 12909 8007
rect 12943 8004 12955 8007
rect 15396 8004 15424 8035
rect 12943 7976 13584 8004
rect 12943 7973 12955 7976
rect 12897 7967 12955 7973
rect 2130 7936 2136 7948
rect 2091 7908 2136 7936
rect 2130 7896 2136 7908
rect 2188 7896 2194 7948
rect 2590 7896 2596 7948
rect 2648 7936 2654 7948
rect 2685 7939 2743 7945
rect 2685 7936 2697 7939
rect 2648 7908 2697 7936
rect 2648 7896 2654 7908
rect 2685 7905 2697 7908
rect 2731 7905 2743 7939
rect 7650 7936 7656 7948
rect 7611 7908 7656 7936
rect 2685 7899 2743 7905
rect 7650 7896 7656 7908
rect 7708 7896 7714 7948
rect 8570 7936 8576 7948
rect 8531 7908 8576 7936
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 9861 7939 9919 7945
rect 9861 7905 9873 7939
rect 9907 7936 9919 7939
rect 10226 7936 10232 7948
rect 9907 7908 10232 7936
rect 9907 7905 9919 7908
rect 9861 7899 9919 7905
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 9766 7828 9772 7880
rect 9824 7868 9830 7880
rect 12989 7871 13047 7877
rect 12989 7868 13001 7871
rect 9824 7840 13001 7868
rect 9824 7828 9830 7840
rect 12989 7837 13001 7840
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 2685 7735 2743 7741
rect 2685 7701 2697 7735
rect 2731 7732 2743 7735
rect 3970 7732 3976 7744
rect 2731 7704 3976 7732
rect 2731 7701 2743 7704
rect 2685 7695 2743 7701
rect 3970 7692 3976 7704
rect 4028 7692 4034 7744
rect 8297 7735 8355 7741
rect 8297 7701 8309 7735
rect 8343 7732 8355 7735
rect 9398 7732 9404 7744
rect 8343 7704 9404 7732
rect 8343 7701 8355 7704
rect 8297 7695 8355 7701
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 9490 7692 9496 7744
rect 9548 7732 9554 7744
rect 9769 7735 9827 7741
rect 9769 7732 9781 7735
rect 9548 7704 9781 7732
rect 9548 7692 9554 7704
rect 9769 7701 9781 7704
rect 9815 7701 9827 7735
rect 9769 7695 9827 7701
rect 12342 7692 12348 7744
rect 12400 7732 12406 7744
rect 12437 7735 12495 7741
rect 12437 7732 12449 7735
rect 12400 7704 12449 7732
rect 12400 7692 12406 7704
rect 12437 7701 12449 7704
rect 12483 7701 12495 7735
rect 13556 7732 13584 7976
rect 14660 7976 15424 8004
rect 16393 8007 16451 8013
rect 14366 7936 14372 7948
rect 14327 7908 14372 7936
rect 14366 7896 14372 7908
rect 14424 7896 14430 7948
rect 14458 7896 14464 7948
rect 14516 7936 14522 7948
rect 14660 7936 14688 7976
rect 16393 7973 16405 8007
rect 16439 8004 16451 8007
rect 16758 8004 16764 8016
rect 16439 7976 16764 8004
rect 16439 7973 16451 7976
rect 16393 7967 16451 7973
rect 16758 7964 16764 7976
rect 16816 7964 16822 8016
rect 14516 7908 14688 7936
rect 14921 7939 14979 7945
rect 14516 7896 14522 7908
rect 14921 7905 14933 7939
rect 14967 7936 14979 7939
rect 15013 7939 15071 7945
rect 15013 7936 15025 7939
rect 14967 7908 15025 7936
rect 14967 7905 14979 7908
rect 14921 7899 14979 7905
rect 15013 7905 15025 7908
rect 15059 7905 15071 7939
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 15013 7899 15071 7905
rect 15120 7908 15669 7936
rect 13722 7828 13728 7880
rect 13780 7868 13786 7880
rect 14936 7868 14964 7899
rect 13780 7840 14964 7868
rect 13780 7828 13786 7840
rect 14366 7760 14372 7812
rect 14424 7800 14430 7812
rect 15120 7800 15148 7908
rect 15657 7905 15669 7908
rect 15703 7936 15715 7939
rect 16209 7939 16267 7945
rect 16209 7936 16221 7939
rect 15703 7908 16221 7936
rect 15703 7905 15715 7908
rect 15657 7899 15715 7905
rect 16209 7905 16221 7908
rect 16255 7905 16267 7939
rect 16209 7899 16267 7905
rect 21266 7868 21272 7880
rect 16546 7840 21272 7868
rect 14424 7772 15148 7800
rect 15381 7803 15439 7809
rect 14424 7760 14430 7772
rect 15381 7769 15393 7803
rect 15427 7800 15439 7803
rect 15473 7803 15531 7809
rect 15473 7800 15485 7803
rect 15427 7772 15485 7800
rect 15427 7769 15439 7772
rect 15381 7763 15439 7769
rect 15473 7769 15485 7772
rect 15519 7769 15531 7803
rect 15473 7763 15531 7769
rect 16546 7732 16574 7840
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 13556 7704 16574 7732
rect 12437 7695 12495 7701
rect 1104 7642 21804 7664
rect 1104 7590 4432 7642
rect 4484 7590 4496 7642
rect 4548 7590 4560 7642
rect 4612 7590 4624 7642
rect 4676 7590 11332 7642
rect 11384 7590 11396 7642
rect 11448 7590 11460 7642
rect 11512 7590 11524 7642
rect 11576 7590 18232 7642
rect 18284 7590 18296 7642
rect 18348 7590 18360 7642
rect 18412 7590 18424 7642
rect 18476 7590 21804 7642
rect 1104 7568 21804 7590
rect 7650 7528 7656 7540
rect 7611 7500 7656 7528
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 12710 7488 12716 7540
rect 12768 7528 12774 7540
rect 12805 7531 12863 7537
rect 12805 7528 12817 7531
rect 12768 7500 12817 7528
rect 12768 7488 12774 7500
rect 12805 7497 12817 7500
rect 12851 7528 12863 7531
rect 13265 7531 13323 7537
rect 13265 7528 13277 7531
rect 12851 7500 13277 7528
rect 12851 7497 12863 7500
rect 12805 7491 12863 7497
rect 13265 7497 13277 7500
rect 13311 7497 13323 7531
rect 13265 7491 13323 7497
rect 2958 7420 2964 7472
rect 3016 7460 3022 7472
rect 3697 7463 3755 7469
rect 3697 7460 3709 7463
rect 3016 7432 3709 7460
rect 3016 7420 3022 7432
rect 3697 7429 3709 7432
rect 3743 7429 3755 7463
rect 3697 7423 3755 7429
rect 8570 7392 8576 7404
rect 8531 7364 8576 7392
rect 8570 7352 8576 7364
rect 8628 7352 8634 7404
rect 9398 7352 9404 7404
rect 9456 7392 9462 7404
rect 9456 7364 9720 7392
rect 9456 7352 9462 7364
rect 7837 7327 7895 7333
rect 7837 7293 7849 7327
rect 7883 7293 7895 7327
rect 9490 7324 9496 7336
rect 9451 7296 9496 7324
rect 7837 7287 7895 7293
rect 3878 7256 3884 7268
rect 3839 7228 3884 7256
rect 3878 7216 3884 7228
rect 3936 7216 3942 7268
rect 7852 7256 7880 7287
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 9692 7333 9720 7364
rect 12342 7352 12348 7404
rect 12400 7392 12406 7404
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 12400 7364 12909 7392
rect 12400 7352 12434 7364
rect 12897 7361 12909 7364
rect 12943 7361 12955 7395
rect 14366 7392 14372 7404
rect 12897 7355 12955 7361
rect 13188 7364 14372 7392
rect 9677 7327 9735 7333
rect 9677 7293 9689 7327
rect 9723 7293 9735 7327
rect 10410 7324 10416 7336
rect 10371 7296 10416 7324
rect 9677 7287 9735 7293
rect 10410 7284 10416 7296
rect 10468 7284 10474 7336
rect 12253 7327 12311 7333
rect 12253 7293 12265 7327
rect 12299 7324 12311 7327
rect 12406 7324 12434 7352
rect 12299 7296 12434 7324
rect 12805 7327 12863 7333
rect 12299 7293 12311 7296
rect 12253 7287 12311 7293
rect 12805 7293 12817 7327
rect 12851 7324 12863 7327
rect 13188 7324 13216 7364
rect 14366 7352 14372 7364
rect 14424 7352 14430 7404
rect 12851 7296 13216 7324
rect 13265 7327 13323 7333
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 13265 7293 13277 7327
rect 13311 7324 13323 7327
rect 14093 7327 14151 7333
rect 14093 7324 14105 7327
rect 13311 7296 14105 7324
rect 13311 7293 13323 7296
rect 13265 7287 13323 7293
rect 14093 7293 14105 7296
rect 14139 7293 14151 7327
rect 14093 7287 14151 7293
rect 14277 7327 14335 7333
rect 14277 7293 14289 7327
rect 14323 7324 14335 7327
rect 14458 7324 14464 7336
rect 14323 7296 14464 7324
rect 14323 7293 14335 7296
rect 14277 7287 14335 7293
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 9217 7259 9275 7265
rect 9217 7256 9229 7259
rect 7852 7228 9229 7256
rect 9217 7225 9229 7228
rect 9263 7256 9275 7259
rect 10428 7256 10456 7284
rect 10594 7256 10600 7268
rect 9263 7228 10456 7256
rect 10555 7228 10600 7256
rect 9263 7225 9275 7228
rect 9217 7219 9275 7225
rect 10594 7216 10600 7228
rect 10652 7216 10658 7268
rect 1104 7098 21804 7120
rect 1104 7046 7882 7098
rect 7934 7046 7946 7098
rect 7998 7046 8010 7098
rect 8062 7046 8074 7098
rect 8126 7046 14782 7098
rect 14834 7046 14846 7098
rect 14898 7046 14910 7098
rect 14962 7046 14974 7098
rect 15026 7046 21804 7098
rect 1104 7024 21804 7046
rect 8294 6984 8300 6996
rect 8255 6956 8300 6984
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 8570 6944 8576 6996
rect 8628 6984 8634 6996
rect 8665 6987 8723 6993
rect 8665 6984 8677 6987
rect 8628 6956 8677 6984
rect 8628 6944 8634 6956
rect 8665 6953 8677 6956
rect 8711 6953 8723 6987
rect 10873 6987 10931 6993
rect 10873 6984 10885 6987
rect 8665 6947 8723 6953
rect 10336 6956 10885 6984
rect 4816 6888 5028 6916
rect 4249 6851 4307 6857
rect 4249 6817 4261 6851
rect 4295 6848 4307 6851
rect 4816 6848 4844 6888
rect 4295 6820 4844 6848
rect 4893 6851 4951 6857
rect 4295 6817 4307 6820
rect 4249 6811 4307 6817
rect 4893 6817 4905 6851
rect 4939 6817 4951 6851
rect 4893 6811 4951 6817
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 4908 6780 4936 6811
rect 3936 6752 4936 6780
rect 5000 6780 5028 6888
rect 10226 6876 10232 6928
rect 10284 6916 10290 6928
rect 10336 6925 10364 6956
rect 10873 6953 10885 6956
rect 10919 6953 10931 6987
rect 10873 6947 10931 6953
rect 10321 6919 10379 6925
rect 10321 6916 10333 6919
rect 10284 6888 10333 6916
rect 10284 6876 10290 6888
rect 10321 6885 10333 6888
rect 10367 6885 10379 6919
rect 10321 6879 10379 6885
rect 5169 6851 5227 6857
rect 5169 6817 5181 6851
rect 5215 6848 5227 6851
rect 5534 6848 5540 6860
rect 5215 6820 5540 6848
rect 5215 6817 5227 6820
rect 5169 6811 5227 6817
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 5813 6851 5871 6857
rect 5813 6817 5825 6851
rect 5859 6848 5871 6851
rect 5905 6851 5963 6857
rect 5905 6848 5917 6851
rect 5859 6820 5917 6848
rect 5859 6817 5871 6820
rect 5813 6811 5871 6817
rect 5905 6817 5917 6820
rect 5951 6817 5963 6851
rect 5905 6811 5963 6817
rect 6089 6851 6147 6857
rect 6089 6817 6101 6851
rect 6135 6848 6147 6851
rect 6178 6848 6184 6860
rect 6135 6820 6184 6848
rect 6135 6817 6147 6820
rect 6089 6811 6147 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 8478 6848 8484 6860
rect 8128 6820 8484 6848
rect 5258 6780 5264 6792
rect 5000 6752 5264 6780
rect 3936 6740 3942 6752
rect 4908 6712 4936 6752
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 8128 6789 8156 6820
rect 8478 6808 8484 6820
rect 8536 6848 8542 6860
rect 9766 6848 9772 6860
rect 8536 6820 9772 6848
rect 8536 6808 8542 6820
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 9861 6851 9919 6857
rect 9861 6817 9873 6851
rect 9907 6848 9919 6851
rect 10134 6848 10140 6860
rect 9907 6820 10140 6848
rect 9907 6817 9919 6820
rect 9861 6811 9919 6817
rect 10134 6808 10140 6820
rect 10192 6848 10198 6860
rect 10425 6851 10483 6857
rect 10192 6820 10364 6848
rect 10192 6808 10198 6820
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6780 8263 6783
rect 10336 6780 10364 6820
rect 10425 6817 10437 6851
rect 10471 6848 10483 6851
rect 10594 6848 10600 6860
rect 10471 6820 10600 6848
rect 10471 6817 10483 6820
rect 10425 6811 10483 6817
rect 10594 6808 10600 6820
rect 10652 6848 10658 6860
rect 11146 6848 11152 6860
rect 10652 6820 11152 6848
rect 10652 6808 10658 6820
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 15930 6848 15936 6860
rect 15891 6820 15936 6848
rect 15930 6808 15936 6820
rect 15988 6808 15994 6860
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6848 16083 6851
rect 17218 6848 17224 6860
rect 16071 6820 17224 6848
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 10505 6783 10563 6789
rect 10505 6780 10517 6783
rect 8251 6752 10272 6780
rect 10336 6752 10517 6780
rect 8251 6749 8263 6752
rect 8205 6743 8263 6749
rect 5721 6715 5779 6721
rect 5721 6712 5733 6715
rect 4908 6684 5733 6712
rect 5721 6681 5733 6684
rect 5767 6681 5779 6715
rect 10244 6712 10272 6752
rect 10505 6749 10517 6752
rect 10551 6749 10563 6783
rect 16206 6780 16212 6792
rect 10505 6743 10563 6749
rect 10796 6752 12434 6780
rect 16167 6752 16212 6780
rect 10796 6712 10824 6752
rect 10244 6684 10824 6712
rect 10873 6715 10931 6721
rect 5721 6675 5779 6681
rect 10873 6681 10885 6715
rect 10919 6712 10931 6715
rect 10965 6715 11023 6721
rect 10965 6712 10977 6715
rect 10919 6684 10977 6712
rect 10919 6681 10931 6684
rect 10873 6675 10931 6681
rect 10965 6681 10977 6684
rect 11011 6681 11023 6715
rect 12406 6712 12434 6752
rect 16206 6740 16212 6752
rect 16264 6740 16270 6792
rect 21913 6715 21971 6721
rect 21913 6712 21925 6715
rect 12406 6684 21925 6712
rect 10965 6675 11023 6681
rect 21913 6681 21925 6684
rect 21959 6681 21971 6715
rect 21913 6675 21971 6681
rect 1670 6604 1676 6656
rect 1728 6644 1734 6656
rect 15565 6647 15623 6653
rect 15565 6644 15577 6647
rect 1728 6616 15577 6644
rect 1728 6604 1734 6616
rect 15565 6613 15577 6616
rect 15611 6613 15623 6647
rect 15565 6607 15623 6613
rect 1104 6554 21804 6576
rect 1104 6502 4432 6554
rect 4484 6502 4496 6554
rect 4548 6502 4560 6554
rect 4612 6502 4624 6554
rect 4676 6502 11332 6554
rect 11384 6502 11396 6554
rect 11448 6502 11460 6554
rect 11512 6502 11524 6554
rect 11576 6502 18232 6554
rect 18284 6502 18296 6554
rect 18348 6502 18360 6554
rect 18412 6502 18424 6554
rect 18476 6502 21804 6554
rect 1104 6480 21804 6502
rect 6825 6375 6883 6381
rect 6825 6341 6837 6375
rect 6871 6372 6883 6375
rect 6917 6375 6975 6381
rect 6917 6372 6929 6375
rect 6871 6344 6929 6372
rect 6871 6341 6883 6344
rect 6825 6335 6883 6341
rect 6917 6341 6929 6344
rect 6963 6341 6975 6375
rect 6917 6335 6975 6341
rect 5552 6276 7144 6304
rect 5552 6248 5580 6276
rect 3478 6239 3536 6245
rect 3478 6205 3490 6239
rect 3524 6236 3536 6239
rect 3878 6236 3884 6248
rect 3524 6208 3884 6236
rect 3524 6205 3536 6208
rect 3478 6199 3536 6205
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 5534 6236 5540 6248
rect 5495 6208 5540 6236
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 5902 6196 5908 6248
rect 5960 6236 5966 6248
rect 6089 6239 6147 6245
rect 6089 6236 6101 6239
rect 5960 6208 6101 6236
rect 5960 6196 5966 6208
rect 6089 6205 6101 6208
rect 6135 6236 6147 6239
rect 6457 6239 6515 6245
rect 6457 6236 6469 6239
rect 6135 6208 6469 6236
rect 6135 6205 6147 6208
rect 6089 6199 6147 6205
rect 6457 6205 6469 6208
rect 6503 6205 6515 6239
rect 6457 6199 6515 6205
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7116 6245 7144 6276
rect 16206 6264 16212 6316
rect 16264 6304 16270 6316
rect 17221 6307 17279 6313
rect 17221 6304 17233 6307
rect 16264 6276 17233 6304
rect 16264 6264 16270 6276
rect 17221 6273 17233 6276
rect 17267 6273 17279 6307
rect 17221 6267 17279 6273
rect 17405 6307 17463 6313
rect 17405 6273 17417 6307
rect 17451 6304 17463 6307
rect 18230 6304 18236 6316
rect 17451 6276 18236 6304
rect 17451 6273 17463 6276
rect 17405 6267 17463 6273
rect 18230 6264 18236 6276
rect 18288 6264 18294 6316
rect 7101 6239 7159 6245
rect 7101 6236 7113 6239
rect 6972 6208 7113 6236
rect 6972 6196 6978 6208
rect 7101 6205 7113 6208
rect 7147 6205 7159 6239
rect 17586 6236 17592 6248
rect 17547 6208 17592 6236
rect 7101 6199 7159 6205
rect 17586 6196 17592 6208
rect 17644 6196 17650 6248
rect 17773 6239 17831 6245
rect 17773 6205 17785 6239
rect 17819 6205 17831 6239
rect 17773 6199 17831 6205
rect 5629 6171 5687 6177
rect 5629 6137 5641 6171
rect 5675 6168 5687 6171
rect 6178 6168 6184 6180
rect 5675 6140 6184 6168
rect 5675 6137 5687 6140
rect 5629 6131 5687 6137
rect 6178 6128 6184 6140
rect 6236 6168 6242 6180
rect 17788 6168 17816 6199
rect 18046 6196 18052 6248
rect 18104 6236 18110 6248
rect 18141 6239 18199 6245
rect 18141 6236 18153 6239
rect 18104 6208 18153 6236
rect 18104 6196 18110 6208
rect 18141 6205 18153 6208
rect 18187 6205 18199 6239
rect 18141 6199 18199 6205
rect 18325 6239 18383 6245
rect 18325 6205 18337 6239
rect 18371 6236 18383 6239
rect 18414 6236 18420 6248
rect 18371 6208 18420 6236
rect 18371 6205 18383 6208
rect 18325 6199 18383 6205
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 18509 6239 18567 6245
rect 18509 6205 18521 6239
rect 18555 6205 18567 6239
rect 18509 6199 18567 6205
rect 18524 6168 18552 6199
rect 18690 6168 18696 6180
rect 6236 6140 6868 6168
rect 6236 6128 6242 6140
rect 2774 6060 2780 6112
rect 2832 6100 2838 6112
rect 6840 6109 6868 6140
rect 17420 6140 18696 6168
rect 17420 6112 17448 6140
rect 18690 6128 18696 6140
rect 18748 6128 18754 6180
rect 3375 6103 3433 6109
rect 3375 6100 3387 6103
rect 2832 6072 3387 6100
rect 2832 6060 2838 6072
rect 3375 6069 3387 6072
rect 3421 6069 3433 6103
rect 3375 6063 3433 6069
rect 6825 6103 6883 6109
rect 6825 6069 6837 6103
rect 6871 6069 6883 6103
rect 6825 6063 6883 6069
rect 17402 6060 17408 6112
rect 17460 6060 17466 6112
rect 18509 6103 18567 6109
rect 18509 6069 18521 6103
rect 18555 6100 18567 6103
rect 18598 6100 18604 6112
rect 18555 6072 18604 6100
rect 18555 6069 18567 6072
rect 18509 6063 18567 6069
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 1104 6010 21804 6032
rect 1104 5958 7882 6010
rect 7934 5958 7946 6010
rect 7998 5958 8010 6010
rect 8062 5958 8074 6010
rect 8126 5958 14782 6010
rect 14834 5958 14846 6010
rect 14898 5958 14910 6010
rect 14962 5958 14974 6010
rect 15026 5958 21804 6010
rect 1104 5936 21804 5958
rect 6914 5896 6920 5908
rect 6875 5868 6920 5896
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 15930 5856 15936 5908
rect 15988 5896 15994 5908
rect 16117 5899 16175 5905
rect 16117 5896 16129 5899
rect 15988 5868 16129 5896
rect 15988 5856 15994 5868
rect 16117 5865 16129 5868
rect 16163 5865 16175 5899
rect 16117 5859 16175 5865
rect 17497 5899 17555 5905
rect 17497 5865 17509 5899
rect 17543 5865 17555 5899
rect 17497 5859 17555 5865
rect 21269 5899 21327 5905
rect 21269 5865 21281 5899
rect 21315 5896 21327 5899
rect 21913 5899 21971 5905
rect 21913 5896 21925 5899
rect 21315 5868 21925 5896
rect 21315 5865 21327 5868
rect 21269 5859 21327 5865
rect 21913 5865 21925 5868
rect 21959 5865 21971 5899
rect 21913 5859 21971 5865
rect 1581 5831 1639 5837
rect 1581 5797 1593 5831
rect 1627 5828 1639 5831
rect 4982 5828 4988 5840
rect 1627 5800 4988 5828
rect 1627 5797 1639 5800
rect 1581 5791 1639 5797
rect 4982 5788 4988 5800
rect 5040 5788 5046 5840
rect 12710 5828 12716 5840
rect 12671 5800 12716 5828
rect 12710 5788 12716 5800
rect 12768 5788 12774 5840
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 7006 5760 7012 5772
rect 2832 5732 2877 5760
rect 6967 5732 7012 5760
rect 2832 5720 2838 5732
rect 7006 5720 7012 5732
rect 7064 5720 7070 5772
rect 14553 5763 14611 5769
rect 14553 5729 14565 5763
rect 14599 5760 14611 5763
rect 14826 5760 14832 5772
rect 14599 5732 14832 5760
rect 14599 5729 14611 5732
rect 14553 5723 14611 5729
rect 14826 5720 14832 5732
rect 14884 5720 14890 5772
rect 15102 5760 15108 5772
rect 15063 5732 15108 5760
rect 15102 5720 15108 5732
rect 15160 5760 15166 5772
rect 15565 5763 15623 5769
rect 15565 5760 15577 5763
rect 15160 5732 15577 5760
rect 15160 5720 15166 5732
rect 15565 5729 15577 5732
rect 15611 5729 15623 5763
rect 15565 5723 15623 5729
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5760 16543 5763
rect 16942 5760 16948 5772
rect 16531 5732 16948 5760
rect 16531 5729 16543 5732
rect 16485 5723 16543 5729
rect 16942 5720 16948 5732
rect 17000 5720 17006 5772
rect 17402 5760 17408 5772
rect 17363 5732 17408 5760
rect 17402 5720 17408 5732
rect 17460 5720 17466 5772
rect 15194 5692 15200 5704
rect 15155 5664 15200 5692
rect 15194 5652 15200 5664
rect 15252 5652 15258 5704
rect 15286 5652 15292 5704
rect 15344 5692 15350 5704
rect 16577 5695 16635 5701
rect 16577 5692 16589 5695
rect 15344 5664 16589 5692
rect 15344 5652 15350 5664
rect 16577 5661 16589 5664
rect 16623 5661 16635 5695
rect 16577 5655 16635 5661
rect 16761 5695 16819 5701
rect 16761 5661 16773 5695
rect 16807 5692 16819 5695
rect 17512 5692 17540 5859
rect 17586 5788 17592 5840
rect 17644 5828 17650 5840
rect 17644 5800 19104 5828
rect 17644 5788 17650 5800
rect 17788 5769 17816 5800
rect 17773 5763 17831 5769
rect 17773 5729 17785 5763
rect 17819 5729 17831 5763
rect 17773 5723 17831 5729
rect 17865 5763 17923 5769
rect 17865 5729 17877 5763
rect 17911 5760 17923 5763
rect 18046 5760 18052 5772
rect 17911 5732 18052 5760
rect 17911 5729 17923 5732
rect 17865 5723 17923 5729
rect 18046 5720 18052 5732
rect 18104 5720 18110 5772
rect 18414 5720 18420 5772
rect 18472 5760 18478 5772
rect 18509 5763 18567 5769
rect 18509 5760 18521 5763
rect 18472 5732 18521 5760
rect 18472 5720 18478 5732
rect 18509 5729 18521 5732
rect 18555 5729 18567 5763
rect 18690 5760 18696 5772
rect 18651 5732 18696 5760
rect 18509 5723 18567 5729
rect 16807 5664 17540 5692
rect 16807 5661 16819 5664
rect 16761 5655 16819 5661
rect 17954 5652 17960 5704
rect 18012 5692 18018 5704
rect 18141 5695 18199 5701
rect 18141 5692 18153 5695
rect 18012 5664 18153 5692
rect 18012 5652 18018 5664
rect 18141 5661 18153 5664
rect 18187 5661 18199 5695
rect 18141 5655 18199 5661
rect 18230 5652 18236 5704
rect 18288 5692 18294 5704
rect 18325 5695 18383 5701
rect 18325 5692 18337 5695
rect 18288 5664 18337 5692
rect 18288 5652 18294 5664
rect 18325 5661 18337 5664
rect 18371 5661 18383 5695
rect 18524 5692 18552 5723
rect 18690 5720 18696 5732
rect 18748 5720 18754 5772
rect 19076 5769 19104 5800
rect 19061 5763 19119 5769
rect 19061 5729 19073 5763
rect 19107 5760 19119 5763
rect 20806 5760 20812 5772
rect 19107 5732 20812 5760
rect 19107 5729 19119 5732
rect 19061 5723 19119 5729
rect 20806 5720 20812 5732
rect 20864 5720 20870 5772
rect 21450 5760 21456 5772
rect 21411 5732 21456 5760
rect 21450 5720 21456 5732
rect 21508 5720 21514 5772
rect 18969 5695 19027 5701
rect 18969 5692 18981 5695
rect 18524 5664 18981 5692
rect 18325 5655 18383 5661
rect 18969 5661 18981 5664
rect 19015 5661 19027 5695
rect 18969 5655 19027 5661
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 12529 5627 12587 5633
rect 12529 5624 12541 5627
rect 9732 5596 12541 5624
rect 9732 5584 9738 5596
rect 12529 5593 12541 5596
rect 12575 5593 12587 5627
rect 18340 5624 18368 5655
rect 18690 5624 18696 5636
rect 18340 5596 18696 5624
rect 12529 5587 12587 5593
rect 18690 5584 18696 5596
rect 18748 5584 18754 5636
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 2682 5556 2688 5568
rect 2643 5528 2688 5556
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 14553 5559 14611 5565
rect 14553 5525 14565 5559
rect 14599 5556 14611 5559
rect 14734 5556 14740 5568
rect 14599 5528 14740 5556
rect 14599 5525 14611 5528
rect 14553 5519 14611 5525
rect 14734 5516 14740 5528
rect 14792 5556 14798 5568
rect 15197 5559 15255 5565
rect 15197 5556 15209 5559
rect 14792 5528 15209 5556
rect 14792 5516 14798 5528
rect 15197 5525 15209 5528
rect 15243 5525 15255 5559
rect 15197 5519 15255 5525
rect 1104 5466 21804 5488
rect 1104 5414 4432 5466
rect 4484 5414 4496 5466
rect 4548 5414 4560 5466
rect 4612 5414 4624 5466
rect 4676 5414 11332 5466
rect 11384 5414 11396 5466
rect 11448 5414 11460 5466
rect 11512 5414 11524 5466
rect 11576 5414 18232 5466
rect 18284 5414 18296 5466
rect 18348 5414 18360 5466
rect 18412 5414 18424 5466
rect 18476 5414 21804 5466
rect 1104 5392 21804 5414
rect 7006 5312 7012 5364
rect 7064 5352 7070 5364
rect 8113 5355 8171 5361
rect 8113 5352 8125 5355
rect 7064 5324 8125 5352
rect 7064 5312 7070 5324
rect 8113 5321 8125 5324
rect 8159 5352 8171 5355
rect 8573 5355 8631 5361
rect 8573 5352 8585 5355
rect 8159 5324 8585 5352
rect 8159 5321 8171 5324
rect 8113 5315 8171 5321
rect 8573 5321 8585 5324
rect 8619 5321 8631 5355
rect 8573 5315 8631 5321
rect 12989 5355 13047 5361
rect 12989 5321 13001 5355
rect 13035 5352 13047 5355
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 13035 5324 13461 5352
rect 13035 5321 13047 5324
rect 12989 5315 13047 5321
rect 13449 5321 13461 5324
rect 13495 5321 13507 5355
rect 13449 5315 13507 5321
rect 15105 5355 15163 5361
rect 15105 5321 15117 5355
rect 15151 5352 15163 5355
rect 15194 5352 15200 5364
rect 15151 5324 15200 5352
rect 15151 5321 15163 5324
rect 15105 5315 15163 5321
rect 3234 5216 3240 5228
rect 3195 5188 3240 5216
rect 3234 5176 3240 5188
rect 3292 5216 3298 5228
rect 7742 5216 7748 5228
rect 3292 5188 5028 5216
rect 3292 5176 3298 5188
rect 2038 5108 2044 5160
rect 2096 5148 2102 5160
rect 2682 5148 2688 5160
rect 2096 5120 2688 5148
rect 2096 5108 2102 5120
rect 2682 5108 2688 5120
rect 2740 5148 2746 5160
rect 5000 5157 5028 5188
rect 7576 5188 7748 5216
rect 2961 5151 3019 5157
rect 2961 5148 2973 5151
rect 2740 5120 2973 5148
rect 2740 5108 2746 5120
rect 2961 5117 2973 5120
rect 3007 5117 3019 5151
rect 2961 5111 3019 5117
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5148 5043 5151
rect 7006 5148 7012 5160
rect 5031 5120 7012 5148
rect 5031 5117 5043 5120
rect 4985 5111 5043 5117
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 7576 5157 7604 5188
rect 7742 5176 7748 5188
rect 7800 5216 7806 5228
rect 8205 5219 8263 5225
rect 8205 5216 8217 5219
rect 7800 5188 8217 5216
rect 7800 5176 7806 5188
rect 8205 5185 8217 5188
rect 8251 5185 8263 5219
rect 9674 5216 9680 5228
rect 8205 5179 8263 5185
rect 8496 5188 9680 5216
rect 7561 5151 7619 5157
rect 7561 5117 7573 5151
rect 7607 5117 7619 5151
rect 7561 5111 7619 5117
rect 8113 5151 8171 5157
rect 8113 5117 8125 5151
rect 8159 5148 8171 5151
rect 8496 5148 8524 5188
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 13004 5216 13032 5315
rect 15194 5312 15200 5324
rect 15252 5312 15258 5364
rect 16942 5352 16948 5364
rect 16903 5324 16948 5352
rect 16942 5312 16948 5324
rect 17000 5312 17006 5364
rect 18046 5352 18052 5364
rect 18007 5324 18052 5352
rect 18046 5312 18052 5324
rect 18104 5312 18110 5364
rect 12268 5188 13032 5216
rect 17589 5219 17647 5225
rect 8159 5120 8524 5148
rect 8573 5151 8631 5157
rect 8159 5117 8171 5120
rect 8113 5111 8171 5117
rect 8573 5117 8585 5151
rect 8619 5148 8631 5151
rect 9122 5148 9128 5160
rect 8619 5120 9128 5148
rect 8619 5117 8631 5120
rect 8573 5111 8631 5117
rect 9122 5108 9128 5120
rect 9180 5108 9186 5160
rect 10318 5148 10324 5160
rect 10279 5120 10324 5148
rect 10318 5108 10324 5120
rect 10376 5108 10382 5160
rect 12268 5157 12296 5188
rect 17589 5185 17601 5219
rect 17635 5216 17647 5219
rect 17954 5216 17960 5228
rect 17635 5188 17960 5216
rect 17635 5185 17647 5188
rect 17589 5179 17647 5185
rect 17954 5176 17960 5188
rect 18012 5176 18018 5228
rect 12253 5151 12311 5157
rect 12253 5117 12265 5151
rect 12299 5117 12311 5151
rect 12253 5111 12311 5117
rect 12342 5108 12348 5160
rect 12400 5148 12406 5160
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 12400 5120 12449 5148
rect 12400 5108 12406 5120
rect 12437 5117 12449 5120
rect 12483 5117 12495 5151
rect 12986 5148 12992 5160
rect 12947 5120 12992 5148
rect 12437 5111 12495 5117
rect 6270 5080 6276 5092
rect 4462 5052 6276 5080
rect 6270 5040 6276 5052
rect 6328 5040 6334 5092
rect 11057 5083 11115 5089
rect 11057 5049 11069 5083
rect 11103 5080 11115 5083
rect 11146 5080 11152 5092
rect 11103 5052 11152 5080
rect 11103 5049 11115 5052
rect 11057 5043 11115 5049
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 11241 5083 11299 5089
rect 11241 5049 11253 5083
rect 11287 5080 11299 5083
rect 11882 5080 11888 5092
rect 11287 5052 11888 5080
rect 11287 5049 11299 5052
rect 11241 5043 11299 5049
rect 11882 5040 11888 5052
rect 11940 5080 11946 5092
rect 12069 5083 12127 5089
rect 12069 5080 12081 5083
rect 11940 5052 12081 5080
rect 11940 5040 11946 5052
rect 12069 5049 12081 5052
rect 12115 5049 12127 5083
rect 12452 5080 12480 5111
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 13081 5151 13139 5157
rect 13081 5117 13093 5151
rect 13127 5117 13139 5151
rect 13081 5111 13139 5117
rect 13449 5151 13507 5157
rect 13449 5117 13461 5151
rect 13495 5148 13507 5151
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 13495 5120 14565 5148
rect 13495 5117 13507 5120
rect 13449 5111 13507 5117
rect 14553 5117 14565 5120
rect 14599 5117 14611 5151
rect 14734 5148 14740 5160
rect 14695 5120 14740 5148
rect 14553 5111 14611 5117
rect 13096 5080 13124 5111
rect 14734 5108 14740 5120
rect 14792 5108 14798 5160
rect 14826 5108 14832 5160
rect 14884 5148 14890 5160
rect 15289 5151 15347 5157
rect 15289 5148 15301 5151
rect 14884 5120 15301 5148
rect 14884 5108 14890 5120
rect 15289 5117 15301 5120
rect 15335 5148 15347 5151
rect 15378 5148 15384 5160
rect 15335 5120 15384 5148
rect 15335 5117 15347 5120
rect 15289 5111 15347 5117
rect 15378 5108 15384 5120
rect 15436 5108 15442 5160
rect 18046 5108 18052 5160
rect 18104 5148 18110 5160
rect 18141 5151 18199 5157
rect 18141 5148 18153 5151
rect 18104 5120 18153 5148
rect 18104 5108 18110 5120
rect 18141 5117 18153 5120
rect 18187 5148 18199 5151
rect 18690 5148 18696 5160
rect 18187 5120 18696 5148
rect 18187 5117 18199 5120
rect 18141 5111 18199 5117
rect 18690 5108 18696 5120
rect 18748 5108 18754 5160
rect 12452 5052 13124 5080
rect 12069 5043 12127 5049
rect 13170 5040 13176 5092
rect 13228 5080 13234 5092
rect 14844 5080 14872 5108
rect 13228 5052 14872 5080
rect 13228 5040 13234 5052
rect 7006 4972 7012 5024
rect 7064 5012 7070 5024
rect 15286 5012 15292 5024
rect 7064 4984 15292 5012
rect 7064 4972 7070 4984
rect 15286 4972 15292 4984
rect 15344 4972 15350 5024
rect 17310 5012 17316 5024
rect 17271 4984 17316 5012
rect 17310 4972 17316 4984
rect 17368 4972 17374 5024
rect 17402 4972 17408 5024
rect 17460 5012 17466 5024
rect 17460 4984 17505 5012
rect 17460 4972 17466 4984
rect 1104 4922 21804 4944
rect 1104 4870 7882 4922
rect 7934 4870 7946 4922
rect 7998 4870 8010 4922
rect 8062 4870 8074 4922
rect 8126 4870 14782 4922
rect 14834 4870 14846 4922
rect 14898 4870 14910 4922
rect 14962 4870 14974 4922
rect 15026 4870 21804 4922
rect 1104 4848 21804 4870
rect 7742 4768 7748 4820
rect 7800 4808 7806 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7800 4780 7849 4808
rect 7800 4768 7806 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 9858 4808 9864 4820
rect 9819 4780 9864 4808
rect 7837 4771 7895 4777
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 10229 4811 10287 4817
rect 10229 4777 10241 4811
rect 10275 4808 10287 4811
rect 12342 4808 12348 4820
rect 10275 4780 12348 4808
rect 10275 4777 10287 4780
rect 10229 4771 10287 4777
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 17310 4768 17316 4820
rect 17368 4808 17374 4820
rect 17957 4811 18015 4817
rect 17957 4808 17969 4811
rect 17368 4780 17969 4808
rect 17368 4768 17374 4780
rect 17957 4777 17969 4780
rect 18003 4777 18015 4811
rect 17957 4771 18015 4777
rect 6270 4700 6276 4752
rect 6328 4740 6334 4752
rect 6822 4740 6828 4752
rect 6328 4712 6828 4740
rect 6328 4700 6334 4712
rect 6822 4700 6828 4712
rect 6880 4700 6886 4752
rect 7374 4700 7380 4752
rect 7432 4740 7438 4752
rect 8205 4743 8263 4749
rect 8205 4740 8217 4743
rect 7432 4712 8217 4740
rect 7432 4700 7438 4712
rect 8205 4709 8217 4712
rect 8251 4709 8263 4743
rect 11146 4740 11152 4752
rect 11107 4712 11152 4740
rect 8205 4703 8263 4709
rect 11146 4700 11152 4712
rect 11204 4700 11210 4752
rect 18417 4743 18475 4749
rect 18417 4709 18429 4743
rect 18463 4740 18475 4743
rect 18966 4740 18972 4752
rect 18463 4712 18972 4740
rect 18463 4709 18475 4712
rect 18417 4703 18475 4709
rect 18966 4700 18972 4712
rect 19024 4700 19030 4752
rect 4982 4672 4988 4684
rect 4895 4644 4988 4672
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 7006 4632 7012 4684
rect 7064 4672 7070 4684
rect 7064 4644 7109 4672
rect 7064 4632 7070 4644
rect 10318 4632 10324 4684
rect 10376 4672 10382 4684
rect 10505 4675 10563 4681
rect 10505 4672 10517 4675
rect 10376 4644 10517 4672
rect 10376 4632 10382 4644
rect 10505 4641 10517 4644
rect 10551 4641 10563 4675
rect 10505 4635 10563 4641
rect 11425 4675 11483 4681
rect 11425 4641 11437 4675
rect 11471 4672 11483 4675
rect 11698 4672 11704 4684
rect 11471 4644 11704 4672
rect 11471 4641 11483 4644
rect 11425 4635 11483 4641
rect 11698 4632 11704 4644
rect 11756 4632 11762 4684
rect 18325 4675 18383 4681
rect 18325 4641 18337 4675
rect 18371 4672 18383 4675
rect 19150 4672 19156 4684
rect 18371 4644 19156 4672
rect 18371 4641 18383 4644
rect 18325 4635 18383 4641
rect 19150 4632 19156 4644
rect 19208 4632 19214 4684
rect 5000 4604 5028 4632
rect 6733 4607 6791 4613
rect 6733 4604 6745 4607
rect 5000 4576 6745 4604
rect 6733 4573 6745 4576
rect 6779 4604 6791 4607
rect 8297 4607 8355 4613
rect 8297 4604 8309 4607
rect 6779 4576 6960 4604
rect 6779 4573 6791 4576
rect 6733 4567 6791 4573
rect 6932 4536 6960 4576
rect 8220 4576 8309 4604
rect 8220 4548 8248 4576
rect 8297 4573 8309 4576
rect 8343 4573 8355 4607
rect 8478 4604 8484 4616
rect 8439 4576 8484 4604
rect 8297 4567 8355 4573
rect 8478 4564 8484 4576
rect 8536 4604 8542 4616
rect 9585 4607 9643 4613
rect 9585 4604 9597 4607
rect 8536 4576 9597 4604
rect 8536 4564 8542 4576
rect 9585 4573 9597 4576
rect 9631 4573 9643 4607
rect 9585 4567 9643 4573
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 9769 4607 9827 4613
rect 9769 4604 9781 4607
rect 9732 4576 9781 4604
rect 9732 4564 9738 4576
rect 9769 4573 9781 4576
rect 9815 4573 9827 4607
rect 18598 4604 18604 4616
rect 18559 4576 18604 4604
rect 9769 4567 9827 4573
rect 18598 4564 18604 4576
rect 18656 4564 18662 4616
rect 7098 4536 7104 4548
rect 6932 4508 7104 4536
rect 7098 4496 7104 4508
rect 7156 4496 7162 4548
rect 8202 4496 8208 4548
rect 8260 4496 8266 4548
rect 1104 4378 21804 4400
rect 1104 4326 4432 4378
rect 4484 4326 4496 4378
rect 4548 4326 4560 4378
rect 4612 4326 4624 4378
rect 4676 4326 11332 4378
rect 11384 4326 11396 4378
rect 11448 4326 11460 4378
rect 11512 4326 11524 4378
rect 11576 4326 18232 4378
rect 18284 4326 18296 4378
rect 18348 4326 18360 4378
rect 18412 4326 18424 4378
rect 18476 4326 21804 4378
rect 1104 4304 21804 4326
rect 7098 4224 7104 4276
rect 7156 4264 7162 4276
rect 16942 4264 16948 4276
rect 7156 4236 16948 4264
rect 7156 4224 7162 4236
rect 16942 4224 16948 4236
rect 17000 4264 17006 4276
rect 17402 4264 17408 4276
rect 17000 4236 17408 4264
rect 17000 4224 17006 4236
rect 17402 4224 17408 4236
rect 17460 4224 17466 4276
rect 15378 4196 15384 4208
rect 15339 4168 15384 4196
rect 15378 4156 15384 4168
rect 15436 4156 15442 4208
rect 18966 4156 18972 4208
rect 19024 4196 19030 4208
rect 21082 4196 21088 4208
rect 19024 4168 21088 4196
rect 19024 4156 19030 4168
rect 21082 4156 21088 4168
rect 21140 4156 21146 4208
rect 15102 3952 15108 4004
rect 15160 3992 15166 4004
rect 15565 3995 15623 4001
rect 15565 3992 15577 3995
rect 15160 3964 15577 3992
rect 15160 3952 15166 3964
rect 15565 3961 15577 3964
rect 15611 3961 15623 3995
rect 15565 3955 15623 3961
rect 7558 3884 7564 3936
rect 7616 3924 7622 3936
rect 11974 3924 11980 3936
rect 7616 3896 11980 3924
rect 7616 3884 7622 3896
rect 11974 3884 11980 3896
rect 12032 3884 12038 3936
rect 1104 3834 21804 3856
rect 1104 3782 7882 3834
rect 7934 3782 7946 3834
rect 7998 3782 8010 3834
rect 8062 3782 8074 3834
rect 8126 3782 14782 3834
rect 14834 3782 14846 3834
rect 14898 3782 14910 3834
rect 14962 3782 14974 3834
rect 15026 3782 21804 3834
rect 1104 3760 21804 3782
rect 8849 3723 8907 3729
rect 8849 3689 8861 3723
rect 8895 3720 8907 3723
rect 9309 3723 9367 3729
rect 9309 3720 9321 3723
rect 8895 3692 9321 3720
rect 8895 3689 8907 3692
rect 8849 3683 8907 3689
rect 9309 3689 9321 3692
rect 9355 3720 9367 3723
rect 9490 3720 9496 3732
rect 9355 3692 9496 3720
rect 9355 3689 9367 3692
rect 9309 3683 9367 3689
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 11333 3723 11391 3729
rect 11333 3720 11345 3723
rect 11204 3692 11345 3720
rect 11204 3680 11210 3692
rect 11333 3689 11345 3692
rect 11379 3720 11391 3723
rect 11425 3723 11483 3729
rect 11425 3720 11437 3723
rect 11379 3692 11437 3720
rect 11379 3689 11391 3692
rect 11333 3683 11391 3689
rect 11425 3689 11437 3692
rect 11471 3689 11483 3723
rect 11425 3683 11483 3689
rect 13909 3723 13967 3729
rect 13909 3689 13921 3723
rect 13955 3720 13967 3723
rect 14458 3720 14464 3732
rect 13955 3692 14464 3720
rect 13955 3689 13967 3692
rect 13909 3683 13967 3689
rect 14458 3680 14464 3692
rect 14516 3720 14522 3732
rect 14829 3723 14887 3729
rect 14829 3720 14841 3723
rect 14516 3692 14841 3720
rect 14516 3680 14522 3692
rect 14829 3689 14841 3692
rect 14875 3689 14887 3723
rect 15102 3720 15108 3732
rect 15063 3692 15108 3720
rect 14829 3683 14887 3689
rect 15102 3680 15108 3692
rect 15160 3680 15166 3732
rect 3970 3652 3976 3664
rect 3931 3624 3976 3652
rect 3970 3612 3976 3624
rect 4028 3612 4034 3664
rect 9122 3652 9128 3664
rect 9083 3624 9128 3652
rect 9122 3612 9128 3624
rect 9180 3612 9186 3664
rect 11609 3655 11667 3661
rect 11609 3621 11621 3655
rect 11655 3652 11667 3655
rect 11698 3652 11704 3664
rect 11655 3624 11704 3652
rect 11655 3621 11667 3624
rect 11609 3615 11667 3621
rect 11698 3612 11704 3624
rect 11756 3612 11762 3664
rect 17954 3652 17960 3664
rect 12406 3624 17960 3652
rect 6730 3584 6736 3596
rect 6691 3556 6736 3584
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 6822 3544 6828 3596
rect 6880 3584 6886 3596
rect 7009 3587 7067 3593
rect 7009 3584 7021 3587
rect 6880 3556 7021 3584
rect 6880 3544 6886 3556
rect 7009 3553 7021 3556
rect 7055 3584 7067 3587
rect 11882 3584 11888 3596
rect 7055 3556 11100 3584
rect 11843 3556 11888 3584
rect 7055 3553 7067 3556
rect 7009 3547 7067 3553
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3516 8539 3519
rect 9030 3516 9036 3528
rect 8527 3488 9036 3516
rect 8527 3485 8539 3488
rect 8481 3479 8539 3485
rect 9030 3476 9036 3488
rect 9088 3476 9094 3528
rect 10962 3516 10968 3528
rect 10923 3488 10968 3516
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11072 3516 11100 3556
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 12406 3516 12434 3624
rect 17954 3612 17960 3624
rect 18012 3612 18018 3664
rect 15013 3587 15071 3593
rect 15013 3553 15025 3587
rect 15059 3584 15071 3587
rect 15105 3587 15163 3593
rect 15105 3584 15117 3587
rect 15059 3556 15117 3584
rect 15059 3553 15071 3556
rect 15013 3547 15071 3553
rect 15105 3553 15117 3556
rect 15151 3553 15163 3587
rect 15105 3547 15163 3553
rect 11072 3488 12434 3516
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13814 3516 13820 3528
rect 13587 3488 13820 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 15473 3519 15531 3525
rect 15473 3485 15485 3519
rect 15519 3516 15531 3519
rect 15562 3516 15568 3528
rect 15519 3488 15568 3516
rect 15519 3485 15531 3488
rect 15473 3479 15531 3485
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 4157 3451 4215 3457
rect 4157 3417 4169 3451
rect 4203 3448 4215 3451
rect 8849 3451 8907 3457
rect 4203 3420 8800 3448
rect 4203 3417 4215 3420
rect 4157 3411 4215 3417
rect 8772 3380 8800 3420
rect 8849 3417 8861 3451
rect 8895 3448 8907 3451
rect 9766 3448 9772 3460
rect 8895 3420 9772 3448
rect 8895 3417 8907 3420
rect 8849 3411 8907 3417
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 11333 3451 11391 3457
rect 11333 3417 11345 3451
rect 11379 3448 11391 3451
rect 11701 3451 11759 3457
rect 11701 3448 11713 3451
rect 11379 3420 11713 3448
rect 11379 3417 11391 3420
rect 11333 3411 11391 3417
rect 11701 3417 11713 3420
rect 11747 3417 11759 3451
rect 11701 3411 11759 3417
rect 13909 3451 13967 3457
rect 13909 3417 13921 3451
rect 13955 3448 13967 3451
rect 14550 3448 14556 3460
rect 13955 3420 14556 3448
rect 13955 3417 13967 3420
rect 13909 3411 13967 3417
rect 14550 3408 14556 3420
rect 14608 3408 14614 3460
rect 11790 3380 11796 3392
rect 8772 3352 11796 3380
rect 11790 3340 11796 3352
rect 11848 3340 11854 3392
rect 11974 3340 11980 3392
rect 12032 3380 12038 3392
rect 15930 3380 15936 3392
rect 12032 3352 15936 3380
rect 12032 3340 12038 3352
rect 15930 3340 15936 3352
rect 15988 3340 15994 3392
rect 1104 3290 21804 3312
rect 1104 3238 4432 3290
rect 4484 3238 4496 3290
rect 4548 3238 4560 3290
rect 4612 3238 4624 3290
rect 4676 3238 11332 3290
rect 11384 3238 11396 3290
rect 11448 3238 11460 3290
rect 11512 3238 11524 3290
rect 11576 3238 18232 3290
rect 18284 3238 18296 3290
rect 18348 3238 18360 3290
rect 18412 3238 18424 3290
rect 18476 3238 21804 3290
rect 1104 3216 21804 3238
rect 9030 3176 9036 3188
rect 8991 3148 9036 3176
rect 9030 3136 9036 3148
rect 9088 3136 9094 3188
rect 9766 3176 9772 3188
rect 9727 3148 9772 3176
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 11146 3136 11152 3188
rect 11204 3176 11210 3188
rect 11425 3179 11483 3185
rect 11425 3176 11437 3179
rect 11204 3148 11437 3176
rect 11204 3136 11210 3148
rect 11425 3145 11437 3148
rect 11471 3145 11483 3179
rect 11425 3139 11483 3145
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 12621 3179 12679 3185
rect 12621 3176 12633 3179
rect 12492 3148 12633 3176
rect 12492 3136 12498 3148
rect 12621 3145 12633 3148
rect 12667 3145 12679 3179
rect 13814 3176 13820 3188
rect 13775 3148 13820 3176
rect 12621 3139 12679 3145
rect 13814 3136 13820 3148
rect 13872 3136 13878 3188
rect 14550 3176 14556 3188
rect 14511 3148 14556 3176
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 14921 3179 14979 3185
rect 14921 3145 14933 3179
rect 14967 3176 14979 3179
rect 15102 3176 15108 3188
rect 14967 3148 15108 3176
rect 14967 3145 14979 3148
rect 14921 3139 14979 3145
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 15562 3176 15568 3188
rect 15523 3148 15568 3176
rect 15562 3136 15568 3148
rect 15620 3136 15626 3188
rect 17208 3179 17266 3185
rect 17208 3145 17220 3179
rect 17254 3176 17266 3179
rect 18966 3176 18972 3188
rect 17254 3148 18972 3176
rect 17254 3145 17266 3148
rect 17208 3139 17266 3145
rect 18966 3136 18972 3148
rect 19024 3136 19030 3188
rect 19150 3176 19156 3188
rect 19111 3148 19156 3176
rect 19150 3136 19156 3148
rect 19208 3136 19214 3188
rect 8478 3040 8484 3052
rect 8439 3012 8484 3040
rect 8478 3000 8484 3012
rect 8536 3000 8542 3052
rect 1394 2972 1400 2984
rect 1355 2944 1400 2972
rect 1394 2932 1400 2944
rect 1452 2932 1458 2984
rect 8496 2904 8524 3000
rect 8665 2975 8723 2981
rect 8665 2941 8677 2975
rect 8711 2972 8723 2975
rect 8938 2972 8944 2984
rect 8711 2944 8944 2972
rect 8711 2941 8723 2944
rect 8665 2935 8723 2941
rect 8938 2932 8944 2944
rect 8996 2932 9002 2984
rect 9048 2972 9076 3136
rect 14458 3108 14464 3120
rect 10428 3080 12296 3108
rect 14419 3080 14464 3108
rect 9490 3040 9496 3052
rect 9451 3012 9496 3040
rect 9490 3000 9496 3012
rect 9548 3000 9554 3052
rect 9125 2975 9183 2981
rect 9125 2972 9137 2975
rect 9048 2944 9137 2972
rect 9125 2941 9137 2944
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 9677 2975 9735 2981
rect 9677 2941 9689 2975
rect 9723 2972 9735 2975
rect 9858 2972 9864 2984
rect 9723 2944 9864 2972
rect 9723 2941 9735 2944
rect 9677 2935 9735 2941
rect 9858 2932 9864 2944
rect 9916 2972 9922 2984
rect 9953 2975 10011 2981
rect 9953 2972 9965 2975
rect 9916 2944 9965 2972
rect 9916 2932 9922 2944
rect 9953 2941 9965 2944
rect 9999 2941 10011 2975
rect 9953 2935 10011 2941
rect 10428 2904 10456 3080
rect 10502 3000 10508 3052
rect 10560 3040 10566 3052
rect 12268 3049 12296 3080
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 12253 3043 12311 3049
rect 10560 3012 12112 3040
rect 10560 3000 10566 3012
rect 10873 2975 10931 2981
rect 10873 2941 10885 2975
rect 10919 2972 10931 2975
rect 10962 2972 10968 2984
rect 10919 2944 10968 2972
rect 10919 2941 10931 2944
rect 10873 2935 10931 2941
rect 8496 2876 10456 2904
rect 10888 2904 10916 2935
rect 10962 2932 10968 2944
rect 11020 2932 11026 2984
rect 11425 2975 11483 2981
rect 11425 2941 11437 2975
rect 11471 2972 11483 2975
rect 11882 2972 11888 2984
rect 11471 2944 11888 2972
rect 11471 2941 11483 2944
rect 11425 2935 11483 2941
rect 11882 2932 11888 2944
rect 11940 2932 11946 2984
rect 12084 2981 12112 3012
rect 12253 3009 12265 3043
rect 12299 3040 12311 3043
rect 13265 3043 13323 3049
rect 13265 3040 13277 3043
rect 12299 3012 13277 3040
rect 12299 3009 12311 3012
rect 12253 3003 12311 3009
rect 13265 3009 13277 3012
rect 13311 3040 13323 3043
rect 13311 3012 15056 3040
rect 13311 3009 13323 3012
rect 13265 3003 13323 3009
rect 12069 2975 12127 2981
rect 12069 2941 12081 2975
rect 12115 2941 12127 2975
rect 12526 2972 12532 2984
rect 12487 2944 12532 2972
rect 12069 2935 12127 2941
rect 12526 2932 12532 2944
rect 12584 2932 12590 2984
rect 13446 2972 13452 2984
rect 13407 2944 13452 2972
rect 13446 2932 13452 2944
rect 13504 2932 13510 2984
rect 13814 2932 13820 2984
rect 13872 2972 13878 2984
rect 13909 2975 13967 2981
rect 13909 2972 13921 2975
rect 13872 2944 13921 2972
rect 13872 2932 13878 2944
rect 13909 2941 13921 2944
rect 13955 2941 13967 2975
rect 13909 2935 13967 2941
rect 14461 2975 14519 2981
rect 14461 2941 14473 2975
rect 14507 2972 14519 2975
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 14507 2944 14749 2972
rect 14507 2941 14519 2944
rect 14461 2935 14519 2941
rect 14737 2941 14749 2944
rect 14783 2972 14795 2975
rect 14921 2975 14979 2981
rect 14921 2972 14933 2975
rect 14783 2944 14933 2972
rect 14783 2941 14795 2944
rect 14737 2935 14795 2941
rect 14921 2941 14933 2944
rect 14967 2941 14979 2975
rect 14921 2935 14979 2941
rect 10888 2876 11744 2904
rect 11716 2845 11744 2876
rect 11790 2864 11796 2916
rect 11848 2904 11854 2916
rect 14476 2904 14504 2935
rect 11848 2876 14504 2904
rect 15028 2904 15056 3012
rect 15473 2975 15531 2981
rect 15473 2941 15485 2975
rect 15519 2972 15531 2975
rect 15580 2972 15608 3136
rect 16114 3040 16120 3052
rect 16075 3012 16120 3040
rect 16114 3000 16120 3012
rect 16172 3000 16178 3052
rect 16942 3040 16948 3052
rect 16903 3012 16948 3040
rect 16942 3000 16948 3012
rect 17000 3000 17006 3052
rect 17954 3000 17960 3052
rect 18012 3040 18018 3052
rect 19168 3040 19196 3136
rect 20898 3040 20904 3052
rect 18012 3012 18460 3040
rect 19168 3012 20904 3040
rect 18012 3000 18018 3012
rect 15930 2972 15936 2984
rect 15519 2944 15608 2972
rect 15891 2944 15936 2972
rect 15519 2941 15531 2944
rect 15473 2935 15531 2941
rect 15930 2932 15936 2944
rect 15988 2932 15994 2984
rect 16114 2904 16120 2916
rect 15028 2876 16120 2904
rect 11848 2864 11854 2876
rect 16114 2864 16120 2876
rect 16172 2864 16178 2916
rect 18432 2904 18460 3012
rect 20898 3000 20904 3012
rect 20956 3000 20962 3052
rect 21174 3040 21180 3052
rect 21135 3012 21180 3040
rect 21174 3000 21180 3012
rect 21232 3000 21238 3052
rect 18966 2972 18972 2984
rect 18927 2944 18972 2972
rect 18966 2932 18972 2944
rect 19024 2932 19030 2984
rect 21450 2972 21456 2984
rect 21411 2944 21456 2972
rect 21450 2932 21456 2944
rect 21508 2932 21514 2984
rect 18432 2890 19734 2904
rect 18446 2876 19734 2890
rect 1581 2839 1639 2845
rect 1581 2805 1593 2839
rect 1627 2836 1639 2839
rect 8573 2839 8631 2845
rect 8573 2836 8585 2839
rect 1627 2808 8585 2836
rect 1627 2805 1639 2808
rect 1581 2799 1639 2805
rect 8573 2805 8585 2808
rect 8619 2805 8631 2839
rect 8573 2799 8631 2805
rect 11701 2839 11759 2845
rect 11701 2805 11713 2839
rect 11747 2805 11759 2839
rect 12158 2836 12164 2848
rect 12119 2808 12164 2836
rect 11701 2799 11759 2805
rect 12158 2796 12164 2808
rect 12216 2796 12222 2848
rect 13357 2839 13415 2845
rect 13357 2805 13369 2839
rect 13403 2836 13415 2839
rect 13814 2836 13820 2848
rect 13403 2808 13820 2836
rect 13403 2805 13415 2808
rect 13357 2799 13415 2805
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 16025 2839 16083 2845
rect 16025 2805 16037 2839
rect 16071 2836 16083 2839
rect 21269 2839 21327 2845
rect 21269 2836 21281 2839
rect 16071 2808 21281 2836
rect 16071 2805 16083 2808
rect 16025 2799 16083 2805
rect 21269 2805 21281 2808
rect 21315 2805 21327 2839
rect 21269 2799 21327 2805
rect 1104 2746 21804 2768
rect 1104 2694 7882 2746
rect 7934 2694 7946 2746
rect 7998 2694 8010 2746
rect 8062 2694 8074 2746
rect 8126 2694 14782 2746
rect 14834 2694 14846 2746
rect 14898 2694 14910 2746
rect 14962 2694 14974 2746
rect 15026 2694 21804 2746
rect 1104 2672 21804 2694
rect 4065 2635 4123 2641
rect 4065 2601 4077 2635
rect 4111 2632 4123 2635
rect 4798 2632 4804 2644
rect 4111 2604 4804 2632
rect 4111 2601 4123 2604
rect 4065 2595 4123 2601
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 5721 2635 5779 2641
rect 5721 2601 5733 2635
rect 5767 2632 5779 2635
rect 6638 2632 6644 2644
rect 5767 2604 6644 2632
rect 5767 2601 5779 2604
rect 5721 2595 5779 2601
rect 6638 2592 6644 2604
rect 6696 2592 6702 2644
rect 6730 2592 6736 2644
rect 6788 2632 6794 2644
rect 7009 2635 7067 2641
rect 7009 2632 7021 2635
rect 6788 2604 7021 2632
rect 6788 2592 6794 2604
rect 7009 2601 7021 2604
rect 7055 2601 7067 2635
rect 7009 2595 7067 2601
rect 8941 2635 8999 2641
rect 8941 2601 8953 2635
rect 8987 2632 8999 2635
rect 9674 2632 9680 2644
rect 8987 2604 9680 2632
rect 8987 2601 8999 2604
rect 8941 2595 8999 2601
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 12158 2632 12164 2644
rect 12119 2604 12164 2632
rect 12158 2592 12164 2604
rect 12216 2592 12222 2644
rect 13814 2632 13820 2644
rect 13775 2604 13820 2632
rect 13814 2592 13820 2604
rect 13872 2592 13878 2644
rect 17405 2635 17463 2641
rect 17405 2601 17417 2635
rect 17451 2632 17463 2635
rect 17494 2632 17500 2644
rect 17451 2604 17500 2632
rect 17451 2601 17463 2604
rect 17405 2595 17463 2601
rect 17494 2592 17500 2604
rect 17552 2592 17558 2644
rect 18874 2632 18880 2644
rect 18835 2604 18880 2632
rect 18874 2592 18880 2604
rect 18932 2592 18938 2644
rect 21269 2635 21327 2641
rect 21269 2601 21281 2635
rect 21315 2601 21327 2635
rect 21269 2595 21327 2601
rect 2038 2564 2044 2576
rect 1999 2536 2044 2564
rect 2038 2524 2044 2536
rect 2096 2524 2102 2576
rect 8202 2524 8208 2576
rect 8260 2564 8266 2576
rect 21284 2564 21312 2595
rect 8260 2536 21312 2564
rect 8260 2524 8266 2536
rect 474 2456 480 2508
rect 532 2496 538 2508
rect 1397 2499 1455 2505
rect 1397 2496 1409 2499
rect 532 2468 1409 2496
rect 532 2456 538 2468
rect 1397 2465 1409 2468
rect 1443 2465 1455 2499
rect 1397 2459 1455 2465
rect 3694 2456 3700 2508
rect 3752 2496 3758 2508
rect 3881 2499 3939 2505
rect 3881 2496 3893 2499
rect 3752 2468 3893 2496
rect 3752 2456 3758 2468
rect 3881 2465 3893 2468
rect 3927 2465 3939 2499
rect 5534 2496 5540 2508
rect 5495 2468 5540 2496
rect 3881 2459 3939 2465
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 7101 2499 7159 2505
rect 7101 2496 7113 2499
rect 6972 2468 7113 2496
rect 6972 2456 6978 2468
rect 7101 2465 7113 2468
rect 7147 2465 7159 2499
rect 8754 2496 8760 2508
rect 8715 2468 8760 2496
rect 7101 2459 7159 2465
rect 8754 2456 8760 2468
rect 8812 2456 8818 2508
rect 10594 2456 10600 2508
rect 10652 2496 10658 2508
rect 10689 2499 10747 2505
rect 10689 2496 10701 2499
rect 10652 2468 10701 2496
rect 10652 2456 10658 2468
rect 10689 2465 10701 2468
rect 10735 2465 10747 2499
rect 11974 2496 11980 2508
rect 11935 2468 11980 2496
rect 10689 2459 10747 2465
rect 11974 2456 11980 2468
rect 12032 2456 12038 2508
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 14001 2499 14059 2505
rect 14001 2496 14013 2499
rect 13872 2468 14013 2496
rect 13872 2456 13878 2468
rect 14001 2465 14013 2468
rect 14047 2465 14059 2499
rect 15654 2496 15660 2508
rect 15615 2468 15660 2496
rect 14001 2459 14059 2465
rect 15654 2456 15660 2468
rect 15712 2456 15718 2508
rect 17034 2456 17040 2508
rect 17092 2496 17098 2508
rect 17313 2499 17371 2505
rect 17313 2496 17325 2499
rect 17092 2468 17325 2496
rect 17092 2456 17098 2468
rect 17313 2465 17325 2468
rect 17359 2465 17371 2499
rect 17313 2459 17371 2465
rect 18874 2456 18880 2508
rect 18932 2496 18938 2508
rect 19061 2499 19119 2505
rect 19061 2496 19073 2499
rect 18932 2468 19073 2496
rect 18932 2456 18938 2468
rect 19061 2465 19073 2468
rect 19107 2465 19119 2499
rect 20898 2496 20904 2508
rect 20859 2468 20904 2496
rect 19061 2459 19119 2465
rect 20898 2456 20904 2468
rect 20956 2456 20962 2508
rect 21453 2499 21511 2505
rect 21453 2465 21465 2499
rect 21499 2496 21511 2499
rect 22094 2496 22100 2508
rect 21499 2468 22100 2496
rect 21499 2465 21511 2468
rect 21453 2459 21511 2465
rect 22094 2456 22100 2468
rect 22152 2456 22158 2508
rect 12526 2428 12532 2440
rect 1596 2400 12532 2428
rect 1596 2369 1624 2400
rect 12526 2388 12532 2400
rect 12584 2388 12590 2440
rect 16114 2428 16120 2440
rect 16075 2400 16120 2428
rect 16114 2388 16120 2400
rect 16172 2388 16178 2440
rect 1581 2363 1639 2369
rect 1581 2329 1593 2363
rect 1627 2329 1639 2363
rect 1854 2360 1860 2372
rect 1815 2332 1860 2360
rect 1581 2323 1639 2329
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 10873 2363 10931 2369
rect 10873 2329 10885 2363
rect 10919 2360 10931 2363
rect 18046 2360 18052 2372
rect 10919 2332 18052 2360
rect 10919 2329 10931 2332
rect 10873 2323 10931 2329
rect 18046 2320 18052 2332
rect 18104 2320 18110 2372
rect 20714 2360 20720 2372
rect 20675 2332 20720 2360
rect 20714 2320 20720 2332
rect 20772 2320 20778 2372
rect 1104 2202 21804 2224
rect 1104 2150 4432 2202
rect 4484 2150 4496 2202
rect 4548 2150 4560 2202
rect 4612 2150 4624 2202
rect 4676 2150 11332 2202
rect 11384 2150 11396 2202
rect 11448 2150 11460 2202
rect 11512 2150 11524 2202
rect 11576 2150 18232 2202
rect 18284 2150 18296 2202
rect 18348 2150 18360 2202
rect 18412 2150 18424 2202
rect 18476 2150 21804 2202
rect 1104 2128 21804 2150
<< via1 >>
rect 4432 22822 4484 22874
rect 4496 22822 4548 22874
rect 4560 22822 4612 22874
rect 4624 22822 4676 22874
rect 11332 22822 11384 22874
rect 11396 22822 11448 22874
rect 11460 22822 11512 22874
rect 11524 22822 11576 22874
rect 18232 22822 18284 22874
rect 18296 22822 18348 22874
rect 18360 22822 18412 22874
rect 18424 22822 18476 22874
rect 1492 22763 1544 22772
rect 1492 22729 1501 22763
rect 1501 22729 1535 22763
rect 1535 22729 1544 22763
rect 1492 22720 1544 22729
rect 4896 22652 4948 22704
rect 11796 22652 11848 22704
rect 940 22516 992 22568
rect 2780 22559 2832 22568
rect 2780 22525 2789 22559
rect 2789 22525 2823 22559
rect 2823 22525 2832 22559
rect 2780 22516 2832 22525
rect 4804 22516 4856 22568
rect 6000 22559 6052 22568
rect 6000 22525 6009 22559
rect 6009 22525 6043 22559
rect 6043 22525 6052 22559
rect 6000 22516 6052 22525
rect 7840 22559 7892 22568
rect 7840 22525 7849 22559
rect 7849 22525 7883 22559
rect 7883 22525 7892 22559
rect 7840 22516 7892 22525
rect 9680 22559 9732 22568
rect 9680 22525 9689 22559
rect 9689 22525 9723 22559
rect 9723 22525 9732 22559
rect 9680 22516 9732 22525
rect 11704 22559 11756 22568
rect 11704 22525 11713 22559
rect 11713 22525 11747 22559
rect 11747 22525 11756 22559
rect 11704 22516 11756 22525
rect 12900 22559 12952 22568
rect 12900 22525 12909 22559
rect 12909 22525 12943 22559
rect 12943 22525 12952 22559
rect 12900 22516 12952 22525
rect 14740 22516 14792 22568
rect 16580 22516 16632 22568
rect 17960 22516 18012 22568
rect 19800 22516 19852 22568
rect 21088 22559 21140 22568
rect 21088 22525 21097 22559
rect 21097 22525 21131 22559
rect 21131 22525 21140 22559
rect 21088 22516 21140 22525
rect 21640 22516 21692 22568
rect 1584 22491 1636 22500
rect 1584 22457 1593 22491
rect 1593 22457 1627 22491
rect 1627 22457 1636 22491
rect 1584 22448 1636 22457
rect 2044 22380 2096 22432
rect 4804 22423 4856 22432
rect 4804 22389 4813 22423
rect 4813 22389 4847 22423
rect 4847 22389 4856 22423
rect 4804 22380 4856 22389
rect 6368 22380 6420 22432
rect 9680 22380 9732 22432
rect 11152 22380 11204 22432
rect 13084 22423 13136 22432
rect 13084 22389 13093 22423
rect 13093 22389 13127 22423
rect 13127 22389 13136 22423
rect 13084 22380 13136 22389
rect 14556 22380 14608 22432
rect 16764 22380 16816 22432
rect 17960 22423 18012 22432
rect 17960 22389 17969 22423
rect 17969 22389 18003 22423
rect 18003 22389 18012 22423
rect 17960 22380 18012 22389
rect 19616 22380 19668 22432
rect 20904 22423 20956 22432
rect 20904 22389 20913 22423
rect 20913 22389 20947 22423
rect 20947 22389 20956 22423
rect 20904 22380 20956 22389
rect 20996 22380 21048 22432
rect 7882 22278 7934 22330
rect 7946 22278 7998 22330
rect 8010 22278 8062 22330
rect 8074 22278 8126 22330
rect 14782 22278 14834 22330
rect 14846 22278 14898 22330
rect 14910 22278 14962 22330
rect 14974 22278 15026 22330
rect 15476 22176 15528 22228
rect 20904 22176 20956 22228
rect 3700 22040 3752 22092
rect 5264 22040 5316 22092
rect 5540 22040 5592 22092
rect 10324 22040 10376 22092
rect 11704 22083 11756 22092
rect 11704 22049 11713 22083
rect 11713 22049 11747 22083
rect 11747 22049 11756 22083
rect 11704 22040 11756 22049
rect 11888 22083 11940 22092
rect 11888 22049 11897 22083
rect 11897 22049 11931 22083
rect 11931 22049 11940 22083
rect 11888 22040 11940 22049
rect 11980 22083 12032 22092
rect 11980 22049 11989 22083
rect 11989 22049 12023 22083
rect 12023 22049 12032 22083
rect 11980 22040 12032 22049
rect 12348 22040 12400 22092
rect 5816 21972 5868 22024
rect 17132 22040 17184 22092
rect 4160 21836 4212 21888
rect 4988 21836 5040 21888
rect 5448 21879 5500 21888
rect 5448 21845 5457 21879
rect 5457 21845 5491 21879
rect 5491 21845 5500 21879
rect 5448 21836 5500 21845
rect 7656 21836 7708 21888
rect 10048 21879 10100 21888
rect 10048 21845 10057 21879
rect 10057 21845 10091 21879
rect 10091 21845 10100 21879
rect 10048 21836 10100 21845
rect 12072 21836 12124 21888
rect 12808 21836 12860 21888
rect 15292 21836 15344 21888
rect 18696 21836 18748 21888
rect 20168 21879 20220 21888
rect 20168 21845 20177 21879
rect 20177 21845 20211 21879
rect 20211 21845 20220 21879
rect 20168 21836 20220 21845
rect 4432 21734 4484 21786
rect 4496 21734 4548 21786
rect 4560 21734 4612 21786
rect 4624 21734 4676 21786
rect 11332 21734 11384 21786
rect 11396 21734 11448 21786
rect 11460 21734 11512 21786
rect 11524 21734 11576 21786
rect 18232 21734 18284 21786
rect 18296 21734 18348 21786
rect 18360 21734 18412 21786
rect 18424 21734 18476 21786
rect 1584 21632 1636 21684
rect 5540 21632 5592 21684
rect 5816 21675 5868 21684
rect 4160 21539 4212 21548
rect 4160 21505 4169 21539
rect 4169 21505 4203 21539
rect 4203 21505 4212 21539
rect 4160 21496 4212 21505
rect 2504 21428 2556 21480
rect 5816 21641 5825 21675
rect 5825 21641 5859 21675
rect 5859 21641 5868 21675
rect 5816 21632 5868 21641
rect 9036 21539 9088 21548
rect 9036 21505 9045 21539
rect 9045 21505 9079 21539
rect 9079 21505 9088 21539
rect 9036 21496 9088 21505
rect 12072 21539 12124 21548
rect 12072 21505 12081 21539
rect 12081 21505 12115 21539
rect 12115 21505 12124 21539
rect 12072 21496 12124 21505
rect 16580 21632 16632 21684
rect 15108 21496 15160 21548
rect 16580 21496 16632 21548
rect 17776 21496 17828 21548
rect 5448 21360 5500 21412
rect 7196 21360 7248 21412
rect 7656 21360 7708 21412
rect 10048 21360 10100 21412
rect 7748 21292 7800 21344
rect 9036 21292 9088 21344
rect 17132 21471 17184 21480
rect 17132 21437 17141 21471
rect 17141 21437 17175 21471
rect 17175 21437 17184 21471
rect 17132 21428 17184 21437
rect 11244 21403 11296 21412
rect 11244 21369 11253 21403
rect 11253 21369 11287 21403
rect 11287 21369 11296 21403
rect 11244 21360 11296 21369
rect 12808 21360 12860 21412
rect 14648 21360 14700 21412
rect 15292 21360 15344 21412
rect 17960 21360 18012 21412
rect 18696 21360 18748 21412
rect 20168 21360 20220 21412
rect 11888 21292 11940 21344
rect 13544 21335 13596 21344
rect 13544 21301 13553 21335
rect 13553 21301 13587 21335
rect 13587 21301 13596 21335
rect 13544 21292 13596 21301
rect 17224 21292 17276 21344
rect 20904 21292 20956 21344
rect 7882 21190 7934 21242
rect 7946 21190 7998 21242
rect 8010 21190 8062 21242
rect 8074 21190 8126 21242
rect 14782 21190 14834 21242
rect 14846 21190 14898 21242
rect 14910 21190 14962 21242
rect 14974 21190 15026 21242
rect 7196 21131 7248 21140
rect 7196 21097 7205 21131
rect 7205 21097 7239 21131
rect 7239 21097 7248 21131
rect 7196 21088 7248 21097
rect 7472 21063 7524 21072
rect 7472 21029 7481 21063
rect 7481 21029 7515 21063
rect 7515 21029 7524 21063
rect 7472 21020 7524 21029
rect 8300 21088 8352 21140
rect 11980 21088 12032 21140
rect 14648 21131 14700 21140
rect 7748 21020 7800 21072
rect 14648 21097 14657 21131
rect 14657 21097 14691 21131
rect 14691 21097 14700 21131
rect 14648 21088 14700 21097
rect 12624 21020 12676 21072
rect 13544 21020 13596 21072
rect 15108 21020 15160 21072
rect 7380 20995 7432 21004
rect 7380 20961 7389 20995
rect 7389 20961 7423 20995
rect 7423 20961 7432 20995
rect 7380 20952 7432 20961
rect 8852 20952 8904 21004
rect 11244 20952 11296 21004
rect 11704 20952 11756 21004
rect 11980 20995 12032 21004
rect 11980 20961 11989 20995
rect 11989 20961 12023 20995
rect 12023 20961 12032 20995
rect 11980 20952 12032 20961
rect 12164 20995 12216 21004
rect 12164 20961 12173 20995
rect 12173 20961 12207 20995
rect 12207 20961 12216 20995
rect 12348 20995 12400 21004
rect 12164 20952 12216 20961
rect 12348 20961 12357 20995
rect 12357 20961 12391 20995
rect 12391 20961 12400 20995
rect 12348 20952 12400 20961
rect 15200 20995 15252 21004
rect 15200 20961 15209 20995
rect 15209 20961 15243 20995
rect 15243 20961 15252 20995
rect 15200 20952 15252 20961
rect 16580 21020 16632 21072
rect 17224 21020 17276 21072
rect 21088 20952 21140 21004
rect 15384 20884 15436 20936
rect 16488 20927 16540 20936
rect 16488 20893 16497 20927
rect 16497 20893 16531 20927
rect 16531 20893 16540 20927
rect 16488 20884 16540 20893
rect 15844 20816 15896 20868
rect 8300 20791 8352 20800
rect 8300 20757 8309 20791
rect 8309 20757 8343 20791
rect 8343 20757 8352 20791
rect 8300 20748 8352 20757
rect 9312 20748 9364 20800
rect 11060 20748 11112 20800
rect 15384 20748 15436 20800
rect 21364 20791 21416 20800
rect 21364 20757 21373 20791
rect 21373 20757 21407 20791
rect 21407 20757 21416 20791
rect 21364 20748 21416 20757
rect 4432 20646 4484 20698
rect 4496 20646 4548 20698
rect 4560 20646 4612 20698
rect 4624 20646 4676 20698
rect 11332 20646 11384 20698
rect 11396 20646 11448 20698
rect 11460 20646 11512 20698
rect 11524 20646 11576 20698
rect 18232 20646 18284 20698
rect 18296 20646 18348 20698
rect 18360 20646 18412 20698
rect 18424 20646 18476 20698
rect 11980 20476 12032 20528
rect 9036 20408 9088 20460
rect 11060 20408 11112 20460
rect 1400 20383 1452 20392
rect 1400 20349 1409 20383
rect 1409 20349 1443 20383
rect 1443 20349 1452 20383
rect 1400 20340 1452 20349
rect 2504 20383 2556 20392
rect 2504 20349 2513 20383
rect 2513 20349 2547 20383
rect 2547 20349 2556 20383
rect 2504 20340 2556 20349
rect 1492 20204 1544 20256
rect 3516 20272 3568 20324
rect 5540 20340 5592 20392
rect 11888 20383 11940 20392
rect 11888 20349 11897 20383
rect 11897 20349 11931 20383
rect 11931 20349 11940 20383
rect 11888 20340 11940 20349
rect 12164 20340 12216 20392
rect 15200 20408 15252 20460
rect 16396 20408 16448 20460
rect 12532 20383 12584 20392
rect 12532 20349 12541 20383
rect 12541 20349 12575 20383
rect 12575 20349 12584 20383
rect 12532 20340 12584 20349
rect 12624 20383 12676 20392
rect 12624 20349 12633 20383
rect 12633 20349 12667 20383
rect 12667 20349 12676 20383
rect 15108 20383 15160 20392
rect 12624 20340 12676 20349
rect 15108 20349 15117 20383
rect 15117 20349 15151 20383
rect 15151 20349 15160 20383
rect 15108 20340 15160 20349
rect 10508 20272 10560 20324
rect 19708 20272 19760 20324
rect 20904 20340 20956 20392
rect 21364 20272 21416 20324
rect 4160 20204 4212 20256
rect 5172 20204 5224 20256
rect 5356 20247 5408 20256
rect 5356 20213 5365 20247
rect 5365 20213 5399 20247
rect 5399 20213 5408 20247
rect 5356 20204 5408 20213
rect 5448 20204 5500 20256
rect 15108 20204 15160 20256
rect 7882 20102 7934 20154
rect 7946 20102 7998 20154
rect 8010 20102 8062 20154
rect 8074 20102 8126 20154
rect 14782 20102 14834 20154
rect 14846 20102 14898 20154
rect 14910 20102 14962 20154
rect 14974 20102 15026 20154
rect 3516 20043 3568 20052
rect 3516 20009 3525 20043
rect 3525 20009 3559 20043
rect 3559 20009 3568 20043
rect 3516 20000 3568 20009
rect 4160 20000 4212 20052
rect 5172 20000 5224 20052
rect 3700 19907 3752 19916
rect 3700 19873 3709 19907
rect 3709 19873 3743 19907
rect 3743 19873 3752 19907
rect 3700 19864 3752 19873
rect 4896 19728 4948 19780
rect 4988 19728 5040 19780
rect 5172 19907 5224 19916
rect 5172 19873 5207 19907
rect 5207 19873 5224 19907
rect 5448 19907 5500 19916
rect 5172 19864 5224 19873
rect 5448 19873 5457 19907
rect 5457 19873 5491 19907
rect 5491 19873 5500 19907
rect 5448 19864 5500 19873
rect 5540 19864 5592 19916
rect 7472 20000 7524 20052
rect 7380 19932 7432 19984
rect 10508 20043 10560 20052
rect 10508 20009 10517 20043
rect 10517 20009 10551 20043
rect 10551 20009 10560 20043
rect 10508 20000 10560 20009
rect 15752 20000 15804 20052
rect 21364 20043 21416 20052
rect 21364 20009 21373 20043
rect 21373 20009 21407 20043
rect 21407 20009 21416 20043
rect 21364 20000 21416 20009
rect 15384 19975 15436 19984
rect 15384 19941 15393 19975
rect 15393 19941 15427 19975
rect 15427 19941 15436 19975
rect 15384 19932 15436 19941
rect 7748 19864 7800 19916
rect 8208 19907 8260 19916
rect 8208 19873 8217 19907
rect 8217 19873 8251 19907
rect 8251 19873 8260 19907
rect 8208 19864 8260 19873
rect 10324 19907 10376 19916
rect 10324 19873 10333 19907
rect 10333 19873 10367 19907
rect 10367 19873 10376 19907
rect 10324 19864 10376 19873
rect 14464 19864 14516 19916
rect 15108 19907 15160 19916
rect 15108 19873 15117 19907
rect 15117 19873 15151 19907
rect 15151 19873 15160 19907
rect 15108 19864 15160 19873
rect 15200 19864 15252 19916
rect 20628 19932 20680 19984
rect 15936 19864 15988 19916
rect 16120 19907 16172 19916
rect 16120 19873 16129 19907
rect 16129 19873 16163 19907
rect 16163 19873 16172 19907
rect 16120 19864 16172 19873
rect 16396 19907 16448 19916
rect 14556 19839 14608 19848
rect 5264 19728 5316 19780
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 8852 19728 8904 19780
rect 14924 19796 14976 19848
rect 16396 19873 16405 19907
rect 16405 19873 16439 19907
rect 16439 19873 16448 19907
rect 16396 19864 16448 19873
rect 17776 19864 17828 19916
rect 5724 19660 5776 19712
rect 14648 19660 14700 19712
rect 15200 19660 15252 19712
rect 15752 19660 15804 19712
rect 20904 19796 20956 19848
rect 16488 19728 16540 19780
rect 4432 19558 4484 19610
rect 4496 19558 4548 19610
rect 4560 19558 4612 19610
rect 4624 19558 4676 19610
rect 11332 19558 11384 19610
rect 11396 19558 11448 19610
rect 11460 19558 11512 19610
rect 11524 19558 11576 19610
rect 18232 19558 18284 19610
rect 18296 19558 18348 19610
rect 18360 19558 18412 19610
rect 18424 19558 18476 19610
rect 5448 19456 5500 19508
rect 4896 19388 4948 19440
rect 5356 19388 5408 19440
rect 7748 19456 7800 19508
rect 14556 19456 14608 19508
rect 15016 19456 15068 19508
rect 20628 19499 20680 19508
rect 20628 19465 20637 19499
rect 20637 19465 20671 19499
rect 20671 19465 20680 19499
rect 20628 19456 20680 19465
rect 6460 19388 6512 19440
rect 5172 19252 5224 19304
rect 5632 19252 5684 19304
rect 5724 19295 5776 19304
rect 5724 19261 5733 19295
rect 5733 19261 5767 19295
rect 5767 19261 5776 19295
rect 5724 19252 5776 19261
rect 6460 19252 6512 19304
rect 7472 19320 7524 19372
rect 8760 19320 8812 19372
rect 14648 19363 14700 19372
rect 7564 19295 7616 19304
rect 7564 19261 7573 19295
rect 7573 19261 7607 19295
rect 7607 19261 7616 19295
rect 7564 19252 7616 19261
rect 8300 19295 8352 19304
rect 7656 19227 7708 19236
rect 7656 19193 7665 19227
rect 7665 19193 7699 19227
rect 7699 19193 7708 19227
rect 7656 19184 7708 19193
rect 5816 19159 5868 19168
rect 5816 19125 5825 19159
rect 5825 19125 5859 19159
rect 5859 19125 5868 19159
rect 5816 19116 5868 19125
rect 7564 19116 7616 19168
rect 8300 19261 8309 19295
rect 8309 19261 8343 19295
rect 8343 19261 8352 19295
rect 8300 19252 8352 19261
rect 9588 19252 9640 19304
rect 12716 19295 12768 19304
rect 12716 19261 12725 19295
rect 12725 19261 12759 19295
rect 12759 19261 12768 19295
rect 12716 19252 12768 19261
rect 13912 19252 13964 19304
rect 14648 19329 14657 19363
rect 14657 19329 14691 19363
rect 14691 19329 14700 19363
rect 14648 19320 14700 19329
rect 14464 19252 14516 19304
rect 14740 19295 14792 19304
rect 14740 19261 14749 19295
rect 14749 19261 14783 19295
rect 14783 19261 14792 19295
rect 14740 19252 14792 19261
rect 14924 19295 14976 19304
rect 14924 19261 14933 19295
rect 14933 19261 14967 19295
rect 14967 19261 14976 19295
rect 14924 19252 14976 19261
rect 17132 19252 17184 19304
rect 20444 19295 20496 19304
rect 20444 19261 20453 19295
rect 20453 19261 20487 19295
rect 20487 19261 20496 19295
rect 20444 19252 20496 19261
rect 9220 19116 9272 19168
rect 12624 19159 12676 19168
rect 12624 19125 12633 19159
rect 12633 19125 12667 19159
rect 12667 19125 12676 19159
rect 12624 19116 12676 19125
rect 12992 19116 13044 19168
rect 13912 19116 13964 19168
rect 14648 19116 14700 19168
rect 15016 19227 15068 19236
rect 15016 19193 15025 19227
rect 15025 19193 15059 19227
rect 15059 19193 15068 19227
rect 15200 19227 15252 19236
rect 15016 19184 15068 19193
rect 15200 19193 15209 19227
rect 15209 19193 15243 19227
rect 15243 19193 15252 19227
rect 15200 19184 15252 19193
rect 15752 19116 15804 19168
rect 17684 19116 17736 19168
rect 7882 19014 7934 19066
rect 7946 19014 7998 19066
rect 8010 19014 8062 19066
rect 8074 19014 8126 19066
rect 14782 19014 14834 19066
rect 14846 19014 14898 19066
rect 14910 19014 14962 19066
rect 14974 19014 15026 19066
rect 12992 18887 13044 18896
rect 12992 18853 13001 18887
rect 13001 18853 13035 18887
rect 13035 18853 13044 18887
rect 12992 18844 13044 18853
rect 6460 18776 6512 18828
rect 8484 18708 8536 18760
rect 8852 18776 8904 18828
rect 9220 18819 9272 18828
rect 9220 18785 9230 18819
rect 9230 18785 9264 18819
rect 9264 18785 9272 18819
rect 9220 18776 9272 18785
rect 9588 18819 9640 18828
rect 9588 18785 9602 18819
rect 9602 18785 9636 18819
rect 9636 18785 9640 18819
rect 9588 18776 9640 18785
rect 12532 18819 12584 18828
rect 12532 18785 12541 18819
rect 12541 18785 12575 18819
rect 12575 18785 12584 18819
rect 12532 18776 12584 18785
rect 12716 18776 12768 18828
rect 17684 18844 17736 18896
rect 13360 18819 13412 18828
rect 13360 18785 13369 18819
rect 13369 18785 13403 18819
rect 13403 18785 13412 18819
rect 15844 18819 15896 18828
rect 13360 18776 13412 18785
rect 15844 18785 15853 18819
rect 15853 18785 15887 18819
rect 15887 18785 15896 18819
rect 15844 18776 15896 18785
rect 16028 18819 16080 18828
rect 16028 18785 16037 18819
rect 16037 18785 16071 18819
rect 16071 18785 16080 18819
rect 16028 18776 16080 18785
rect 16120 18819 16172 18828
rect 16120 18785 16129 18819
rect 16129 18785 16163 18819
rect 16163 18785 16172 18819
rect 16120 18776 16172 18785
rect 16488 18776 16540 18828
rect 19156 18819 19208 18828
rect 19156 18785 19165 18819
rect 19165 18785 19199 18819
rect 19199 18785 19208 18819
rect 19156 18776 19208 18785
rect 12808 18751 12860 18760
rect 12808 18717 12817 18751
rect 12817 18717 12851 18751
rect 12851 18717 12860 18751
rect 12808 18708 12860 18717
rect 16212 18751 16264 18760
rect 16212 18717 16221 18751
rect 16221 18717 16255 18751
rect 16255 18717 16264 18751
rect 16212 18708 16264 18717
rect 17684 18708 17736 18760
rect 18420 18751 18472 18760
rect 18420 18717 18429 18751
rect 18429 18717 18463 18751
rect 18463 18717 18472 18751
rect 18420 18708 18472 18717
rect 18788 18751 18840 18760
rect 18788 18717 18797 18751
rect 18797 18717 18831 18751
rect 18831 18717 18840 18751
rect 18788 18708 18840 18717
rect 19064 18708 19116 18760
rect 19340 18776 19392 18828
rect 19616 18819 19668 18828
rect 19616 18785 19625 18819
rect 19625 18785 19659 18819
rect 19659 18785 19668 18819
rect 19616 18776 19668 18785
rect 19432 18708 19484 18760
rect 8852 18640 8904 18692
rect 5632 18572 5684 18624
rect 7564 18572 7616 18624
rect 8944 18572 8996 18624
rect 9404 18572 9456 18624
rect 13176 18615 13228 18624
rect 13176 18581 13185 18615
rect 13185 18581 13219 18615
rect 13219 18581 13228 18615
rect 13176 18572 13228 18581
rect 16488 18572 16540 18624
rect 19800 18572 19852 18624
rect 4432 18470 4484 18522
rect 4496 18470 4548 18522
rect 4560 18470 4612 18522
rect 4624 18470 4676 18522
rect 11332 18470 11384 18522
rect 11396 18470 11448 18522
rect 11460 18470 11512 18522
rect 11524 18470 11576 18522
rect 18232 18470 18284 18522
rect 18296 18470 18348 18522
rect 18360 18470 18412 18522
rect 18424 18470 18476 18522
rect 8484 18411 8536 18420
rect 8484 18377 8493 18411
rect 8493 18377 8527 18411
rect 8527 18377 8536 18411
rect 8484 18368 8536 18377
rect 8944 18411 8996 18420
rect 8944 18377 8953 18411
rect 8953 18377 8987 18411
rect 8987 18377 8996 18411
rect 8944 18368 8996 18377
rect 16120 18368 16172 18420
rect 12992 18300 13044 18352
rect 13360 18300 13412 18352
rect 19156 18300 19208 18352
rect 2504 18232 2556 18284
rect 4620 18232 4672 18284
rect 9404 18275 9456 18284
rect 9404 18241 9413 18275
rect 9413 18241 9447 18275
rect 9447 18241 9456 18275
rect 9404 18232 9456 18241
rect 9128 18207 9180 18216
rect 3976 18096 4028 18148
rect 9128 18173 9137 18207
rect 9137 18173 9171 18207
rect 9171 18173 9180 18207
rect 9128 18164 9180 18173
rect 9312 18164 9364 18216
rect 10324 18207 10376 18216
rect 10324 18173 10333 18207
rect 10333 18173 10367 18207
rect 10367 18173 10376 18207
rect 10324 18164 10376 18173
rect 10968 18164 11020 18216
rect 12624 18207 12676 18216
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 12624 18164 12676 18173
rect 13176 18232 13228 18284
rect 12992 18207 13044 18216
rect 12992 18173 13001 18207
rect 13001 18173 13035 18207
rect 13035 18173 13044 18207
rect 12992 18164 13044 18173
rect 13268 18207 13320 18216
rect 13268 18173 13277 18207
rect 13277 18173 13311 18207
rect 13311 18173 13320 18207
rect 13268 18164 13320 18173
rect 19064 18232 19116 18284
rect 16580 18207 16632 18216
rect 16580 18173 16589 18207
rect 16589 18173 16623 18207
rect 16623 18173 16632 18207
rect 16580 18164 16632 18173
rect 5172 18028 5224 18080
rect 16212 18096 16264 18148
rect 16856 18096 16908 18148
rect 19340 18164 19392 18216
rect 19432 18207 19484 18216
rect 19432 18173 19441 18207
rect 19441 18173 19475 18207
rect 19475 18173 19484 18207
rect 21272 18232 21324 18284
rect 19432 18164 19484 18173
rect 19800 18207 19852 18216
rect 19800 18173 19809 18207
rect 19809 18173 19843 18207
rect 19843 18173 19852 18207
rect 19800 18164 19852 18173
rect 8668 18028 8720 18080
rect 8760 18028 8812 18080
rect 9588 18028 9640 18080
rect 10600 18028 10652 18080
rect 16488 18028 16540 18080
rect 18788 18028 18840 18080
rect 7882 17926 7934 17978
rect 7946 17926 7998 17978
rect 8010 17926 8062 17978
rect 8074 17926 8126 17978
rect 14782 17926 14834 17978
rect 14846 17926 14898 17978
rect 14910 17926 14962 17978
rect 14974 17926 15026 17978
rect 3976 17824 4028 17876
rect 4620 17867 4672 17876
rect 4620 17833 4629 17867
rect 4629 17833 4663 17867
rect 4663 17833 4672 17867
rect 4620 17824 4672 17833
rect 6000 17867 6052 17876
rect 6000 17833 6009 17867
rect 6009 17833 6043 17867
rect 6043 17833 6052 17867
rect 6000 17824 6052 17833
rect 4988 17799 5040 17808
rect 4988 17765 4997 17799
rect 4997 17765 5031 17799
rect 5031 17765 5040 17799
rect 4988 17756 5040 17765
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 3700 17688 3752 17740
rect 1584 17527 1636 17536
rect 1584 17493 1593 17527
rect 1593 17493 1627 17527
rect 1627 17493 1636 17527
rect 1584 17484 1636 17493
rect 5172 17688 5224 17740
rect 5264 17731 5316 17740
rect 5264 17697 5273 17731
rect 5273 17697 5307 17731
rect 5307 17697 5316 17731
rect 5816 17756 5868 17808
rect 9588 17799 9640 17808
rect 5724 17731 5776 17740
rect 5264 17688 5316 17697
rect 5724 17697 5733 17731
rect 5733 17697 5767 17731
rect 5767 17697 5776 17731
rect 5724 17688 5776 17697
rect 6276 17688 6328 17740
rect 9588 17765 9597 17799
rect 9597 17765 9631 17799
rect 9631 17765 9640 17799
rect 9588 17756 9640 17765
rect 10600 17756 10652 17808
rect 7748 17688 7800 17740
rect 8760 17688 8812 17740
rect 9036 17688 9088 17740
rect 11796 17688 11848 17740
rect 12348 17688 12400 17740
rect 12440 17688 12492 17740
rect 13912 17688 13964 17740
rect 15844 17824 15896 17876
rect 17316 17824 17368 17876
rect 16212 17756 16264 17808
rect 6736 17620 6788 17672
rect 8208 17663 8260 17672
rect 8208 17629 8217 17663
rect 8217 17629 8251 17663
rect 8251 17629 8260 17663
rect 8208 17620 8260 17629
rect 8300 17663 8352 17672
rect 8300 17629 8309 17663
rect 8309 17629 8343 17663
rect 8343 17629 8352 17663
rect 15200 17688 15252 17740
rect 16396 17688 16448 17740
rect 20444 17688 20496 17740
rect 21456 17731 21508 17740
rect 21456 17697 21465 17731
rect 21465 17697 21499 17731
rect 21499 17697 21508 17731
rect 21456 17688 21508 17697
rect 8300 17620 8352 17629
rect 16580 17620 16632 17672
rect 6644 17552 6696 17604
rect 8484 17552 8536 17604
rect 12716 17552 12768 17604
rect 8392 17484 8444 17536
rect 8668 17484 8720 17536
rect 10140 17484 10192 17536
rect 12624 17527 12676 17536
rect 12624 17493 12633 17527
rect 12633 17493 12667 17527
rect 12667 17493 12676 17527
rect 12624 17484 12676 17493
rect 14740 17484 14792 17536
rect 20996 17484 21048 17536
rect 21180 17484 21232 17536
rect 4432 17382 4484 17434
rect 4496 17382 4548 17434
rect 4560 17382 4612 17434
rect 4624 17382 4676 17434
rect 11332 17382 11384 17434
rect 11396 17382 11448 17434
rect 11460 17382 11512 17434
rect 11524 17382 11576 17434
rect 18232 17382 18284 17434
rect 18296 17382 18348 17434
rect 18360 17382 18412 17434
rect 18424 17382 18476 17434
rect 8208 17280 8260 17332
rect 9128 17280 9180 17332
rect 9496 17280 9548 17332
rect 12624 17280 12676 17332
rect 13268 17280 13320 17332
rect 16212 17323 16264 17332
rect 5908 17212 5960 17264
rect 5172 17076 5224 17128
rect 5632 17119 5684 17128
rect 5632 17085 5641 17119
rect 5641 17085 5675 17119
rect 5675 17085 5684 17119
rect 5632 17076 5684 17085
rect 5816 17076 5868 17128
rect 6460 17119 6512 17128
rect 5724 17008 5776 17060
rect 6460 17085 6469 17119
rect 6469 17085 6503 17119
rect 6503 17085 6512 17119
rect 6460 17076 6512 17085
rect 7380 17212 7432 17264
rect 12808 17212 12860 17264
rect 6736 17187 6788 17196
rect 6736 17153 6745 17187
rect 6745 17153 6779 17187
rect 6779 17153 6788 17187
rect 6736 17144 6788 17153
rect 12440 17187 12492 17196
rect 12440 17153 12449 17187
rect 12449 17153 12483 17187
rect 12483 17153 12492 17187
rect 12624 17187 12676 17196
rect 12440 17144 12492 17153
rect 12624 17153 12633 17187
rect 12633 17153 12667 17187
rect 12667 17153 12676 17187
rect 12624 17144 12676 17153
rect 16212 17289 16221 17323
rect 16221 17289 16255 17323
rect 16255 17289 16264 17323
rect 16212 17280 16264 17289
rect 14740 17187 14792 17196
rect 14740 17153 14749 17187
rect 14749 17153 14783 17187
rect 14783 17153 14792 17187
rect 14740 17144 14792 17153
rect 17684 17144 17736 17196
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 10140 17119 10192 17128
rect 6276 17008 6328 17060
rect 10140 17085 10149 17119
rect 10149 17085 10183 17119
rect 10183 17085 10192 17119
rect 10140 17076 10192 17085
rect 12164 17076 12216 17128
rect 12348 17119 12400 17128
rect 12348 17085 12357 17119
rect 12357 17085 12391 17119
rect 12391 17085 12400 17119
rect 12348 17076 12400 17085
rect 12716 17119 12768 17128
rect 12716 17085 12725 17119
rect 12725 17085 12759 17119
rect 12759 17085 12768 17119
rect 12716 17076 12768 17085
rect 17132 17008 17184 17060
rect 17592 17008 17644 17060
rect 19984 17051 20036 17060
rect 19984 17017 19993 17051
rect 19993 17017 20027 17051
rect 20027 17017 20036 17051
rect 19984 17008 20036 17017
rect 20996 17008 21048 17060
rect 17316 16940 17368 16992
rect 19708 16940 19760 16992
rect 7882 16838 7934 16890
rect 7946 16838 7998 16890
rect 8010 16838 8062 16890
rect 8074 16838 8126 16890
rect 14782 16838 14834 16890
rect 14846 16838 14898 16890
rect 14910 16838 14962 16890
rect 14974 16838 15026 16890
rect 16580 16736 16632 16788
rect 16948 16736 17000 16788
rect 5816 16643 5868 16652
rect 5816 16609 5825 16643
rect 5825 16609 5859 16643
rect 5859 16609 5868 16643
rect 5816 16600 5868 16609
rect 6000 16600 6052 16652
rect 6920 16600 6972 16652
rect 8392 16668 8444 16720
rect 16856 16668 16908 16720
rect 17132 16711 17184 16720
rect 17132 16677 17141 16711
rect 17141 16677 17175 16711
rect 17175 16677 17184 16711
rect 17132 16668 17184 16677
rect 17960 16736 18012 16788
rect 19984 16736 20036 16788
rect 8852 16600 8904 16652
rect 15016 16600 15068 16652
rect 15200 16600 15252 16652
rect 16028 16600 16080 16652
rect 17040 16643 17092 16652
rect 17040 16609 17049 16643
rect 17049 16609 17083 16643
rect 17083 16609 17092 16643
rect 17040 16600 17092 16609
rect 18604 16668 18656 16720
rect 18696 16668 18748 16720
rect 17592 16643 17644 16652
rect 17592 16609 17601 16643
rect 17601 16609 17635 16643
rect 17635 16609 17644 16643
rect 19616 16643 19668 16652
rect 17592 16600 17644 16609
rect 19616 16609 19625 16643
rect 19625 16609 19659 16643
rect 19659 16609 19668 16643
rect 19616 16600 19668 16609
rect 19708 16600 19760 16652
rect 5908 16507 5960 16516
rect 5908 16473 5917 16507
rect 5917 16473 5951 16507
rect 5951 16473 5960 16507
rect 5908 16464 5960 16473
rect 6552 16396 6604 16448
rect 17224 16396 17276 16448
rect 19524 16396 19576 16448
rect 19892 16396 19944 16448
rect 4432 16294 4484 16346
rect 4496 16294 4548 16346
rect 4560 16294 4612 16346
rect 4624 16294 4676 16346
rect 11332 16294 11384 16346
rect 11396 16294 11448 16346
rect 11460 16294 11512 16346
rect 11524 16294 11576 16346
rect 18232 16294 18284 16346
rect 18296 16294 18348 16346
rect 18360 16294 18412 16346
rect 18424 16294 18476 16346
rect 1952 15988 2004 16040
rect 2872 15988 2924 16040
rect 5264 15988 5316 16040
rect 15108 16192 15160 16244
rect 6644 16124 6696 16176
rect 9312 16124 9364 16176
rect 14556 16124 14608 16176
rect 6552 16031 6604 16040
rect 6552 15997 6562 16031
rect 6562 15997 6596 16031
rect 6596 15997 6604 16031
rect 6828 16056 6880 16108
rect 6552 15988 6604 15997
rect 6920 16031 6972 16040
rect 6920 15997 6934 16031
rect 6934 15997 6968 16031
rect 6968 15997 6972 16031
rect 6920 15988 6972 15997
rect 8852 16031 8904 16040
rect 2688 15920 2740 15972
rect 8852 15997 8861 16031
rect 8861 15997 8895 16031
rect 8895 15997 8904 16031
rect 8852 15988 8904 15997
rect 8944 16031 8996 16040
rect 8944 15997 8958 16031
rect 8958 15997 8992 16031
rect 8992 15997 8996 16031
rect 10968 16031 11020 16040
rect 8944 15988 8996 15997
rect 10968 15997 10977 16031
rect 10977 15997 11011 16031
rect 11011 15997 11020 16031
rect 10968 15988 11020 15997
rect 6920 15852 6972 15904
rect 8392 15852 8444 15904
rect 9128 15895 9180 15904
rect 9128 15861 9137 15895
rect 9137 15861 9171 15895
rect 9171 15861 9180 15895
rect 9128 15852 9180 15861
rect 11244 15852 11296 15904
rect 16212 16056 16264 16108
rect 17592 16192 17644 16244
rect 18696 16235 18748 16244
rect 18696 16201 18705 16235
rect 18705 16201 18739 16235
rect 18739 16201 18748 16235
rect 18696 16192 18748 16201
rect 19064 16235 19116 16244
rect 19064 16201 19073 16235
rect 19073 16201 19107 16235
rect 19107 16201 19116 16235
rect 19064 16192 19116 16201
rect 17224 16099 17276 16108
rect 17224 16065 17233 16099
rect 17233 16065 17267 16099
rect 17267 16065 17276 16099
rect 17224 16056 17276 16065
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 16856 15988 16908 16040
rect 19524 16031 19576 16040
rect 19524 15997 19533 16031
rect 19533 15997 19567 16031
rect 19567 15997 19576 16031
rect 19524 15988 19576 15997
rect 19892 16031 19944 16040
rect 17960 15920 18012 15972
rect 18604 15920 18656 15972
rect 18972 15920 19024 15972
rect 19892 15997 19901 16031
rect 19901 15997 19935 16031
rect 19935 15997 19944 16031
rect 19892 15988 19944 15997
rect 19984 15963 20036 15972
rect 19984 15929 19993 15963
rect 19993 15929 20027 15963
rect 20027 15929 20036 15963
rect 19984 15920 20036 15929
rect 7882 15750 7934 15802
rect 7946 15750 7998 15802
rect 8010 15750 8062 15802
rect 8074 15750 8126 15802
rect 14782 15750 14834 15802
rect 14846 15750 14898 15802
rect 14910 15750 14962 15802
rect 14974 15750 15026 15802
rect 8944 15648 8996 15700
rect 9036 15648 9088 15700
rect 12164 15691 12216 15700
rect 12164 15657 12173 15691
rect 12173 15657 12207 15691
rect 12207 15657 12216 15691
rect 12164 15648 12216 15657
rect 12992 15648 13044 15700
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 3240 15555 3292 15564
rect 3240 15521 3249 15555
rect 3249 15521 3283 15555
rect 3283 15521 3292 15555
rect 3240 15512 3292 15521
rect 1952 15444 2004 15496
rect 2688 15376 2740 15428
rect 8484 15512 8536 15564
rect 8760 15580 8812 15632
rect 11244 15580 11296 15632
rect 17132 15691 17184 15700
rect 9588 15512 9640 15564
rect 14556 15555 14608 15564
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 9312 15487 9364 15496
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 12532 15444 12584 15496
rect 14556 15521 14562 15555
rect 14562 15521 14596 15555
rect 14596 15521 14608 15555
rect 14556 15512 14608 15521
rect 17132 15657 17141 15691
rect 17141 15657 17175 15691
rect 17175 15657 17184 15691
rect 17132 15648 17184 15657
rect 17316 15691 17368 15700
rect 17316 15657 17325 15691
rect 17325 15657 17359 15691
rect 17359 15657 17368 15691
rect 17316 15648 17368 15657
rect 17684 15648 17736 15700
rect 19432 15648 19484 15700
rect 16948 15623 17000 15632
rect 16948 15589 16957 15623
rect 16957 15589 16991 15623
rect 16991 15589 17000 15623
rect 16948 15580 17000 15589
rect 17040 15580 17092 15632
rect 15200 15512 15252 15564
rect 20168 15648 20220 15700
rect 21272 15691 21324 15700
rect 21272 15657 21281 15691
rect 21281 15657 21315 15691
rect 21315 15657 21324 15691
rect 21272 15648 21324 15657
rect 21456 15555 21508 15564
rect 19984 15444 20036 15496
rect 21456 15521 21465 15555
rect 21465 15521 21499 15555
rect 21499 15521 21508 15555
rect 21456 15512 21508 15521
rect 9864 15376 9916 15428
rect 1860 15308 1912 15360
rect 5632 15308 5684 15360
rect 7288 15308 7340 15360
rect 10876 15308 10928 15360
rect 18604 15308 18656 15360
rect 4432 15206 4484 15258
rect 4496 15206 4548 15258
rect 4560 15206 4612 15258
rect 4624 15206 4676 15258
rect 11332 15206 11384 15258
rect 11396 15206 11448 15258
rect 11460 15206 11512 15258
rect 11524 15206 11576 15258
rect 18232 15206 18284 15258
rect 18296 15206 18348 15258
rect 18360 15206 18412 15258
rect 18424 15206 18476 15258
rect 1952 15104 2004 15156
rect 6644 15147 6696 15156
rect 6644 15113 6653 15147
rect 6653 15113 6687 15147
rect 6687 15113 6696 15147
rect 6644 15104 6696 15113
rect 6828 15147 6880 15156
rect 6828 15113 6837 15147
rect 6837 15113 6871 15147
rect 6871 15113 6880 15147
rect 6828 15104 6880 15113
rect 7288 15147 7340 15156
rect 7288 15113 7297 15147
rect 7297 15113 7331 15147
rect 7331 15113 7340 15147
rect 7288 15104 7340 15113
rect 12440 15104 12492 15156
rect 2044 15011 2096 15020
rect 2044 14977 2053 15011
rect 2053 14977 2087 15011
rect 2087 14977 2096 15011
rect 2044 14968 2096 14977
rect 1768 14900 1820 14952
rect 2872 14943 2924 14952
rect 2872 14909 2881 14943
rect 2881 14909 2915 14943
rect 2915 14909 2924 14943
rect 9588 15036 9640 15088
rect 6920 14968 6972 15020
rect 2872 14900 2924 14909
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 3332 14832 3384 14884
rect 5264 14900 5316 14952
rect 7012 14943 7064 14952
rect 7012 14909 7021 14943
rect 7021 14909 7055 14943
rect 7055 14909 7064 14943
rect 7012 14900 7064 14909
rect 8484 14968 8536 15020
rect 12072 14968 12124 15020
rect 7564 14900 7616 14952
rect 9864 14900 9916 14952
rect 9772 14875 9824 14884
rect 9772 14841 9781 14875
rect 9781 14841 9815 14875
rect 9815 14841 9824 14875
rect 9772 14832 9824 14841
rect 3240 14764 3292 14816
rect 4896 14807 4948 14816
rect 4896 14773 4905 14807
rect 4905 14773 4939 14807
rect 4939 14773 4948 14807
rect 4896 14764 4948 14773
rect 5632 14764 5684 14816
rect 11152 14832 11204 14884
rect 14648 14900 14700 14952
rect 15200 14832 15252 14884
rect 19984 14943 20036 14952
rect 15568 14764 15620 14816
rect 15752 14764 15804 14816
rect 19984 14909 19993 14943
rect 19993 14909 20027 14943
rect 20027 14909 20036 14943
rect 19984 14900 20036 14909
rect 20168 14943 20220 14952
rect 20168 14909 20177 14943
rect 20177 14909 20211 14943
rect 20211 14909 20220 14943
rect 20168 14900 20220 14909
rect 19892 14875 19944 14884
rect 19892 14841 19901 14875
rect 19901 14841 19935 14875
rect 19935 14841 19944 14875
rect 19892 14832 19944 14841
rect 20352 14764 20404 14816
rect 7882 14662 7934 14714
rect 7946 14662 7998 14714
rect 8010 14662 8062 14714
rect 8074 14662 8126 14714
rect 14782 14662 14834 14714
rect 14846 14662 14898 14714
rect 14910 14662 14962 14714
rect 14974 14662 15026 14714
rect 5264 14560 5316 14612
rect 7288 14560 7340 14612
rect 10968 14560 11020 14612
rect 14556 14603 14608 14612
rect 14556 14569 14565 14603
rect 14565 14569 14599 14603
rect 14599 14569 14608 14603
rect 14556 14560 14608 14569
rect 14648 14560 14700 14612
rect 4896 14492 4948 14544
rect 5632 14535 5684 14544
rect 5632 14501 5641 14535
rect 5641 14501 5675 14535
rect 5675 14501 5684 14535
rect 5632 14492 5684 14501
rect 17132 14560 17184 14612
rect 18972 14603 19024 14612
rect 18972 14569 18981 14603
rect 18981 14569 19015 14603
rect 19015 14569 19024 14603
rect 18972 14560 19024 14569
rect 20168 14603 20220 14612
rect 20168 14569 20177 14603
rect 20177 14569 20211 14603
rect 20211 14569 20220 14603
rect 20168 14560 20220 14569
rect 20352 14603 20404 14612
rect 20352 14569 20361 14603
rect 20361 14569 20395 14603
rect 20395 14569 20404 14603
rect 20352 14560 20404 14569
rect 8484 14424 8536 14476
rect 9036 14424 9088 14476
rect 13912 14424 13964 14476
rect 13820 14356 13872 14408
rect 5264 14220 5316 14272
rect 6828 14220 6880 14272
rect 7748 14220 7800 14272
rect 8668 14220 8720 14272
rect 15200 14467 15252 14476
rect 15200 14433 15209 14467
rect 15209 14433 15243 14467
rect 15243 14433 15252 14467
rect 15200 14424 15252 14433
rect 15568 14424 15620 14476
rect 15752 14467 15804 14476
rect 15752 14433 15761 14467
rect 15761 14433 15795 14467
rect 15795 14433 15804 14467
rect 15752 14424 15804 14433
rect 18052 14424 18104 14476
rect 18696 14424 18748 14476
rect 19156 14424 19208 14476
rect 19340 14424 19392 14476
rect 19892 14424 19944 14476
rect 15568 14220 15620 14272
rect 20076 14220 20128 14272
rect 20352 14220 20404 14272
rect 4432 14118 4484 14170
rect 4496 14118 4548 14170
rect 4560 14118 4612 14170
rect 4624 14118 4676 14170
rect 11332 14118 11384 14170
rect 11396 14118 11448 14170
rect 11460 14118 11512 14170
rect 11524 14118 11576 14170
rect 18232 14118 18284 14170
rect 18296 14118 18348 14170
rect 18360 14118 18412 14170
rect 18424 14118 18476 14170
rect 1952 14016 2004 14068
rect 7472 14016 7524 14068
rect 8024 14016 8076 14068
rect 8576 14016 8628 14068
rect 9772 14016 9824 14068
rect 13820 14016 13872 14068
rect 15108 14016 15160 14068
rect 18972 14016 19024 14068
rect 5816 13948 5868 14000
rect 5172 13812 5224 13864
rect 6460 13812 6512 13864
rect 6644 13855 6696 13864
rect 6644 13821 6653 13855
rect 6653 13821 6687 13855
rect 6687 13821 6696 13855
rect 6644 13812 6696 13821
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 18052 13948 18104 14000
rect 6736 13676 6788 13728
rect 7564 13812 7616 13864
rect 9588 13880 9640 13932
rect 7196 13744 7248 13796
rect 8024 13855 8076 13864
rect 8024 13821 8033 13855
rect 8033 13821 8067 13855
rect 8067 13821 8076 13855
rect 9496 13855 9548 13864
rect 8024 13812 8076 13821
rect 9496 13821 9505 13855
rect 9505 13821 9539 13855
rect 9539 13821 9548 13855
rect 9496 13812 9548 13821
rect 7656 13719 7708 13728
rect 7656 13685 7665 13719
rect 7665 13685 7699 13719
rect 7699 13685 7708 13719
rect 7656 13676 7708 13685
rect 8208 13676 8260 13728
rect 10140 13812 10192 13864
rect 17868 13855 17920 13864
rect 17868 13821 17877 13855
rect 17877 13821 17911 13855
rect 17911 13821 17920 13855
rect 17868 13812 17920 13821
rect 19340 13812 19392 13864
rect 18696 13744 18748 13796
rect 9864 13676 9916 13728
rect 17960 13719 18012 13728
rect 17960 13685 17969 13719
rect 17969 13685 18003 13719
rect 18003 13685 18012 13719
rect 17960 13676 18012 13685
rect 7882 13574 7934 13626
rect 7946 13574 7998 13626
rect 8010 13574 8062 13626
rect 8074 13574 8126 13626
rect 14782 13574 14834 13626
rect 14846 13574 14898 13626
rect 14910 13574 14962 13626
rect 14974 13574 15026 13626
rect 1584 13472 1636 13524
rect 3332 13515 3384 13524
rect 3332 13481 3341 13515
rect 3341 13481 3375 13515
rect 3375 13481 3384 13515
rect 3332 13472 3384 13481
rect 7380 13515 7432 13524
rect 7380 13481 7389 13515
rect 7389 13481 7423 13515
rect 7423 13481 7432 13515
rect 7380 13472 7432 13481
rect 8300 13515 8352 13524
rect 8300 13481 8309 13515
rect 8309 13481 8343 13515
rect 8343 13481 8352 13515
rect 8300 13472 8352 13481
rect 5540 13404 5592 13456
rect 12072 13447 12124 13456
rect 12072 13413 12081 13447
rect 12081 13413 12115 13447
rect 12115 13413 12124 13447
rect 12072 13404 12124 13413
rect 1768 13311 1820 13320
rect 1768 13277 1777 13311
rect 1777 13277 1811 13311
rect 1811 13277 1820 13311
rect 1768 13268 1820 13277
rect 3148 13336 3200 13388
rect 6644 13336 6696 13388
rect 4896 13268 4948 13320
rect 8116 13336 8168 13388
rect 10968 13336 11020 13388
rect 14372 13404 14424 13456
rect 14648 13447 14700 13456
rect 14648 13413 14657 13447
rect 14657 13413 14691 13447
rect 14691 13413 14700 13447
rect 14648 13404 14700 13413
rect 12808 13379 12860 13388
rect 10048 13268 10100 13320
rect 12808 13345 12817 13379
rect 12817 13345 12851 13379
rect 12851 13345 12860 13379
rect 12808 13336 12860 13345
rect 4804 13200 4856 13252
rect 12164 13311 12216 13320
rect 12164 13277 12173 13311
rect 12173 13277 12207 13311
rect 12207 13277 12216 13311
rect 13912 13336 13964 13388
rect 15108 13336 15160 13388
rect 12164 13268 12216 13277
rect 10416 13200 10468 13252
rect 10876 13200 10928 13252
rect 12256 13200 12308 13252
rect 15568 13268 15620 13320
rect 16672 13404 16724 13456
rect 17684 13404 17736 13456
rect 18052 13379 18104 13388
rect 18052 13345 18061 13379
rect 18061 13345 18095 13379
rect 18095 13345 18104 13379
rect 18052 13336 18104 13345
rect 18696 13379 18748 13388
rect 18696 13345 18705 13379
rect 18705 13345 18739 13379
rect 18739 13345 18748 13379
rect 18696 13336 18748 13345
rect 18972 13404 19024 13456
rect 19340 13404 19392 13456
rect 20076 13404 20128 13456
rect 19616 13379 19668 13388
rect 13728 13200 13780 13252
rect 2136 13132 2188 13184
rect 13268 13132 13320 13184
rect 15844 13132 15896 13184
rect 17684 13311 17736 13320
rect 17684 13277 17693 13311
rect 17693 13277 17727 13311
rect 17727 13277 17736 13311
rect 17960 13311 18012 13320
rect 17684 13268 17736 13277
rect 17960 13277 17969 13311
rect 17969 13277 18003 13311
rect 18003 13277 18012 13311
rect 17960 13268 18012 13277
rect 18604 13268 18656 13320
rect 19156 13268 19208 13320
rect 19616 13345 19625 13379
rect 19625 13345 19659 13379
rect 19659 13345 19668 13379
rect 19616 13336 19668 13345
rect 19800 13379 19852 13388
rect 19800 13345 19809 13379
rect 19809 13345 19843 13379
rect 19843 13345 19852 13379
rect 19800 13336 19852 13345
rect 20444 13336 20496 13388
rect 21456 13379 21508 13388
rect 21456 13345 21465 13379
rect 21465 13345 21499 13379
rect 21499 13345 21508 13379
rect 21456 13336 21508 13345
rect 17316 13132 17368 13184
rect 18880 13132 18932 13184
rect 19984 13132 20036 13184
rect 20720 13132 20772 13184
rect 4432 13030 4484 13082
rect 4496 13030 4548 13082
rect 4560 13030 4612 13082
rect 4624 13030 4676 13082
rect 11332 13030 11384 13082
rect 11396 13030 11448 13082
rect 11460 13030 11512 13082
rect 11524 13030 11576 13082
rect 18232 13030 18284 13082
rect 18296 13030 18348 13082
rect 18360 13030 18412 13082
rect 18424 13030 18476 13082
rect 1492 12971 1544 12980
rect 1492 12937 1501 12971
rect 1501 12937 1535 12971
rect 1535 12937 1544 12971
rect 1492 12928 1544 12937
rect 3148 12971 3200 12980
rect 3148 12937 3157 12971
rect 3157 12937 3191 12971
rect 3191 12937 3200 12971
rect 3148 12928 3200 12937
rect 4896 12971 4948 12980
rect 4896 12937 4905 12971
rect 4905 12937 4939 12971
rect 4939 12937 4948 12971
rect 4896 12928 4948 12937
rect 5264 12971 5316 12980
rect 5264 12937 5273 12971
rect 5273 12937 5307 12971
rect 5307 12937 5316 12971
rect 5264 12928 5316 12937
rect 6184 12928 6236 12980
rect 6644 12928 6696 12980
rect 8668 12928 8720 12980
rect 9864 12971 9916 12980
rect 9864 12937 9873 12971
rect 9873 12937 9907 12971
rect 9907 12937 9916 12971
rect 9864 12928 9916 12937
rect 10048 12971 10100 12980
rect 10048 12937 10057 12971
rect 10057 12937 10091 12971
rect 10091 12937 10100 12971
rect 10048 12928 10100 12937
rect 12072 12928 12124 12980
rect 2136 12767 2188 12776
rect 2136 12733 2145 12767
rect 2145 12733 2179 12767
rect 2179 12733 2188 12767
rect 2136 12724 2188 12733
rect 2964 12724 3016 12776
rect 3332 12724 3384 12776
rect 5172 12767 5224 12776
rect 5172 12733 5181 12767
rect 5181 12733 5215 12767
rect 5215 12733 5224 12767
rect 5172 12724 5224 12733
rect 5356 12792 5408 12844
rect 8116 12835 8168 12844
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 8116 12792 8168 12801
rect 9588 12860 9640 12912
rect 9496 12792 9548 12844
rect 11244 12860 11296 12912
rect 12808 12860 12860 12912
rect 6460 12767 6512 12776
rect 6460 12733 6469 12767
rect 6469 12733 6503 12767
rect 6503 12733 6512 12767
rect 6460 12724 6512 12733
rect 7748 12767 7800 12776
rect 7748 12733 7757 12767
rect 7757 12733 7791 12767
rect 7791 12733 7800 12767
rect 7748 12724 7800 12733
rect 8300 12767 8352 12776
rect 8300 12733 8309 12767
rect 8309 12733 8343 12767
rect 8343 12733 8352 12767
rect 8300 12724 8352 12733
rect 8484 12767 8536 12776
rect 8484 12733 8493 12767
rect 8493 12733 8527 12767
rect 8527 12733 8536 12767
rect 8484 12724 8536 12733
rect 10140 12767 10192 12776
rect 3240 12656 3292 12708
rect 6184 12656 6236 12708
rect 7196 12656 7248 12708
rect 7472 12656 7524 12708
rect 7656 12656 7708 12708
rect 10140 12733 10149 12767
rect 10149 12733 10183 12767
rect 10183 12733 10192 12767
rect 10140 12724 10192 12733
rect 12256 12835 12308 12844
rect 12256 12801 12265 12835
rect 12265 12801 12299 12835
rect 12299 12801 12308 12835
rect 16672 12928 16724 12980
rect 17868 12928 17920 12980
rect 20076 12928 20128 12980
rect 12256 12792 12308 12801
rect 13268 12767 13320 12776
rect 9496 12656 9548 12708
rect 9128 12588 9180 12640
rect 11060 12699 11112 12708
rect 11060 12665 11069 12699
rect 11069 12665 11103 12699
rect 11103 12665 11112 12699
rect 11244 12699 11296 12708
rect 11060 12656 11112 12665
rect 11244 12665 11253 12699
rect 11253 12665 11287 12699
rect 11287 12665 11296 12699
rect 11244 12656 11296 12665
rect 11336 12588 11388 12640
rect 11704 12631 11756 12640
rect 11704 12597 11713 12631
rect 11713 12597 11747 12631
rect 11747 12597 11756 12631
rect 11704 12588 11756 12597
rect 13268 12733 13277 12767
rect 13277 12733 13311 12767
rect 13311 12733 13320 12767
rect 13268 12724 13320 12733
rect 16764 12860 16816 12912
rect 19340 12860 19392 12912
rect 17684 12792 17736 12844
rect 19156 12792 19208 12844
rect 19984 12835 20036 12844
rect 19984 12801 19993 12835
rect 19993 12801 20027 12835
rect 20027 12801 20036 12835
rect 19984 12792 20036 12801
rect 17316 12767 17368 12776
rect 17316 12733 17325 12767
rect 17325 12733 17359 12767
rect 17359 12733 17368 12767
rect 17316 12724 17368 12733
rect 18880 12767 18932 12776
rect 18880 12733 18889 12767
rect 18889 12733 18923 12767
rect 18923 12733 18932 12767
rect 18880 12724 18932 12733
rect 17960 12656 18012 12708
rect 18604 12656 18656 12708
rect 20720 12656 20772 12708
rect 12900 12631 12952 12640
rect 12900 12597 12909 12631
rect 12909 12597 12943 12631
rect 12943 12597 12952 12631
rect 12900 12588 12952 12597
rect 15108 12588 15160 12640
rect 19248 12631 19300 12640
rect 19248 12597 19257 12631
rect 19257 12597 19291 12631
rect 19291 12597 19300 12631
rect 19248 12588 19300 12597
rect 19340 12588 19392 12640
rect 20352 12588 20404 12640
rect 7882 12486 7934 12538
rect 7946 12486 7998 12538
rect 8010 12486 8062 12538
rect 8074 12486 8126 12538
rect 14782 12486 14834 12538
rect 14846 12486 14898 12538
rect 14910 12486 14962 12538
rect 14974 12486 15026 12538
rect 5172 12384 5224 12436
rect 5540 12427 5592 12436
rect 5540 12393 5549 12427
rect 5549 12393 5583 12427
rect 5583 12393 5592 12427
rect 5540 12384 5592 12393
rect 3332 12359 3384 12368
rect 3332 12325 3341 12359
rect 3341 12325 3375 12359
rect 3375 12325 3384 12359
rect 3332 12316 3384 12325
rect 4804 12316 4856 12368
rect 6736 12384 6788 12436
rect 10324 12384 10376 12436
rect 12164 12384 12216 12436
rect 14372 12427 14424 12436
rect 14372 12393 14381 12427
rect 14381 12393 14415 12427
rect 14415 12393 14424 12427
rect 14372 12384 14424 12393
rect 3516 12291 3568 12300
rect 3516 12257 3525 12291
rect 3525 12257 3559 12291
rect 3559 12257 3568 12291
rect 3516 12248 3568 12257
rect 5172 12248 5224 12300
rect 5816 12248 5868 12300
rect 7472 12316 7524 12368
rect 11336 12316 11388 12368
rect 15108 12316 15160 12368
rect 15844 12359 15896 12368
rect 15844 12325 15853 12359
rect 15853 12325 15887 12359
rect 15887 12325 15896 12359
rect 15844 12316 15896 12325
rect 6644 12248 6696 12300
rect 11704 12291 11756 12300
rect 11704 12257 11713 12291
rect 11713 12257 11747 12291
rect 11747 12257 11756 12291
rect 11704 12248 11756 12257
rect 11796 12291 11848 12300
rect 11796 12257 11805 12291
rect 11805 12257 11839 12291
rect 11839 12257 11848 12291
rect 11796 12248 11848 12257
rect 17684 12248 17736 12300
rect 6184 12223 6236 12232
rect 6184 12189 6193 12223
rect 6193 12189 6227 12223
rect 6227 12189 6236 12223
rect 6184 12180 6236 12189
rect 6460 12112 6512 12164
rect 5264 12044 5316 12096
rect 4432 11942 4484 11994
rect 4496 11942 4548 11994
rect 4560 11942 4612 11994
rect 4624 11942 4676 11994
rect 11332 11942 11384 11994
rect 11396 11942 11448 11994
rect 11460 11942 11512 11994
rect 11524 11942 11576 11994
rect 18232 11942 18284 11994
rect 18296 11942 18348 11994
rect 18360 11942 18412 11994
rect 18424 11942 18476 11994
rect 10140 11840 10192 11892
rect 10508 11840 10560 11892
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 6828 11772 6880 11824
rect 7748 11772 7800 11824
rect 6644 11704 6696 11756
rect 5724 11679 5776 11688
rect 5724 11645 5733 11679
rect 5733 11645 5767 11679
rect 5767 11645 5776 11679
rect 5724 11636 5776 11645
rect 6184 11636 6236 11688
rect 8484 11704 8536 11756
rect 7748 11636 7800 11688
rect 8668 11636 8720 11688
rect 10048 11704 10100 11756
rect 10048 11611 10100 11620
rect 10048 11577 10057 11611
rect 10057 11577 10091 11611
rect 10091 11577 10100 11611
rect 10048 11568 10100 11577
rect 4988 11500 5040 11552
rect 6828 11500 6880 11552
rect 8208 11500 8260 11552
rect 9128 11500 9180 11552
rect 18420 11500 18472 11552
rect 7882 11398 7934 11450
rect 7946 11398 7998 11450
rect 8010 11398 8062 11450
rect 8074 11398 8126 11450
rect 14782 11398 14834 11450
rect 14846 11398 14898 11450
rect 14910 11398 14962 11450
rect 14974 11398 15026 11450
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 3516 11296 3568 11348
rect 7196 11296 7248 11348
rect 7564 11296 7616 11348
rect 2964 11203 3016 11212
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 2964 11169 2973 11203
rect 2973 11169 3007 11203
rect 3007 11169 3016 11203
rect 2964 11160 3016 11169
rect 6644 11160 6696 11212
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 7196 11160 7248 11169
rect 8208 11228 8260 11280
rect 7380 11160 7432 11212
rect 7748 11203 7800 11212
rect 7748 11169 7757 11203
rect 7757 11169 7791 11203
rect 7791 11169 7800 11203
rect 10508 11296 10560 11348
rect 18420 11339 18472 11348
rect 7748 11160 7800 11169
rect 2412 11024 2464 11076
rect 4160 11024 4212 11076
rect 8116 11092 8168 11144
rect 8668 11160 8720 11212
rect 10140 11228 10192 11280
rect 12072 11228 12124 11280
rect 13084 11228 13136 11280
rect 10416 11160 10468 11212
rect 11060 11160 11112 11212
rect 15016 11203 15068 11212
rect 15016 11169 15025 11203
rect 15025 11169 15059 11203
rect 15059 11169 15068 11203
rect 15016 11160 15068 11169
rect 17868 11228 17920 11280
rect 18420 11305 18429 11339
rect 18429 11305 18463 11339
rect 18463 11305 18472 11339
rect 18420 11296 18472 11305
rect 21272 11228 21324 11280
rect 17684 11160 17736 11212
rect 19340 11160 19392 11212
rect 11796 11135 11848 11144
rect 11796 11101 11805 11135
rect 11805 11101 11839 11135
rect 11839 11101 11848 11135
rect 11796 11092 11848 11101
rect 12072 11092 12124 11144
rect 15292 11092 15344 11144
rect 18052 11092 18104 11144
rect 21180 11092 21232 11144
rect 7380 11067 7432 11076
rect 7380 11033 7389 11067
rect 7389 11033 7423 11067
rect 7423 11033 7432 11067
rect 7380 11024 7432 11033
rect 7564 11024 7616 11076
rect 14832 11024 14884 11076
rect 15384 11024 15436 11076
rect 18788 11067 18840 11076
rect 18788 11033 18797 11067
rect 18797 11033 18831 11067
rect 18831 11033 18840 11067
rect 18788 11024 18840 11033
rect 20168 11024 20220 11076
rect 8300 10999 8352 11008
rect 8300 10965 8309 10999
rect 8309 10965 8343 10999
rect 8343 10965 8352 10999
rect 8300 10956 8352 10965
rect 10968 10956 11020 11008
rect 17224 10999 17276 11008
rect 17224 10965 17233 10999
rect 17233 10965 17267 10999
rect 17267 10965 17276 10999
rect 17224 10956 17276 10965
rect 4432 10854 4484 10906
rect 4496 10854 4548 10906
rect 4560 10854 4612 10906
rect 4624 10854 4676 10906
rect 11332 10854 11384 10906
rect 11396 10854 11448 10906
rect 11460 10854 11512 10906
rect 11524 10854 11576 10906
rect 18232 10854 18284 10906
rect 18296 10854 18348 10906
rect 18360 10854 18412 10906
rect 18424 10854 18476 10906
rect 4160 10752 4212 10804
rect 5356 10752 5408 10804
rect 6460 10684 6512 10736
rect 6736 10659 6788 10668
rect 6736 10625 6745 10659
rect 6745 10625 6779 10659
rect 6779 10625 6788 10659
rect 6736 10616 6788 10625
rect 11060 10752 11112 10804
rect 13820 10752 13872 10804
rect 15016 10752 15068 10804
rect 10048 10616 10100 10668
rect 12900 10616 12952 10668
rect 2688 10591 2740 10600
rect 2688 10557 2697 10591
rect 2697 10557 2731 10591
rect 2731 10557 2740 10591
rect 2688 10548 2740 10557
rect 4804 10591 4856 10600
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 6644 10591 6696 10600
rect 2872 10523 2924 10532
rect 2872 10489 2881 10523
rect 2881 10489 2915 10523
rect 2915 10489 2924 10523
rect 2872 10480 2924 10489
rect 6644 10557 6653 10591
rect 6653 10557 6687 10591
rect 6687 10557 6696 10591
rect 6644 10548 6696 10557
rect 6828 10591 6880 10600
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 8208 10548 8260 10600
rect 9128 10591 9180 10600
rect 9128 10557 9137 10591
rect 9137 10557 9171 10591
rect 9171 10557 9180 10591
rect 9128 10548 9180 10557
rect 5724 10480 5776 10532
rect 9496 10591 9548 10600
rect 9496 10557 9505 10591
rect 9505 10557 9539 10591
rect 9539 10557 9548 10591
rect 9496 10548 9548 10557
rect 13636 10548 13688 10600
rect 14832 10591 14884 10600
rect 14832 10557 14841 10591
rect 14841 10557 14875 10591
rect 14875 10557 14884 10591
rect 14832 10548 14884 10557
rect 15384 10591 15436 10600
rect 15384 10557 15393 10591
rect 15393 10557 15427 10591
rect 15427 10557 15436 10591
rect 15384 10548 15436 10557
rect 5448 10412 5500 10464
rect 8944 10455 8996 10464
rect 8944 10421 8953 10455
rect 8953 10421 8987 10455
rect 8987 10421 8996 10455
rect 8944 10412 8996 10421
rect 9588 10455 9640 10464
rect 9588 10421 9597 10455
rect 9597 10421 9631 10455
rect 9631 10421 9640 10455
rect 9588 10412 9640 10421
rect 17224 10795 17276 10804
rect 17224 10761 17233 10795
rect 17233 10761 17267 10795
rect 17267 10761 17276 10795
rect 17224 10752 17276 10761
rect 17684 10795 17736 10804
rect 17684 10761 17693 10795
rect 17693 10761 17727 10795
rect 17727 10761 17736 10795
rect 17684 10752 17736 10761
rect 19248 10752 19300 10804
rect 19800 10752 19852 10804
rect 17868 10684 17920 10736
rect 18052 10616 18104 10668
rect 19156 10659 19208 10668
rect 19156 10625 19165 10659
rect 19165 10625 19199 10659
rect 19199 10625 19208 10659
rect 19156 10616 19208 10625
rect 17960 10480 18012 10532
rect 20168 10480 20220 10532
rect 16764 10412 16816 10464
rect 18880 10412 18932 10464
rect 7882 10310 7934 10362
rect 7946 10310 7998 10362
rect 8010 10310 8062 10362
rect 8074 10310 8126 10362
rect 14782 10310 14834 10362
rect 14846 10310 14898 10362
rect 14910 10310 14962 10362
rect 14974 10310 15026 10362
rect 1492 10251 1544 10260
rect 1492 10217 1501 10251
rect 1501 10217 1535 10251
rect 1535 10217 1544 10251
rect 1492 10208 1544 10217
rect 5080 10208 5132 10260
rect 6368 10251 6420 10260
rect 6368 10217 6377 10251
rect 6377 10217 6411 10251
rect 6411 10217 6420 10251
rect 6368 10208 6420 10217
rect 9772 10208 9824 10260
rect 12072 10208 12124 10260
rect 13636 10251 13688 10260
rect 13636 10217 13645 10251
rect 13645 10217 13679 10251
rect 13679 10217 13688 10251
rect 13636 10208 13688 10217
rect 17224 10208 17276 10260
rect 19156 10208 19208 10260
rect 21272 10251 21324 10260
rect 21272 10217 21281 10251
rect 21281 10217 21315 10251
rect 21315 10217 21324 10251
rect 21272 10208 21324 10217
rect 5448 10183 5500 10192
rect 5448 10149 5457 10183
rect 5457 10149 5491 10183
rect 5491 10149 5500 10183
rect 5448 10140 5500 10149
rect 9128 10140 9180 10192
rect 1676 10072 1728 10124
rect 6828 10072 6880 10124
rect 9772 10115 9824 10124
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 9220 10047 9272 10056
rect 9220 10013 9229 10047
rect 9229 10013 9263 10047
rect 9263 10013 9272 10047
rect 9220 10004 9272 10013
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 10048 10115 10100 10124
rect 10048 10081 10057 10115
rect 10057 10081 10091 10115
rect 10091 10081 10100 10115
rect 10048 10072 10100 10081
rect 13820 10140 13872 10192
rect 12900 10115 12952 10124
rect 12900 10081 12909 10115
rect 12909 10081 12943 10115
rect 12943 10081 12952 10115
rect 12900 10072 12952 10081
rect 13452 10115 13504 10124
rect 13452 10081 13461 10115
rect 13461 10081 13495 10115
rect 13495 10081 13504 10115
rect 13452 10072 13504 10081
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 21456 10115 21508 10124
rect 13544 10072 13596 10081
rect 21456 10081 21465 10115
rect 21465 10081 21499 10115
rect 21499 10081 21508 10115
rect 21456 10072 21508 10081
rect 10324 9936 10376 9988
rect 5908 9911 5960 9920
rect 5908 9877 5917 9911
rect 5917 9877 5951 9911
rect 5951 9877 5960 9911
rect 5908 9868 5960 9877
rect 13360 9868 13412 9920
rect 4432 9766 4484 9818
rect 4496 9766 4548 9818
rect 4560 9766 4612 9818
rect 4624 9766 4676 9818
rect 11332 9766 11384 9818
rect 11396 9766 11448 9818
rect 11460 9766 11512 9818
rect 11524 9766 11576 9818
rect 18232 9766 18284 9818
rect 18296 9766 18348 9818
rect 18360 9766 18412 9818
rect 18424 9766 18476 9818
rect 2412 9571 2464 9580
rect 2412 9537 2421 9571
rect 2421 9537 2455 9571
rect 2455 9537 2464 9571
rect 2412 9528 2464 9537
rect 7288 9528 7340 9580
rect 2596 9460 2648 9512
rect 2872 9460 2924 9512
rect 4988 9503 5040 9512
rect 4988 9469 4997 9503
rect 4997 9469 5031 9503
rect 5031 9469 5040 9503
rect 4988 9460 5040 9469
rect 9220 9528 9272 9580
rect 9680 9571 9732 9580
rect 2228 9435 2280 9444
rect 2228 9401 2237 9435
rect 2237 9401 2271 9435
rect 2271 9401 2280 9435
rect 2228 9392 2280 9401
rect 4620 9392 4672 9444
rect 5172 9392 5224 9444
rect 8392 9392 8444 9444
rect 9680 9537 9689 9571
rect 9689 9537 9723 9571
rect 9723 9537 9732 9571
rect 9680 9528 9732 9537
rect 9588 9460 9640 9512
rect 10968 9528 11020 9580
rect 10416 9503 10468 9512
rect 10416 9469 10425 9503
rect 10425 9469 10459 9503
rect 10459 9469 10468 9503
rect 10416 9460 10468 9469
rect 9680 9392 9732 9444
rect 12440 9460 12492 9512
rect 13452 9460 13504 9512
rect 12072 9392 12124 9444
rect 2734 9367 2786 9376
rect 2734 9333 2743 9367
rect 2743 9333 2777 9367
rect 2777 9333 2786 9367
rect 2734 9324 2786 9333
rect 4804 9367 4856 9376
rect 4804 9333 4813 9367
rect 4813 9333 4847 9367
rect 4847 9333 4856 9367
rect 4804 9324 4856 9333
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10140 9324 10192 9333
rect 13544 9324 13596 9376
rect 7882 9222 7934 9274
rect 7946 9222 7998 9274
rect 8010 9222 8062 9274
rect 8074 9222 8126 9274
rect 14782 9222 14834 9274
rect 14846 9222 14898 9274
rect 14910 9222 14962 9274
rect 14974 9222 15026 9274
rect 2228 9120 2280 9172
rect 2688 9163 2740 9172
rect 2688 9129 2697 9163
rect 2697 9129 2731 9163
rect 2731 9129 2740 9163
rect 2688 9120 2740 9129
rect 6736 9120 6788 9172
rect 1584 9052 1636 9104
rect 4620 8848 4672 8900
rect 5356 8984 5408 9036
rect 6736 8984 6788 9036
rect 10416 9120 10468 9172
rect 15476 9120 15528 9172
rect 10968 9052 11020 9104
rect 12440 9052 12492 9104
rect 16764 9095 16816 9104
rect 16764 9061 16773 9095
rect 16773 9061 16807 9095
rect 16807 9061 16816 9095
rect 16764 9052 16816 9061
rect 10416 8984 10468 9036
rect 12072 8984 12124 9036
rect 18604 8984 18656 9036
rect 8392 8916 8444 8968
rect 15292 8916 15344 8968
rect 8300 8848 8352 8900
rect 1768 8780 1820 8832
rect 2688 8780 2740 8832
rect 3516 8780 3568 8832
rect 3608 8780 3660 8832
rect 9588 8823 9640 8832
rect 9588 8789 9597 8823
rect 9597 8789 9631 8823
rect 9631 8789 9640 8823
rect 9588 8780 9640 8789
rect 9864 8823 9916 8832
rect 9864 8789 9873 8823
rect 9873 8789 9907 8823
rect 9907 8789 9916 8823
rect 9864 8780 9916 8789
rect 15108 8780 15160 8832
rect 16856 8823 16908 8832
rect 16856 8789 16865 8823
rect 16865 8789 16899 8823
rect 16899 8789 16908 8823
rect 16856 8780 16908 8789
rect 17316 8780 17368 8832
rect 4432 8678 4484 8730
rect 4496 8678 4548 8730
rect 4560 8678 4612 8730
rect 4624 8678 4676 8730
rect 11332 8678 11384 8730
rect 11396 8678 11448 8730
rect 11460 8678 11512 8730
rect 11524 8678 11576 8730
rect 18232 8678 18284 8730
rect 18296 8678 18348 8730
rect 18360 8678 18412 8730
rect 18424 8678 18476 8730
rect 2136 8619 2188 8628
rect 2136 8585 2145 8619
rect 2145 8585 2179 8619
rect 2179 8585 2188 8619
rect 16764 8619 16816 8628
rect 2136 8576 2188 8585
rect 16764 8585 16773 8619
rect 16773 8585 16807 8619
rect 16807 8585 16816 8619
rect 16764 8576 16816 8585
rect 2688 8483 2740 8492
rect 2688 8449 2697 8483
rect 2697 8449 2731 8483
rect 2731 8449 2740 8483
rect 2688 8440 2740 8449
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 10416 8440 10468 8492
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 3608 8372 3660 8424
rect 5172 8372 5224 8424
rect 8392 8372 8444 8424
rect 10968 8372 11020 8424
rect 12072 8415 12124 8424
rect 12072 8381 12081 8415
rect 12081 8381 12115 8415
rect 12115 8381 12124 8415
rect 12072 8372 12124 8381
rect 17316 8483 17368 8492
rect 17316 8449 17325 8483
rect 17325 8449 17359 8483
rect 17359 8449 17368 8483
rect 17316 8440 17368 8449
rect 16856 8372 16908 8424
rect 18788 8483 18840 8492
rect 18788 8449 18797 8483
rect 18797 8449 18831 8483
rect 18831 8449 18840 8483
rect 18788 8440 18840 8449
rect 21456 8415 21508 8424
rect 21456 8381 21465 8415
rect 21465 8381 21499 8415
rect 21499 8381 21508 8415
rect 21456 8372 21508 8381
rect 3976 8304 4028 8356
rect 6644 8347 6696 8356
rect 6644 8313 6653 8347
rect 6653 8313 6687 8347
rect 6687 8313 6696 8347
rect 6644 8304 6696 8313
rect 12808 8304 12860 8356
rect 18604 8304 18656 8356
rect 21272 8279 21324 8288
rect 21272 8245 21281 8279
rect 21281 8245 21315 8279
rect 21315 8245 21324 8279
rect 21272 8236 21324 8245
rect 7882 8134 7934 8186
rect 7946 8134 7998 8186
rect 8010 8134 8062 8186
rect 8074 8134 8126 8186
rect 14782 8134 14834 8186
rect 14846 8134 14898 8186
rect 14910 8134 14962 8186
rect 14974 8134 15026 8186
rect 8576 8032 8628 8084
rect 12808 8075 12860 8084
rect 12808 8041 12817 8075
rect 12817 8041 12851 8075
rect 12851 8041 12860 8075
rect 12808 8032 12860 8041
rect 8392 8007 8444 8016
rect 8392 7973 8401 8007
rect 8401 7973 8435 8007
rect 8435 7973 8444 8007
rect 8392 7964 8444 7973
rect 2136 7939 2188 7948
rect 2136 7905 2145 7939
rect 2145 7905 2179 7939
rect 2179 7905 2188 7939
rect 2136 7896 2188 7905
rect 2596 7896 2648 7948
rect 7656 7939 7708 7948
rect 7656 7905 7665 7939
rect 7665 7905 7699 7939
rect 7699 7905 7708 7939
rect 7656 7896 7708 7905
rect 8576 7939 8628 7948
rect 8576 7905 8585 7939
rect 8585 7905 8619 7939
rect 8619 7905 8628 7939
rect 8576 7896 8628 7905
rect 10232 7896 10284 7948
rect 9772 7828 9824 7880
rect 3976 7692 4028 7744
rect 9404 7692 9456 7744
rect 9496 7692 9548 7744
rect 12348 7692 12400 7744
rect 14372 7939 14424 7948
rect 14372 7905 14381 7939
rect 14381 7905 14415 7939
rect 14415 7905 14424 7939
rect 14372 7896 14424 7905
rect 14464 7939 14516 7948
rect 14464 7905 14473 7939
rect 14473 7905 14507 7939
rect 14507 7905 14516 7939
rect 16764 7964 16816 8016
rect 14464 7896 14516 7905
rect 13728 7828 13780 7880
rect 14372 7760 14424 7812
rect 21272 7828 21324 7880
rect 4432 7590 4484 7642
rect 4496 7590 4548 7642
rect 4560 7590 4612 7642
rect 4624 7590 4676 7642
rect 11332 7590 11384 7642
rect 11396 7590 11448 7642
rect 11460 7590 11512 7642
rect 11524 7590 11576 7642
rect 18232 7590 18284 7642
rect 18296 7590 18348 7642
rect 18360 7590 18412 7642
rect 18424 7590 18476 7642
rect 7656 7531 7708 7540
rect 7656 7497 7665 7531
rect 7665 7497 7699 7531
rect 7699 7497 7708 7531
rect 7656 7488 7708 7497
rect 12716 7488 12768 7540
rect 2964 7420 3016 7472
rect 8576 7395 8628 7404
rect 8576 7361 8585 7395
rect 8585 7361 8619 7395
rect 8619 7361 8628 7395
rect 8576 7352 8628 7361
rect 9404 7352 9456 7404
rect 9496 7327 9548 7336
rect 3884 7259 3936 7268
rect 3884 7225 3893 7259
rect 3893 7225 3927 7259
rect 3927 7225 3936 7259
rect 3884 7216 3936 7225
rect 9496 7293 9505 7327
rect 9505 7293 9539 7327
rect 9539 7293 9548 7327
rect 9496 7284 9548 7293
rect 12348 7352 12400 7404
rect 10416 7327 10468 7336
rect 10416 7293 10425 7327
rect 10425 7293 10459 7327
rect 10459 7293 10468 7327
rect 10416 7284 10468 7293
rect 14372 7352 14424 7404
rect 14464 7284 14516 7336
rect 10600 7259 10652 7268
rect 10600 7225 10609 7259
rect 10609 7225 10643 7259
rect 10643 7225 10652 7259
rect 10600 7216 10652 7225
rect 7882 7046 7934 7098
rect 7946 7046 7998 7098
rect 8010 7046 8062 7098
rect 8074 7046 8126 7098
rect 14782 7046 14834 7098
rect 14846 7046 14898 7098
rect 14910 7046 14962 7098
rect 14974 7046 15026 7098
rect 8300 6987 8352 6996
rect 8300 6953 8309 6987
rect 8309 6953 8343 6987
rect 8343 6953 8352 6987
rect 8300 6944 8352 6953
rect 8576 6944 8628 6996
rect 3884 6740 3936 6792
rect 10232 6876 10284 6928
rect 5540 6808 5592 6860
rect 6184 6808 6236 6860
rect 5264 6783 5316 6792
rect 5264 6749 5273 6783
rect 5273 6749 5307 6783
rect 5307 6749 5316 6783
rect 5264 6740 5316 6749
rect 8484 6808 8536 6860
rect 9772 6808 9824 6860
rect 10140 6808 10192 6860
rect 10600 6808 10652 6860
rect 11152 6851 11204 6860
rect 11152 6817 11161 6851
rect 11161 6817 11195 6851
rect 11195 6817 11204 6851
rect 11152 6808 11204 6817
rect 15936 6851 15988 6860
rect 15936 6817 15945 6851
rect 15945 6817 15979 6851
rect 15979 6817 15988 6851
rect 15936 6808 15988 6817
rect 17224 6808 17276 6860
rect 16212 6783 16264 6792
rect 16212 6749 16221 6783
rect 16221 6749 16255 6783
rect 16255 6749 16264 6783
rect 16212 6740 16264 6749
rect 1676 6604 1728 6656
rect 4432 6502 4484 6554
rect 4496 6502 4548 6554
rect 4560 6502 4612 6554
rect 4624 6502 4676 6554
rect 11332 6502 11384 6554
rect 11396 6502 11448 6554
rect 11460 6502 11512 6554
rect 11524 6502 11576 6554
rect 18232 6502 18284 6554
rect 18296 6502 18348 6554
rect 18360 6502 18412 6554
rect 18424 6502 18476 6554
rect 3884 6196 3936 6248
rect 5540 6239 5592 6248
rect 5540 6205 5549 6239
rect 5549 6205 5583 6239
rect 5583 6205 5592 6239
rect 5540 6196 5592 6205
rect 5908 6196 5960 6248
rect 6920 6196 6972 6248
rect 16212 6264 16264 6316
rect 18236 6264 18288 6316
rect 17592 6239 17644 6248
rect 17592 6205 17601 6239
rect 17601 6205 17635 6239
rect 17635 6205 17644 6239
rect 17592 6196 17644 6205
rect 6184 6128 6236 6180
rect 18052 6196 18104 6248
rect 18420 6196 18472 6248
rect 2780 6060 2832 6112
rect 18696 6128 18748 6180
rect 17408 6060 17460 6112
rect 18604 6060 18656 6112
rect 7882 5958 7934 6010
rect 7946 5958 7998 6010
rect 8010 5958 8062 6010
rect 8074 5958 8126 6010
rect 14782 5958 14834 6010
rect 14846 5958 14898 6010
rect 14910 5958 14962 6010
rect 14974 5958 15026 6010
rect 6920 5899 6972 5908
rect 6920 5865 6929 5899
rect 6929 5865 6963 5899
rect 6963 5865 6972 5899
rect 6920 5856 6972 5865
rect 15936 5856 15988 5908
rect 4988 5788 5040 5840
rect 12716 5831 12768 5840
rect 12716 5797 12725 5831
rect 12725 5797 12759 5831
rect 12759 5797 12768 5831
rect 12716 5788 12768 5797
rect 2780 5763 2832 5772
rect 2780 5729 2789 5763
rect 2789 5729 2823 5763
rect 2823 5729 2832 5763
rect 7012 5763 7064 5772
rect 2780 5720 2832 5729
rect 7012 5729 7021 5763
rect 7021 5729 7055 5763
rect 7055 5729 7064 5763
rect 7012 5720 7064 5729
rect 14832 5720 14884 5772
rect 15108 5763 15160 5772
rect 15108 5729 15117 5763
rect 15117 5729 15151 5763
rect 15151 5729 15160 5763
rect 15108 5720 15160 5729
rect 16948 5720 17000 5772
rect 17408 5763 17460 5772
rect 17408 5729 17417 5763
rect 17417 5729 17451 5763
rect 17451 5729 17460 5763
rect 17408 5720 17460 5729
rect 15200 5695 15252 5704
rect 15200 5661 15209 5695
rect 15209 5661 15243 5695
rect 15243 5661 15252 5695
rect 15200 5652 15252 5661
rect 15292 5652 15344 5704
rect 17592 5788 17644 5840
rect 18052 5720 18104 5772
rect 18420 5720 18472 5772
rect 18696 5763 18748 5772
rect 17960 5652 18012 5704
rect 18236 5652 18288 5704
rect 18696 5729 18705 5763
rect 18705 5729 18739 5763
rect 18739 5729 18748 5763
rect 18696 5720 18748 5729
rect 20812 5720 20864 5772
rect 21456 5763 21508 5772
rect 21456 5729 21465 5763
rect 21465 5729 21499 5763
rect 21499 5729 21508 5763
rect 21456 5720 21508 5729
rect 9680 5584 9732 5636
rect 18696 5584 18748 5636
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 2688 5559 2740 5568
rect 2688 5525 2697 5559
rect 2697 5525 2731 5559
rect 2731 5525 2740 5559
rect 2688 5516 2740 5525
rect 14740 5516 14792 5568
rect 4432 5414 4484 5466
rect 4496 5414 4548 5466
rect 4560 5414 4612 5466
rect 4624 5414 4676 5466
rect 11332 5414 11384 5466
rect 11396 5414 11448 5466
rect 11460 5414 11512 5466
rect 11524 5414 11576 5466
rect 18232 5414 18284 5466
rect 18296 5414 18348 5466
rect 18360 5414 18412 5466
rect 18424 5414 18476 5466
rect 7012 5312 7064 5364
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3240 5176 3292 5185
rect 2044 5108 2096 5160
rect 2688 5108 2740 5160
rect 7012 5108 7064 5160
rect 7748 5176 7800 5228
rect 9680 5176 9732 5228
rect 15200 5312 15252 5364
rect 16948 5355 17000 5364
rect 16948 5321 16957 5355
rect 16957 5321 16991 5355
rect 16991 5321 17000 5355
rect 16948 5312 17000 5321
rect 18052 5355 18104 5364
rect 18052 5321 18061 5355
rect 18061 5321 18095 5355
rect 18095 5321 18104 5355
rect 18052 5312 18104 5321
rect 9128 5108 9180 5160
rect 10324 5151 10376 5160
rect 10324 5117 10333 5151
rect 10333 5117 10367 5151
rect 10367 5117 10376 5151
rect 10324 5108 10376 5117
rect 17960 5176 18012 5228
rect 12348 5108 12400 5160
rect 12992 5151 13044 5160
rect 6276 5040 6328 5092
rect 11152 5040 11204 5092
rect 11888 5040 11940 5092
rect 12992 5117 13001 5151
rect 13001 5117 13035 5151
rect 13035 5117 13044 5151
rect 12992 5108 13044 5117
rect 14740 5151 14792 5160
rect 14740 5117 14749 5151
rect 14749 5117 14783 5151
rect 14783 5117 14792 5151
rect 14740 5108 14792 5117
rect 14832 5108 14884 5160
rect 15384 5108 15436 5160
rect 18052 5108 18104 5160
rect 18696 5108 18748 5160
rect 13176 5040 13228 5092
rect 7012 4972 7064 5024
rect 15292 4972 15344 5024
rect 17316 5015 17368 5024
rect 17316 4981 17325 5015
rect 17325 4981 17359 5015
rect 17359 4981 17368 5015
rect 17316 4972 17368 4981
rect 17408 5015 17460 5024
rect 17408 4981 17417 5015
rect 17417 4981 17451 5015
rect 17451 4981 17460 5015
rect 17408 4972 17460 4981
rect 7882 4870 7934 4922
rect 7946 4870 7998 4922
rect 8010 4870 8062 4922
rect 8074 4870 8126 4922
rect 14782 4870 14834 4922
rect 14846 4870 14898 4922
rect 14910 4870 14962 4922
rect 14974 4870 15026 4922
rect 7748 4768 7800 4820
rect 9864 4811 9916 4820
rect 9864 4777 9873 4811
rect 9873 4777 9907 4811
rect 9907 4777 9916 4811
rect 9864 4768 9916 4777
rect 12348 4768 12400 4820
rect 17316 4768 17368 4820
rect 6276 4700 6328 4752
rect 6828 4700 6880 4752
rect 7380 4700 7432 4752
rect 11152 4743 11204 4752
rect 11152 4709 11161 4743
rect 11161 4709 11195 4743
rect 11195 4709 11204 4743
rect 11152 4700 11204 4709
rect 18972 4700 19024 4752
rect 4988 4675 5040 4684
rect 4988 4641 4997 4675
rect 4997 4641 5031 4675
rect 5031 4641 5040 4675
rect 4988 4632 5040 4641
rect 7012 4675 7064 4684
rect 7012 4641 7021 4675
rect 7021 4641 7055 4675
rect 7055 4641 7064 4675
rect 7012 4632 7064 4641
rect 10324 4632 10376 4684
rect 11704 4632 11756 4684
rect 19156 4632 19208 4684
rect 8484 4607 8536 4616
rect 8484 4573 8493 4607
rect 8493 4573 8527 4607
rect 8527 4573 8536 4607
rect 8484 4564 8536 4573
rect 9680 4564 9732 4616
rect 18604 4607 18656 4616
rect 18604 4573 18613 4607
rect 18613 4573 18647 4607
rect 18647 4573 18656 4607
rect 18604 4564 18656 4573
rect 7104 4496 7156 4548
rect 8208 4496 8260 4548
rect 4432 4326 4484 4378
rect 4496 4326 4548 4378
rect 4560 4326 4612 4378
rect 4624 4326 4676 4378
rect 11332 4326 11384 4378
rect 11396 4326 11448 4378
rect 11460 4326 11512 4378
rect 11524 4326 11576 4378
rect 18232 4326 18284 4378
rect 18296 4326 18348 4378
rect 18360 4326 18412 4378
rect 18424 4326 18476 4378
rect 7104 4224 7156 4276
rect 16948 4224 17000 4276
rect 17408 4224 17460 4276
rect 15384 4199 15436 4208
rect 15384 4165 15393 4199
rect 15393 4165 15427 4199
rect 15427 4165 15436 4199
rect 15384 4156 15436 4165
rect 18972 4156 19024 4208
rect 21088 4156 21140 4208
rect 15108 3952 15160 4004
rect 7564 3884 7616 3936
rect 11980 3884 12032 3936
rect 7882 3782 7934 3834
rect 7946 3782 7998 3834
rect 8010 3782 8062 3834
rect 8074 3782 8126 3834
rect 14782 3782 14834 3834
rect 14846 3782 14898 3834
rect 14910 3782 14962 3834
rect 14974 3782 15026 3834
rect 9496 3680 9548 3732
rect 11152 3680 11204 3732
rect 14464 3680 14516 3732
rect 15108 3723 15160 3732
rect 15108 3689 15117 3723
rect 15117 3689 15151 3723
rect 15151 3689 15160 3723
rect 15108 3680 15160 3689
rect 3976 3655 4028 3664
rect 3976 3621 3985 3655
rect 3985 3621 4019 3655
rect 4019 3621 4028 3655
rect 3976 3612 4028 3621
rect 9128 3655 9180 3664
rect 9128 3621 9137 3655
rect 9137 3621 9171 3655
rect 9171 3621 9180 3655
rect 9128 3612 9180 3621
rect 11704 3612 11756 3664
rect 6736 3587 6788 3596
rect 6736 3553 6745 3587
rect 6745 3553 6779 3587
rect 6779 3553 6788 3587
rect 6736 3544 6788 3553
rect 6828 3544 6880 3596
rect 11888 3587 11940 3596
rect 9036 3476 9088 3528
rect 10968 3519 11020 3528
rect 10968 3485 10977 3519
rect 10977 3485 11011 3519
rect 11011 3485 11020 3519
rect 10968 3476 11020 3485
rect 11888 3553 11897 3587
rect 11897 3553 11931 3587
rect 11931 3553 11940 3587
rect 11888 3544 11940 3553
rect 17960 3612 18012 3664
rect 13820 3476 13872 3528
rect 15568 3476 15620 3528
rect 9772 3408 9824 3460
rect 14556 3408 14608 3460
rect 11796 3340 11848 3392
rect 11980 3340 12032 3392
rect 15936 3340 15988 3392
rect 4432 3238 4484 3290
rect 4496 3238 4548 3290
rect 4560 3238 4612 3290
rect 4624 3238 4676 3290
rect 11332 3238 11384 3290
rect 11396 3238 11448 3290
rect 11460 3238 11512 3290
rect 11524 3238 11576 3290
rect 18232 3238 18284 3290
rect 18296 3238 18348 3290
rect 18360 3238 18412 3290
rect 18424 3238 18476 3290
rect 9036 3179 9088 3188
rect 9036 3145 9045 3179
rect 9045 3145 9079 3179
rect 9079 3145 9088 3179
rect 9036 3136 9088 3145
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 11152 3136 11204 3188
rect 12440 3136 12492 3188
rect 13820 3179 13872 3188
rect 13820 3145 13829 3179
rect 13829 3145 13863 3179
rect 13863 3145 13872 3179
rect 13820 3136 13872 3145
rect 14556 3179 14608 3188
rect 14556 3145 14565 3179
rect 14565 3145 14599 3179
rect 14599 3145 14608 3179
rect 14556 3136 14608 3145
rect 15108 3136 15160 3188
rect 15568 3179 15620 3188
rect 15568 3145 15577 3179
rect 15577 3145 15611 3179
rect 15611 3145 15620 3179
rect 15568 3136 15620 3145
rect 18972 3136 19024 3188
rect 19156 3179 19208 3188
rect 19156 3145 19165 3179
rect 19165 3145 19199 3179
rect 19199 3145 19208 3179
rect 19156 3136 19208 3145
rect 8484 3043 8536 3052
rect 8484 3009 8493 3043
rect 8493 3009 8527 3043
rect 8527 3009 8536 3043
rect 8484 3000 8536 3009
rect 1400 2975 1452 2984
rect 1400 2941 1409 2975
rect 1409 2941 1443 2975
rect 1443 2941 1452 2975
rect 1400 2932 1452 2941
rect 8944 2932 8996 2984
rect 14464 3111 14516 3120
rect 9496 3043 9548 3052
rect 9496 3009 9505 3043
rect 9505 3009 9539 3043
rect 9539 3009 9548 3043
rect 9496 3000 9548 3009
rect 9864 2932 9916 2984
rect 10508 3000 10560 3052
rect 14464 3077 14473 3111
rect 14473 3077 14507 3111
rect 14507 3077 14516 3111
rect 14464 3068 14516 3077
rect 10968 2932 11020 2984
rect 11888 2932 11940 2984
rect 12532 2975 12584 2984
rect 12532 2941 12541 2975
rect 12541 2941 12575 2975
rect 12575 2941 12584 2975
rect 12532 2932 12584 2941
rect 13452 2975 13504 2984
rect 13452 2941 13461 2975
rect 13461 2941 13495 2975
rect 13495 2941 13504 2975
rect 13452 2932 13504 2941
rect 13820 2932 13872 2984
rect 11796 2864 11848 2916
rect 16120 3043 16172 3052
rect 16120 3009 16129 3043
rect 16129 3009 16163 3043
rect 16163 3009 16172 3043
rect 16120 3000 16172 3009
rect 16948 3043 17000 3052
rect 16948 3009 16957 3043
rect 16957 3009 16991 3043
rect 16991 3009 17000 3043
rect 16948 3000 17000 3009
rect 17960 3000 18012 3052
rect 20904 3043 20956 3052
rect 15936 2975 15988 2984
rect 15936 2941 15945 2975
rect 15945 2941 15979 2975
rect 15979 2941 15988 2975
rect 15936 2932 15988 2941
rect 16120 2864 16172 2916
rect 20904 3009 20913 3043
rect 20913 3009 20947 3043
rect 20947 3009 20956 3043
rect 20904 3000 20956 3009
rect 21180 3043 21232 3052
rect 21180 3009 21189 3043
rect 21189 3009 21223 3043
rect 21223 3009 21232 3043
rect 21180 3000 21232 3009
rect 18972 2975 19024 2984
rect 18972 2941 18981 2975
rect 18981 2941 19015 2975
rect 19015 2941 19024 2975
rect 18972 2932 19024 2941
rect 21456 2975 21508 2984
rect 21456 2941 21465 2975
rect 21465 2941 21499 2975
rect 21499 2941 21508 2975
rect 21456 2932 21508 2941
rect 12164 2839 12216 2848
rect 12164 2805 12173 2839
rect 12173 2805 12207 2839
rect 12207 2805 12216 2839
rect 12164 2796 12216 2805
rect 13820 2796 13872 2848
rect 7882 2694 7934 2746
rect 7946 2694 7998 2746
rect 8010 2694 8062 2746
rect 8074 2694 8126 2746
rect 14782 2694 14834 2746
rect 14846 2694 14898 2746
rect 14910 2694 14962 2746
rect 14974 2694 15026 2746
rect 4804 2592 4856 2644
rect 6644 2592 6696 2644
rect 6736 2592 6788 2644
rect 9680 2592 9732 2644
rect 12164 2635 12216 2644
rect 12164 2601 12173 2635
rect 12173 2601 12207 2635
rect 12207 2601 12216 2635
rect 12164 2592 12216 2601
rect 13820 2635 13872 2644
rect 13820 2601 13829 2635
rect 13829 2601 13863 2635
rect 13863 2601 13872 2635
rect 13820 2592 13872 2601
rect 17500 2592 17552 2644
rect 18880 2635 18932 2644
rect 18880 2601 18889 2635
rect 18889 2601 18923 2635
rect 18923 2601 18932 2635
rect 18880 2592 18932 2601
rect 2044 2567 2096 2576
rect 2044 2533 2053 2567
rect 2053 2533 2087 2567
rect 2087 2533 2096 2567
rect 2044 2524 2096 2533
rect 8208 2524 8260 2576
rect 480 2456 532 2508
rect 3700 2456 3752 2508
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 6920 2456 6972 2508
rect 8760 2499 8812 2508
rect 8760 2465 8769 2499
rect 8769 2465 8803 2499
rect 8803 2465 8812 2499
rect 8760 2456 8812 2465
rect 10600 2456 10652 2508
rect 11980 2499 12032 2508
rect 11980 2465 11989 2499
rect 11989 2465 12023 2499
rect 12023 2465 12032 2499
rect 11980 2456 12032 2465
rect 13820 2456 13872 2508
rect 15660 2499 15712 2508
rect 15660 2465 15669 2499
rect 15669 2465 15703 2499
rect 15703 2465 15712 2499
rect 15660 2456 15712 2465
rect 17040 2456 17092 2508
rect 18880 2456 18932 2508
rect 20904 2499 20956 2508
rect 20904 2465 20913 2499
rect 20913 2465 20947 2499
rect 20947 2465 20956 2499
rect 20904 2456 20956 2465
rect 22100 2456 22152 2508
rect 12532 2388 12584 2440
rect 16120 2431 16172 2440
rect 16120 2397 16129 2431
rect 16129 2397 16163 2431
rect 16163 2397 16172 2431
rect 16120 2388 16172 2397
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 18052 2320 18104 2372
rect 20720 2363 20772 2372
rect 20720 2329 20729 2363
rect 20729 2329 20763 2363
rect 20763 2329 20772 2363
rect 20720 2320 20772 2329
rect 4432 2150 4484 2202
rect 4496 2150 4548 2202
rect 4560 2150 4612 2202
rect 4624 2150 4676 2202
rect 11332 2150 11384 2202
rect 11396 2150 11448 2202
rect 11460 2150 11512 2202
rect 11524 2150 11576 2202
rect 18232 2150 18284 2202
rect 18296 2150 18348 2202
rect 18360 2150 18412 2202
rect 18424 2150 18476 2202
<< metal2 >>
rect 938 24323 994 25123
rect 2778 24323 2834 25123
rect 4618 24323 4674 25123
rect 5998 24323 6054 25123
rect 7838 24323 7894 25123
rect 9678 24323 9734 25123
rect 11518 24323 11574 25123
rect 12898 24323 12954 25123
rect 14738 24323 14794 25123
rect 16578 24323 16634 25123
rect 17958 24323 18014 25123
rect 19798 24323 19854 25123
rect 21638 24323 21694 25123
rect 952 22574 980 24323
rect 1490 23216 1546 23225
rect 1490 23151 1546 23160
rect 1504 22778 1532 23151
rect 1492 22772 1544 22778
rect 1492 22714 1544 22720
rect 2792 22574 2820 24323
rect 4632 23066 4660 24323
rect 4632 23038 4844 23066
rect 4406 22876 4702 22896
rect 4462 22874 4486 22876
rect 4542 22874 4566 22876
rect 4622 22874 4646 22876
rect 4484 22822 4486 22874
rect 4548 22822 4560 22874
rect 4622 22822 4624 22874
rect 4462 22820 4486 22822
rect 4542 22820 4566 22822
rect 4622 22820 4646 22822
rect 4406 22800 4702 22820
rect 4816 22574 4844 23038
rect 4896 22704 4948 22710
rect 4896 22646 4948 22652
rect 940 22568 992 22574
rect 940 22510 992 22516
rect 2780 22568 2832 22574
rect 2780 22510 2832 22516
rect 4804 22568 4856 22574
rect 4804 22510 4856 22516
rect 1584 22500 1636 22506
rect 1584 22442 1636 22448
rect 1596 21690 1624 22442
rect 2044 22432 2096 22438
rect 2044 22374 2096 22380
rect 4804 22432 4856 22438
rect 4804 22374 4856 22380
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1398 20496 1454 20505
rect 1398 20431 1454 20440
rect 1412 20398 1440 20431
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1492 20256 1544 20262
rect 1492 20198 1544 20204
rect 1398 17776 1454 17785
rect 1398 17711 1400 17720
rect 1452 17711 1454 17720
rect 1400 17682 1452 17688
rect 1398 15736 1454 15745
rect 1398 15671 1454 15680
rect 1412 15570 1440 15671
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1504 13138 1532 20198
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 1596 13530 1624 17478
rect 1952 16040 2004 16046
rect 1952 15982 2004 15988
rect 1964 15502 1992 15982
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1780 13326 1808 14894
rect 1768 13320 1820 13326
rect 1768 13262 1820 13268
rect 1504 13110 1624 13138
rect 1490 13016 1546 13025
rect 1490 12951 1492 12960
rect 1544 12951 1546 12960
rect 1492 12922 1544 12928
rect 1490 10296 1546 10305
rect 1490 10231 1492 10240
rect 1544 10231 1546 10240
rect 1492 10202 1544 10208
rect 1596 9110 1624 13110
rect 1780 11150 1808 13262
rect 1872 11354 1900 15302
rect 1964 15162 1992 15438
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 2056 15026 2084 22374
rect 3700 22092 3752 22098
rect 3700 22034 3752 22040
rect 2504 21480 2556 21486
rect 2504 21422 2556 21428
rect 2516 20398 2544 21422
rect 2504 20392 2556 20398
rect 2504 20334 2556 20340
rect 2516 18290 2544 20334
rect 3516 20324 3568 20330
rect 3516 20266 3568 20272
rect 3528 20058 3556 20266
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3712 19922 3740 22034
rect 4160 21888 4212 21894
rect 4160 21830 4212 21836
rect 4172 21554 4200 21830
rect 4406 21788 4702 21808
rect 4462 21786 4486 21788
rect 4542 21786 4566 21788
rect 4622 21786 4646 21788
rect 4484 21734 4486 21786
rect 4548 21734 4560 21786
rect 4622 21734 4624 21786
rect 4462 21732 4486 21734
rect 4542 21732 4566 21734
rect 4622 21732 4646 21734
rect 4406 21712 4702 21732
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4406 20700 4702 20720
rect 4462 20698 4486 20700
rect 4542 20698 4566 20700
rect 4622 20698 4646 20700
rect 4484 20646 4486 20698
rect 4548 20646 4560 20698
rect 4622 20646 4624 20698
rect 4462 20644 4486 20646
rect 4542 20644 4566 20646
rect 4622 20644 4646 20646
rect 4406 20624 4702 20644
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 4172 20058 4200 20198
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 3700 19916 3752 19922
rect 3700 19858 3752 19864
rect 2504 18284 2556 18290
rect 2504 18226 2556 18232
rect 3712 17746 3740 19858
rect 4406 19612 4702 19632
rect 4462 19610 4486 19612
rect 4542 19610 4566 19612
rect 4622 19610 4646 19612
rect 4484 19558 4486 19610
rect 4548 19558 4560 19610
rect 4622 19558 4624 19610
rect 4462 19556 4486 19558
rect 4542 19556 4566 19558
rect 4622 19556 4646 19558
rect 4406 19536 4702 19556
rect 4406 18524 4702 18544
rect 4462 18522 4486 18524
rect 4542 18522 4566 18524
rect 4622 18522 4646 18524
rect 4484 18470 4486 18522
rect 4548 18470 4560 18522
rect 4622 18470 4624 18522
rect 4462 18468 4486 18470
rect 4542 18468 4566 18470
rect 4622 18468 4646 18470
rect 4406 18448 4702 18468
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 3976 18148 4028 18154
rect 3976 18090 4028 18096
rect 3988 17882 4016 18090
rect 4632 17882 4660 18226
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 3700 17740 3752 17746
rect 3700 17682 3752 17688
rect 4406 17436 4702 17456
rect 4462 17434 4486 17436
rect 4542 17434 4566 17436
rect 4622 17434 4646 17436
rect 4484 17382 4486 17434
rect 4548 17382 4560 17434
rect 4622 17382 4624 17434
rect 4462 17380 4486 17382
rect 4542 17380 4566 17382
rect 4622 17380 4646 17382
rect 4406 17360 4702 17380
rect 4406 16348 4702 16368
rect 4462 16346 4486 16348
rect 4542 16346 4566 16348
rect 4622 16346 4646 16348
rect 4484 16294 4486 16346
rect 4548 16294 4560 16346
rect 4622 16294 4624 16346
rect 4462 16292 4486 16294
rect 4542 16292 4566 16294
rect 4622 16292 4646 16294
rect 4406 16272 4702 16292
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 2700 15434 2728 15914
rect 2688 15428 2740 15434
rect 2688 15370 2740 15376
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1964 14074 1992 14758
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2148 12782 2176 13126
rect 2136 12776 2188 12782
rect 2136 12718 2188 12724
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1584 9104 1636 9110
rect 1584 9046 1636 9052
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 8265 1440 8366
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1688 6662 1716 10066
rect 1780 8838 1808 11086
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2424 9586 2452 11018
rect 2700 10606 2728 15370
rect 2884 14958 2912 15982
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 3252 14822 3280 15506
rect 4406 15260 4702 15280
rect 4462 15258 4486 15260
rect 4542 15258 4566 15260
rect 4622 15258 4646 15260
rect 4484 15206 4486 15258
rect 4548 15206 4560 15258
rect 4622 15206 4624 15258
rect 4462 15204 4486 15206
rect 4542 15204 4566 15206
rect 4622 15204 4646 15206
rect 4406 15184 4702 15204
rect 3332 14884 3384 14890
rect 3332 14826 3384 14832
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 3344 13530 3372 14826
rect 4406 14172 4702 14192
rect 4462 14170 4486 14172
rect 4542 14170 4566 14172
rect 4622 14170 4646 14172
rect 4484 14118 4486 14170
rect 4548 14118 4560 14170
rect 4622 14118 4624 14170
rect 4462 14116 4486 14118
rect 4542 14116 4566 14118
rect 4622 14116 4646 14118
rect 4406 14096 4702 14116
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 3160 12986 3188 13330
rect 4816 13258 4844 22374
rect 4908 22094 4936 22646
rect 6012 22574 6040 24323
rect 7852 22574 7880 24323
rect 9692 22574 9720 24323
rect 11532 23474 11560 24323
rect 11532 23446 11744 23474
rect 11306 22876 11602 22896
rect 11362 22874 11386 22876
rect 11442 22874 11466 22876
rect 11522 22874 11546 22876
rect 11384 22822 11386 22874
rect 11448 22822 11460 22874
rect 11522 22822 11524 22874
rect 11362 22820 11386 22822
rect 11442 22820 11466 22822
rect 11522 22820 11546 22822
rect 11306 22800 11602 22820
rect 11716 22574 11744 23446
rect 11796 22704 11848 22710
rect 11796 22646 11848 22652
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 7840 22568 7892 22574
rect 7840 22510 7892 22516
rect 9680 22568 9732 22574
rect 9680 22510 9732 22516
rect 11704 22568 11756 22574
rect 11704 22510 11756 22516
rect 6368 22432 6420 22438
rect 6368 22374 6420 22380
rect 9680 22432 9732 22438
rect 9680 22374 9732 22380
rect 11152 22432 11204 22438
rect 11152 22374 11204 22380
rect 4908 22066 5120 22094
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 5000 19786 5028 21830
rect 4896 19780 4948 19786
rect 4896 19722 4948 19728
rect 4988 19780 5040 19786
rect 4988 19722 5040 19728
rect 4908 19446 4936 19722
rect 4896 19440 4948 19446
rect 4896 19382 4948 19388
rect 5000 17814 5028 19722
rect 4988 17808 5040 17814
rect 4988 17750 5040 17756
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4908 14550 4936 14758
rect 4896 14544 4948 14550
rect 4896 14486 4948 14492
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4804 13252 4856 13258
rect 4804 13194 4856 13200
rect 4406 13084 4702 13104
rect 4462 13082 4486 13084
rect 4542 13082 4566 13084
rect 4622 13082 4646 13084
rect 4484 13030 4486 13082
rect 4548 13030 4560 13082
rect 4622 13030 4624 13082
rect 4462 13028 4486 13030
rect 4542 13028 4566 13030
rect 4622 13028 4646 13030
rect 4406 13008 4702 13028
rect 4908 12986 4936 13262
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 2976 11218 3004 12718
rect 3240 12708 3292 12714
rect 3240 12650 3292 12656
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2872 10532 2924 10538
rect 2872 10474 2924 10480
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2884 9518 2912 10474
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2228 9444 2280 9450
rect 2228 9386 2280 9392
rect 2240 9178 2268 9386
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2148 7954 2176 8570
rect 2608 7954 2636 9454
rect 2734 9376 2786 9382
rect 2700 9324 2734 9330
rect 2700 9318 2786 9324
rect 2700 9302 2774 9318
rect 2700 9178 2728 9302
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2700 8498 2728 8774
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 2596 7948 2648 7954
rect 2596 7890 2648 7896
rect 2976 7478 3004 11154
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2792 5778 2820 6054
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 1492 5568 1544 5574
rect 1490 5536 1492 5545
rect 2688 5568 2740 5574
rect 1544 5536 1546 5545
rect 2688 5510 2740 5516
rect 1490 5471 1546 5480
rect 2700 5166 2728 5510
rect 3252 5234 3280 12650
rect 3344 12374 3372 12718
rect 3332 12368 3384 12374
rect 3332 12310 3384 12316
rect 4804 12368 4856 12374
rect 4804 12310 4856 12316
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3528 11354 3556 12242
rect 4406 11996 4702 12016
rect 4462 11994 4486 11996
rect 4542 11994 4566 11996
rect 4622 11994 4646 11996
rect 4484 11942 4486 11994
rect 4548 11942 4560 11994
rect 4622 11942 4624 11994
rect 4462 11940 4486 11942
rect 4542 11940 4566 11942
rect 4622 11940 4646 11942
rect 4406 11920 4702 11940
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 4172 10810 4200 11018
rect 4406 10908 4702 10928
rect 4462 10906 4486 10908
rect 4542 10906 4566 10908
rect 4622 10906 4646 10908
rect 4484 10854 4486 10906
rect 4548 10854 4560 10906
rect 4622 10854 4624 10906
rect 4462 10852 4486 10854
rect 4542 10852 4566 10854
rect 4622 10852 4646 10854
rect 4406 10832 4702 10852
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4816 10606 4844 12310
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4406 9820 4702 9840
rect 4462 9818 4486 9820
rect 4542 9818 4566 9820
rect 4622 9818 4646 9820
rect 4484 9766 4486 9818
rect 4548 9766 4560 9818
rect 4622 9766 4624 9818
rect 4462 9764 4486 9766
rect 4542 9764 4566 9766
rect 4622 9764 4646 9766
rect 4406 9744 4702 9764
rect 5000 9518 5028 11494
rect 5092 10266 5120 22066
rect 5264 22092 5316 22098
rect 5264 22034 5316 22040
rect 5540 22092 5592 22098
rect 5540 22034 5592 22040
rect 5172 20256 5224 20262
rect 5172 20198 5224 20204
rect 5184 20058 5212 20198
rect 5172 20052 5224 20058
rect 5172 19994 5224 20000
rect 5184 19922 5212 19994
rect 5172 19916 5224 19922
rect 5172 19858 5224 19864
rect 5184 19310 5212 19858
rect 5276 19786 5304 22034
rect 5448 21888 5500 21894
rect 5448 21830 5500 21836
rect 5460 21418 5488 21830
rect 5552 21690 5580 22034
rect 5816 22024 5868 22030
rect 5816 21966 5868 21972
rect 5828 21690 5856 21966
rect 5540 21684 5592 21690
rect 5540 21626 5592 21632
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5448 21412 5500 21418
rect 5448 21354 5500 21360
rect 5552 20398 5580 21626
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 5264 19780 5316 19786
rect 5264 19722 5316 19728
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5184 17746 5212 18022
rect 5276 17746 5304 19722
rect 5368 19446 5396 20198
rect 5460 19922 5488 20198
rect 5552 19922 5580 20334
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5460 19514 5488 19858
rect 5724 19712 5776 19718
rect 5724 19654 5776 19660
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5356 19440 5408 19446
rect 5356 19382 5408 19388
rect 5736 19310 5764 19654
rect 5632 19304 5684 19310
rect 5632 19246 5684 19252
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 5644 18630 5672 19246
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5632 18624 5684 18630
rect 5632 18566 5684 18572
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 5184 17134 5212 17682
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 5184 13870 5212 17070
rect 5276 16046 5304 17682
rect 5644 17134 5672 18566
rect 5828 17814 5856 19110
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 5816 17808 5868 17814
rect 5816 17750 5868 17756
rect 5724 17740 5776 17746
rect 5724 17682 5776 17688
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 5644 15366 5672 17070
rect 5736 17066 5764 17682
rect 5908 17264 5960 17270
rect 5908 17206 5960 17212
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 5724 17060 5776 17066
rect 5724 17002 5776 17008
rect 5828 16658 5856 17070
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5276 14618 5304 14894
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5644 14550 5672 14758
rect 5632 14544 5684 14550
rect 5632 14486 5684 14492
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5276 12986 5304 14214
rect 5828 14006 5856 16594
rect 5920 16522 5948 17206
rect 6012 16658 6040 17818
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6288 17066 6316 17682
rect 6276 17060 6328 17066
rect 6276 17002 6328 17008
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 5908 16516 5960 16522
rect 5908 16458 5960 16464
rect 5816 14000 5868 14006
rect 5816 13942 5868 13948
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 5184 12442 5212 12718
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 5184 10062 5212 12242
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 5184 9450 5212 9998
rect 4620 9444 4672 9450
rect 4620 9386 4672 9392
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 4632 8906 4660 9386
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3528 8498 3556 8774
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3620 8430 3648 8774
rect 4406 8732 4702 8752
rect 4462 8730 4486 8732
rect 4542 8730 4566 8732
rect 4622 8730 4646 8732
rect 4484 8678 4486 8730
rect 4548 8678 4560 8730
rect 4622 8678 4624 8730
rect 4462 8676 4486 8678
rect 4542 8676 4566 8678
rect 4622 8676 4646 8678
rect 4406 8656 4702 8676
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 3988 7750 4016 8298
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 3896 6798 3924 7210
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3896 6254 3924 6734
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1412 2825 1440 2926
rect 1398 2816 1454 2825
rect 1398 2751 1454 2760
rect 2056 2582 2084 5102
rect 3988 3670 4016 7686
rect 4406 7644 4702 7664
rect 4462 7642 4486 7644
rect 4542 7642 4566 7644
rect 4622 7642 4646 7644
rect 4484 7590 4486 7642
rect 4548 7590 4560 7642
rect 4622 7590 4624 7642
rect 4462 7588 4486 7590
rect 4542 7588 4566 7590
rect 4622 7588 4646 7590
rect 4406 7568 4702 7588
rect 4406 6556 4702 6576
rect 4462 6554 4486 6556
rect 4542 6554 4566 6556
rect 4622 6554 4646 6556
rect 4484 6502 4486 6554
rect 4548 6502 4560 6554
rect 4622 6502 4624 6554
rect 4462 6500 4486 6502
rect 4542 6500 4566 6502
rect 4622 6500 4646 6502
rect 4406 6480 4702 6500
rect 4406 5468 4702 5488
rect 4462 5466 4486 5468
rect 4542 5466 4566 5468
rect 4622 5466 4646 5468
rect 4484 5414 4486 5466
rect 4548 5414 4560 5466
rect 4622 5414 4624 5466
rect 4462 5412 4486 5414
rect 4542 5412 4566 5414
rect 4622 5412 4646 5414
rect 4406 5392 4702 5412
rect 4406 4380 4702 4400
rect 4462 4378 4486 4380
rect 4542 4378 4566 4380
rect 4622 4378 4646 4380
rect 4484 4326 4486 4378
rect 4548 4326 4560 4378
rect 4622 4326 4624 4378
rect 4462 4324 4486 4326
rect 4542 4324 4566 4326
rect 4622 4324 4646 4326
rect 4406 4304 4702 4324
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 4406 3292 4702 3312
rect 4462 3290 4486 3292
rect 4542 3290 4566 3292
rect 4622 3290 4646 3292
rect 4484 3238 4486 3290
rect 4548 3238 4560 3290
rect 4622 3238 4624 3290
rect 4462 3236 4486 3238
rect 4542 3236 4566 3238
rect 4622 3236 4646 3238
rect 4406 3216 4702 3236
rect 4816 2650 4844 9318
rect 5184 8430 5212 9386
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 5276 6798 5304 12038
rect 5368 10810 5396 12786
rect 5552 12442 5580 13398
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6196 12714 6224 12922
rect 6184 12708 6236 12714
rect 6184 12650 6236 12656
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 5828 11762 5856 12242
rect 6196 12238 6224 12650
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 6196 11694 6224 12174
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5368 9042 5396 10746
rect 5736 10538 5764 11630
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5460 10198 5488 10406
rect 6380 10266 6408 22374
rect 7856 22332 8152 22352
rect 7912 22330 7936 22332
rect 7992 22330 8016 22332
rect 8072 22330 8096 22332
rect 7934 22278 7936 22330
rect 7998 22278 8010 22330
rect 8072 22278 8074 22330
rect 7912 22276 7936 22278
rect 7992 22276 8016 22278
rect 8072 22276 8096 22278
rect 7856 22256 8152 22276
rect 7656 21888 7708 21894
rect 7656 21830 7708 21836
rect 7668 21418 7696 21830
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 7196 21412 7248 21418
rect 7196 21354 7248 21360
rect 7656 21412 7708 21418
rect 7656 21354 7708 21360
rect 7208 21146 7236 21354
rect 9048 21350 9076 21490
rect 7748 21344 7800 21350
rect 7748 21286 7800 21292
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 7196 21140 7248 21146
rect 7196 21082 7248 21088
rect 7760 21078 7788 21286
rect 7856 21244 8152 21264
rect 7912 21242 7936 21244
rect 7992 21242 8016 21244
rect 8072 21242 8096 21244
rect 7934 21190 7936 21242
rect 7998 21190 8010 21242
rect 8072 21190 8074 21242
rect 7912 21188 7936 21190
rect 7992 21188 8016 21190
rect 8072 21188 8096 21190
rect 7856 21168 8152 21188
rect 8300 21140 8352 21146
rect 8300 21082 8352 21088
rect 7472 21072 7524 21078
rect 7748 21072 7800 21078
rect 7472 21014 7524 21020
rect 7668 21032 7748 21060
rect 7380 21004 7432 21010
rect 7380 20946 7432 20952
rect 7392 19990 7420 20946
rect 7484 20058 7512 21014
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7380 19984 7432 19990
rect 7380 19926 7432 19932
rect 6460 19440 6512 19446
rect 6460 19382 6512 19388
rect 6472 19310 6500 19382
rect 7484 19378 7512 19994
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 6460 19304 6512 19310
rect 7564 19304 7616 19310
rect 6460 19246 6512 19252
rect 7562 19272 7564 19281
rect 7616 19272 7618 19281
rect 6472 18834 6500 19246
rect 7668 19242 7696 21032
rect 7748 21014 7800 21020
rect 8312 20806 8340 21082
rect 8852 21004 8904 21010
rect 8852 20946 8904 20952
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 7856 20156 8152 20176
rect 7912 20154 7936 20156
rect 7992 20154 8016 20156
rect 8072 20154 8096 20156
rect 7934 20102 7936 20154
rect 7998 20102 8010 20154
rect 8072 20102 8074 20154
rect 7912 20100 7936 20102
rect 7992 20100 8016 20102
rect 8072 20100 8096 20102
rect 7856 20080 8152 20100
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 8208 19916 8260 19922
rect 8208 19858 8260 19864
rect 7760 19514 7788 19858
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7562 19207 7618 19216
rect 7656 19236 7708 19242
rect 7656 19178 7708 19184
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 6460 18828 6512 18834
rect 6460 18770 6512 18776
rect 6472 17134 6500 18770
rect 7576 18630 7604 19110
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 6644 17604 6696 17610
rect 6644 17546 6696 17552
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6552 16448 6604 16454
rect 6552 16390 6604 16396
rect 6564 16046 6592 16390
rect 6656 16182 6684 17546
rect 6748 17202 6776 17614
rect 7380 17264 7432 17270
rect 7380 17206 7432 17212
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6644 16176 6696 16182
rect 6644 16118 6696 16124
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6656 15162 6684 16118
rect 6840 16114 6868 17070
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6840 15162 6868 16050
rect 6932 16046 6960 16594
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6932 15026 6960 15846
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7300 15162 7328 15302
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 7012 14952 7064 14958
rect 7064 14912 7236 14940
rect 7012 14894 7064 14900
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6840 13870 6868 14214
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6472 12782 6500 13806
rect 6656 13394 6684 13806
rect 7208 13802 7236 14912
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6656 12986 6684 13330
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 6472 12170 6500 12718
rect 6748 12442 6776 13670
rect 7208 12714 7236 13738
rect 7196 12708 7248 12714
rect 7196 12650 7248 12656
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6748 12322 6776 12378
rect 6644 12300 6696 12306
rect 6748 12294 6868 12322
rect 6644 12242 6696 12248
rect 6460 12164 6512 12170
rect 6460 12106 6512 12112
rect 6472 10742 6500 12106
rect 6656 11762 6684 12242
rect 6840 11830 6868 12294
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6656 11218 6684 11698
rect 6840 11558 6868 11766
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7208 11218 7236 11290
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 6460 10736 6512 10742
rect 6460 10678 6512 10684
rect 6656 10606 6684 11154
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5552 6254 5580 6802
rect 5920 6254 5948 9862
rect 6656 8498 6684 10542
rect 6748 9178 6776 10610
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6840 10130 6868 10542
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 7300 9586 7328 14554
rect 7392 13530 7420 17206
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7392 11218 7420 13466
rect 7484 12714 7512 14010
rect 7576 13870 7604 14894
rect 7668 14600 7696 19178
rect 7760 17746 7788 19450
rect 7856 19068 8152 19088
rect 7912 19066 7936 19068
rect 7992 19066 8016 19068
rect 8072 19066 8096 19068
rect 7934 19014 7936 19066
rect 7998 19014 8010 19066
rect 8072 19014 8074 19066
rect 7912 19012 7936 19014
rect 7992 19012 8016 19014
rect 8072 19012 8096 19014
rect 7856 18992 8152 19012
rect 7856 17980 8152 18000
rect 7912 17978 7936 17980
rect 7992 17978 8016 17980
rect 8072 17978 8096 17980
rect 7934 17926 7936 17978
rect 7998 17926 8010 17978
rect 8072 17926 8074 17978
rect 7912 17924 7936 17926
rect 7992 17924 8016 17926
rect 8072 17924 8096 17926
rect 7856 17904 8152 17924
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 8220 17678 8248 19858
rect 8864 19786 8892 20946
rect 9048 20466 9076 21286
rect 9312 20800 9364 20806
rect 9312 20742 9364 20748
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 8852 19780 8904 19786
rect 8852 19722 8904 19728
rect 8760 19372 8812 19378
rect 8760 19314 8812 19320
rect 8300 19304 8352 19310
rect 8298 19272 8300 19281
rect 8352 19272 8354 19281
rect 8298 19207 8354 19216
rect 8574 19272 8630 19281
rect 8574 19207 8630 19216
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8496 18426 8524 18702
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 8220 17338 8248 17614
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 7856 16892 8152 16912
rect 7912 16890 7936 16892
rect 7992 16890 8016 16892
rect 8072 16890 8096 16892
rect 7934 16838 7936 16890
rect 7998 16838 8010 16890
rect 8072 16838 8074 16890
rect 7912 16836 7936 16838
rect 7992 16836 8016 16838
rect 8072 16836 8096 16838
rect 7856 16816 8152 16836
rect 7856 15804 8152 15824
rect 7912 15802 7936 15804
rect 7992 15802 8016 15804
rect 8072 15802 8096 15804
rect 7934 15750 7936 15802
rect 7998 15750 8010 15802
rect 8072 15750 8074 15802
rect 7912 15748 7936 15750
rect 7992 15748 8016 15750
rect 8072 15748 8096 15750
rect 7856 15728 8152 15748
rect 7856 14716 8152 14736
rect 7912 14714 7936 14716
rect 7992 14714 8016 14716
rect 8072 14714 8096 14716
rect 7934 14662 7936 14714
rect 7998 14662 8010 14714
rect 8072 14662 8074 14714
rect 7912 14660 7936 14662
rect 7992 14660 8016 14662
rect 8072 14660 8096 14662
rect 7856 14640 8152 14660
rect 7668 14572 8064 14600
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7484 12374 7512 12650
rect 7472 12368 7524 12374
rect 7472 12310 7524 12316
rect 7576 11354 7604 13806
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7668 12714 7696 13670
rect 7760 12782 7788 14214
rect 8036 14074 8064 14572
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8036 13870 8064 14010
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 8036 13716 8064 13806
rect 8208 13728 8260 13734
rect 8036 13688 8208 13716
rect 8208 13670 8260 13676
rect 7856 13628 8152 13648
rect 7912 13626 7936 13628
rect 7992 13626 8016 13628
rect 8072 13626 8096 13628
rect 7934 13574 7936 13626
rect 7998 13574 8010 13626
rect 8072 13574 8074 13626
rect 7912 13572 7936 13574
rect 7992 13572 8016 13574
rect 8072 13572 8096 13574
rect 7856 13552 8152 13572
rect 8312 13530 8340 17614
rect 8496 17610 8524 18362
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8404 16726 8432 17478
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8404 15910 8432 16662
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8496 15026 8524 15506
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8496 13818 8524 14418
rect 8588 14074 8616 19207
rect 8772 18272 8800 19314
rect 8864 18834 8892 19722
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 8864 18698 8892 18770
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8956 18426 8984 18566
rect 8944 18420 8996 18426
rect 8944 18362 8996 18368
rect 8772 18244 8892 18272
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8760 18080 8812 18086
rect 8864 18068 8892 18244
rect 8812 18040 8892 18068
rect 8760 18022 8812 18028
rect 8680 17542 8708 18022
rect 8772 17746 8800 18022
rect 9048 17746 9076 20402
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9232 18834 9260 19110
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9324 18222 9352 20742
rect 9588 19304 9640 19310
rect 9588 19246 9640 19252
rect 9600 18834 9628 19246
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9416 18290 9444 18566
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 8760 17740 8812 17746
rect 8760 17682 8812 17688
rect 9036 17740 9088 17746
rect 9036 17682 9088 17688
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8680 14278 8708 17478
rect 8772 15638 8800 17682
rect 8852 16652 8904 16658
rect 8852 16594 8904 16600
rect 8864 16046 8892 16594
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 8944 16040 8996 16046
rect 8944 15982 8996 15988
rect 8956 15706 8984 15982
rect 9048 15706 9076 17682
rect 9140 17338 9168 18158
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9324 16182 9352 18158
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9600 17814 9628 18022
rect 9588 17808 9640 17814
rect 9588 17750 9640 17756
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9312 16176 9364 16182
rect 9312 16118 9364 16124
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 9048 14482 9076 15642
rect 9140 15502 9168 15846
rect 9324 15502 9352 16118
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8576 14068 8628 14074
rect 8628 14028 8708 14056
rect 8576 14010 8628 14016
rect 8496 13790 8616 13818
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 8128 12850 8156 13330
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8312 12782 8340 13466
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 7760 11830 7788 12718
rect 7856 12540 8152 12560
rect 7912 12538 7936 12540
rect 7992 12538 8016 12540
rect 8072 12538 8096 12540
rect 7934 12486 7936 12538
rect 7998 12486 8010 12538
rect 8072 12486 8074 12538
rect 7912 12484 7936 12486
rect 7992 12484 8016 12486
rect 8072 12484 8096 12486
rect 7856 12464 8152 12484
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 8496 11762 8524 12718
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7760 11218 7788 11630
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 7856 11452 8152 11472
rect 7912 11450 7936 11452
rect 7992 11450 8016 11452
rect 8072 11450 8096 11452
rect 7934 11398 7936 11450
rect 7998 11398 8010 11450
rect 8072 11398 8074 11450
rect 7912 11396 7936 11398
rect 7992 11396 8016 11398
rect 8072 11396 8096 11398
rect 7856 11376 8152 11396
rect 8220 11286 8248 11494
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 8116 11144 8168 11150
rect 8220 11098 8248 11222
rect 8168 11092 8248 11098
rect 8116 11086 8248 11092
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7564 11076 7616 11082
rect 8128 11070 8248 11086
rect 7564 11018 7616 11024
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 6196 6186 6224 6802
rect 6184 6180 6236 6186
rect 6184 6122 6236 6128
rect 4988 5840 5040 5846
rect 4988 5782 5040 5788
rect 5000 4690 5028 5782
rect 6276 5092 6328 5098
rect 6276 5034 6328 5040
rect 6288 4758 6316 5034
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 6656 2650 6684 8298
rect 6748 3602 6776 8978
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6932 5914 6960 6190
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 7024 5370 7052 5714
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 7024 5030 7052 5102
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6840 3602 6868 4694
rect 7024 4690 7052 4966
rect 7392 4758 7420 11018
rect 7380 4752 7432 4758
rect 7380 4694 7432 4700
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7116 4282 7144 4490
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7576 3942 7604 11018
rect 8220 10606 8248 11070
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 7856 10364 8152 10384
rect 7912 10362 7936 10364
rect 7992 10362 8016 10364
rect 8072 10362 8096 10364
rect 7934 10310 7936 10362
rect 7998 10310 8010 10362
rect 8072 10310 8074 10362
rect 7912 10308 7936 10310
rect 7992 10308 8016 10310
rect 8072 10308 8096 10310
rect 7856 10288 8152 10308
rect 7856 9276 8152 9296
rect 7912 9274 7936 9276
rect 7992 9274 8016 9276
rect 8072 9274 8096 9276
rect 7934 9222 7936 9274
rect 7998 9222 8010 9274
rect 8072 9222 8074 9274
rect 7912 9220 7936 9222
rect 7992 9220 8016 9222
rect 8072 9220 8096 9222
rect 7856 9200 8152 9220
rect 8312 8906 8340 10950
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8404 8974 8432 9386
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 7856 8188 8152 8208
rect 7912 8186 7936 8188
rect 7992 8186 8016 8188
rect 8072 8186 8096 8188
rect 7934 8134 7936 8186
rect 7998 8134 8010 8186
rect 8072 8134 8074 8186
rect 7912 8132 7936 8134
rect 7992 8132 8016 8134
rect 8072 8132 8096 8134
rect 7856 8112 8152 8132
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7668 7546 7696 7890
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7856 7100 8152 7120
rect 7912 7098 7936 7100
rect 7992 7098 8016 7100
rect 8072 7098 8096 7100
rect 7934 7046 7936 7098
rect 7998 7046 8010 7098
rect 8072 7046 8074 7098
rect 7912 7044 7936 7046
rect 7992 7044 8016 7046
rect 8072 7044 8096 7046
rect 7856 7024 8152 7044
rect 8312 7002 8340 8842
rect 8404 8430 8432 8910
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8404 8022 8432 8366
rect 8588 8090 8616 13790
rect 8680 12986 8708 14028
rect 9508 13870 9536 17274
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9600 15094 9628 15506
rect 9588 15088 9640 15094
rect 9588 15030 9640 15036
rect 9600 13938 9628 15030
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8680 11694 8708 12922
rect 9508 12850 9536 13806
rect 9600 12918 9628 13874
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8680 11218 8708 11630
rect 9140 11558 9168 12582
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 9140 10606 9168 11494
rect 9508 10606 9536 12650
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8588 7410 8616 7890
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 8588 7002 8616 7346
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 7856 6012 8152 6032
rect 7912 6010 7936 6012
rect 7992 6010 8016 6012
rect 8072 6010 8096 6012
rect 7934 5958 7936 6010
rect 7998 5958 8010 6010
rect 8072 5958 8074 6010
rect 7912 5956 7936 5958
rect 7992 5956 8016 5958
rect 8072 5956 8096 5958
rect 7856 5936 8152 5956
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7760 4826 7788 5170
rect 7856 4924 8152 4944
rect 7912 4922 7936 4924
rect 7992 4922 8016 4924
rect 8072 4922 8096 4924
rect 7934 4870 7936 4922
rect 7998 4870 8010 4922
rect 8072 4870 8074 4922
rect 7912 4868 7936 4870
rect 7992 4868 8016 4870
rect 8072 4868 8096 4870
rect 7856 4848 8152 4868
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 8496 4622 8524 6802
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7856 3836 8152 3856
rect 7912 3834 7936 3836
rect 7992 3834 8016 3836
rect 8072 3834 8096 3836
rect 7934 3782 7936 3834
rect 7998 3782 8010 3834
rect 8072 3782 8074 3834
rect 7912 3780 7936 3782
rect 7992 3780 8016 3782
rect 8072 3780 8096 3782
rect 7856 3760 8152 3780
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6748 2650 6776 3538
rect 7856 2748 8152 2768
rect 7912 2746 7936 2748
rect 7992 2746 8016 2748
rect 8072 2746 8096 2748
rect 7934 2694 7936 2746
rect 7998 2694 8010 2746
rect 8072 2694 8074 2746
rect 7912 2692 7936 2694
rect 7992 2692 8016 2694
rect 8072 2692 8096 2694
rect 7856 2672 8152 2692
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 8220 2582 8248 4490
rect 8496 3058 8524 4558
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8956 2990 8984 10406
rect 9140 10198 9168 10542
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9128 10192 9180 10198
rect 9128 10134 9180 10140
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9232 9586 9260 9998
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9600 9518 9628 10406
rect 9692 9586 9720 22374
rect 10324 22092 10376 22098
rect 10324 22034 10376 22040
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 10060 21418 10088 21830
rect 10048 21412 10100 21418
rect 10048 21354 10100 21360
rect 10336 19922 10364 22034
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 11072 20466 11100 20742
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 10508 20324 10560 20330
rect 10508 20266 10560 20272
rect 10520 20058 10548 20266
rect 10508 20052 10560 20058
rect 10508 19994 10560 20000
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 10336 18222 10364 19858
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10612 17814 10640 18022
rect 10600 17808 10652 17814
rect 10600 17750 10652 17756
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10152 17134 10180 17478
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10980 16046 11008 18158
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 9864 15428 9916 15434
rect 9864 15370 9916 15376
rect 9876 14958 9904 15370
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9772 14884 9824 14890
rect 9772 14826 9824 14832
rect 9784 14074 9812 14826
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9876 12986 9904 13670
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 10060 12986 10088 13262
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10060 11762 10088 12922
rect 10152 12782 10180 13806
rect 10888 13258 10916 15302
rect 10980 14618 11008 15982
rect 11164 14890 11192 22374
rect 11704 22092 11756 22098
rect 11704 22034 11756 22040
rect 11306 21788 11602 21808
rect 11362 21786 11386 21788
rect 11442 21786 11466 21788
rect 11522 21786 11546 21788
rect 11384 21734 11386 21786
rect 11448 21734 11460 21786
rect 11522 21734 11524 21786
rect 11362 21732 11386 21734
rect 11442 21732 11466 21734
rect 11522 21732 11546 21734
rect 11306 21712 11602 21732
rect 11244 21412 11296 21418
rect 11244 21354 11296 21360
rect 11256 21010 11284 21354
rect 11716 21010 11744 22034
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 11704 21004 11756 21010
rect 11704 20946 11756 20952
rect 11306 20700 11602 20720
rect 11362 20698 11386 20700
rect 11442 20698 11466 20700
rect 11522 20698 11546 20700
rect 11384 20646 11386 20698
rect 11448 20646 11460 20698
rect 11522 20646 11524 20698
rect 11362 20644 11386 20646
rect 11442 20644 11466 20646
rect 11522 20644 11546 20646
rect 11306 20624 11602 20644
rect 11306 19612 11602 19632
rect 11362 19610 11386 19612
rect 11442 19610 11466 19612
rect 11522 19610 11546 19612
rect 11384 19558 11386 19610
rect 11448 19558 11460 19610
rect 11522 19558 11524 19610
rect 11362 19556 11386 19558
rect 11442 19556 11466 19558
rect 11522 19556 11546 19558
rect 11306 19536 11602 19556
rect 11306 18524 11602 18544
rect 11362 18522 11386 18524
rect 11442 18522 11466 18524
rect 11522 18522 11546 18524
rect 11384 18470 11386 18522
rect 11448 18470 11460 18522
rect 11522 18470 11524 18522
rect 11362 18468 11386 18470
rect 11442 18468 11466 18470
rect 11522 18468 11546 18470
rect 11306 18448 11602 18468
rect 11808 17746 11836 22646
rect 12912 22574 12940 24323
rect 14752 22574 14780 24323
rect 16592 22574 16620 24323
rect 17972 22574 18000 24323
rect 18206 22876 18502 22896
rect 18262 22874 18286 22876
rect 18342 22874 18366 22876
rect 18422 22874 18446 22876
rect 18284 22822 18286 22874
rect 18348 22822 18360 22874
rect 18422 22822 18424 22874
rect 18262 22820 18286 22822
rect 18342 22820 18366 22822
rect 18422 22820 18446 22822
rect 18206 22800 18502 22820
rect 19812 22574 19840 24323
rect 21086 23216 21142 23225
rect 21086 23151 21142 23160
rect 21100 22574 21128 23151
rect 21652 22574 21680 24323
rect 12900 22568 12952 22574
rect 12900 22510 12952 22516
rect 14740 22568 14792 22574
rect 14740 22510 14792 22516
rect 16580 22568 16632 22574
rect 16580 22510 16632 22516
rect 17960 22568 18012 22574
rect 17960 22510 18012 22516
rect 19800 22568 19852 22574
rect 19800 22510 19852 22516
rect 21088 22568 21140 22574
rect 21088 22510 21140 22516
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 13084 22432 13136 22438
rect 13084 22374 13136 22380
rect 14556 22432 14608 22438
rect 14556 22374 14608 22380
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 19616 22432 19668 22438
rect 19616 22374 19668 22380
rect 20904 22432 20956 22438
rect 20904 22374 20956 22380
rect 20996 22432 21048 22438
rect 20996 22374 21048 22380
rect 11888 22092 11940 22098
rect 11888 22034 11940 22040
rect 11980 22092 12032 22098
rect 11980 22034 12032 22040
rect 12348 22092 12400 22098
rect 12348 22034 12400 22040
rect 11900 21350 11928 22034
rect 11888 21344 11940 21350
rect 11888 21286 11940 21292
rect 11900 20398 11928 21286
rect 11992 21146 12020 22034
rect 12072 21888 12124 21894
rect 12072 21830 12124 21836
rect 12084 21554 12112 21830
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 11980 21140 12032 21146
rect 11980 21082 12032 21088
rect 12360 21010 12388 22034
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12820 21418 12848 21830
rect 12808 21412 12860 21418
rect 12808 21354 12860 21360
rect 12624 21072 12676 21078
rect 12624 21014 12676 21020
rect 11980 21004 12032 21010
rect 11980 20946 12032 20952
rect 12164 21004 12216 21010
rect 12164 20946 12216 20952
rect 12348 21004 12400 21010
rect 12348 20946 12400 20952
rect 11992 20534 12020 20946
rect 11980 20528 12032 20534
rect 11980 20470 12032 20476
rect 12176 20398 12204 20946
rect 12636 20398 12664 21014
rect 11888 20392 11940 20398
rect 11888 20334 11940 20340
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12544 18834 12572 20334
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12636 18222 12664 19110
rect 12728 18834 12756 19246
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13004 18902 13032 19110
rect 12992 18896 13044 18902
rect 12992 18838 13044 18844
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 11306 17436 11602 17456
rect 11362 17434 11386 17436
rect 11442 17434 11466 17436
rect 11522 17434 11546 17436
rect 11384 17382 11386 17434
rect 11448 17382 11460 17434
rect 11522 17382 11524 17434
rect 11362 17380 11386 17382
rect 11442 17380 11466 17382
rect 11522 17380 11546 17382
rect 11306 17360 11602 17380
rect 12360 17134 12388 17682
rect 12452 17202 12480 17682
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12636 17338 12664 17478
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12636 17202 12664 17274
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 11306 16348 11602 16368
rect 11362 16346 11386 16348
rect 11442 16346 11466 16348
rect 11522 16346 11546 16348
rect 11384 16294 11386 16346
rect 11448 16294 11460 16346
rect 11522 16294 11524 16346
rect 11362 16292 11386 16294
rect 11442 16292 11466 16294
rect 11522 16292 11546 16294
rect 11306 16272 11602 16292
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11256 15638 11284 15846
rect 12176 15706 12204 17070
rect 12164 15700 12216 15706
rect 12164 15642 12216 15648
rect 11244 15632 11296 15638
rect 11244 15574 11296 15580
rect 11306 15260 11602 15280
rect 11362 15258 11386 15260
rect 11442 15258 11466 15260
rect 11522 15258 11546 15260
rect 11384 15206 11386 15258
rect 11448 15206 11460 15258
rect 11522 15206 11524 15258
rect 11362 15204 11386 15206
rect 11442 15204 11466 15206
rect 11522 15204 11546 15206
rect 11306 15184 11602 15204
rect 12452 15162 12480 17138
rect 12728 17134 12756 17546
rect 12820 17270 12848 18702
rect 13004 18358 13032 18838
rect 12992 18352 13044 18358
rect 12992 18294 13044 18300
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 13004 15706 13032 18158
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 11152 14884 11204 14890
rect 11152 14826 11204 14832
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 11306 14172 11602 14192
rect 11362 14170 11386 14172
rect 11442 14170 11466 14172
rect 11522 14170 11546 14172
rect 11384 14118 11386 14170
rect 11448 14118 11460 14170
rect 11522 14118 11524 14170
rect 11362 14116 11386 14118
rect 11442 14116 11466 14118
rect 11522 14116 11546 14118
rect 11306 14096 11602 14116
rect 12084 13462 12112 14962
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10152 11898 10180 12718
rect 10324 12436 10376 12442
rect 10428 12434 10456 13194
rect 10376 12406 10456 12434
rect 10980 12730 11008 13330
rect 11306 13084 11602 13104
rect 11362 13082 11386 13084
rect 11442 13082 11466 13084
rect 11522 13082 11546 13084
rect 11384 13030 11386 13082
rect 11448 13030 11460 13082
rect 11522 13030 11524 13082
rect 11362 13028 11386 13030
rect 11442 13028 11466 13030
rect 11522 13028 11546 13030
rect 11306 13008 11602 13028
rect 12084 12986 12112 13398
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 11244 12912 11296 12918
rect 11244 12854 11296 12860
rect 10980 12714 11100 12730
rect 11256 12714 11284 12854
rect 10980 12708 11112 12714
rect 10980 12702 11060 12708
rect 10324 12378 10376 12384
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10048 11620 10100 11626
rect 10048 11562 10100 11568
rect 10060 11234 10088 11562
rect 10140 11280 10192 11286
rect 10060 11228 10140 11234
rect 10060 11222 10192 11228
rect 10336 11234 10364 12378
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10520 11354 10548 11834
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10060 11206 10180 11222
rect 10336 11218 10456 11234
rect 10336 11212 10468 11218
rect 10336 11206 10416 11212
rect 10060 10674 10088 11206
rect 10416 11154 10468 11160
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9784 10130 9812 10202
rect 10060 10130 10088 10610
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9588 9512 9640 9518
rect 9784 9466 9812 10066
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 9588 9454 9640 9460
rect 9600 8838 9628 9454
rect 9692 9450 9812 9466
rect 9680 9444 9812 9450
rect 9732 9438 9812 9444
rect 9680 9386 9732 9392
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9784 7886 9812 9438
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9416 7410 9444 7686
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9508 7342 9536 7686
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9784 6866 9812 7822
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9692 5234 9720 5578
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 9140 3670 9168 5102
rect 9692 4706 9720 5170
rect 9876 4826 9904 8774
rect 10152 6866 10180 9318
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10244 6934 10272 7890
rect 10232 6928 10284 6934
rect 10232 6870 10284 6876
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10336 5166 10364 9930
rect 10428 9518 10456 11154
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10428 9178 10456 9454
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10428 8498 10456 8978
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10428 7342 10456 8434
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9692 4678 9904 4706
rect 10336 4690 10364 5102
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9128 3664 9180 3670
rect 9128 3606 9180 3612
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9048 3194 9076 3470
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 9508 3058 9536 3674
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 9692 2650 9720 4558
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9784 3194 9812 3402
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9876 2990 9904 4678
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10520 3058 10548 11290
rect 10980 11014 11008 12702
rect 11060 12650 11112 12656
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11348 12374 11376 12582
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11716 12306 11744 12582
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11306 11996 11602 12016
rect 11362 11994 11386 11996
rect 11442 11994 11466 11996
rect 11522 11994 11546 11996
rect 11384 11942 11386 11994
rect 11448 11942 11460 11994
rect 11522 11942 11524 11994
rect 11362 11940 11386 11942
rect 11442 11940 11466 11942
rect 11522 11940 11546 11942
rect 11306 11920 11602 11940
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 10980 9586 11008 10950
rect 11072 10810 11100 11154
rect 11808 11150 11836 12242
rect 12084 11286 12112 12922
rect 12176 12442 12204 13262
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12268 12850 12296 13194
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 12084 11150 12112 11222
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 11306 10908 11602 10928
rect 11362 10906 11386 10908
rect 11442 10906 11466 10908
rect 11522 10906 11546 10908
rect 11384 10854 11386 10906
rect 11448 10854 11460 10906
rect 11522 10854 11524 10906
rect 11362 10852 11386 10854
rect 11442 10852 11466 10854
rect 11522 10852 11546 10854
rect 11306 10832 11602 10852
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 12084 10266 12112 11086
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11306 9820 11602 9840
rect 11362 9818 11386 9820
rect 11442 9818 11466 9820
rect 11522 9818 11546 9820
rect 11384 9766 11386 9818
rect 11448 9766 11460 9818
rect 11522 9766 11524 9818
rect 11362 9764 11386 9766
rect 11442 9764 11466 9766
rect 11522 9764 11546 9766
rect 11306 9744 11602 9764
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10980 9110 11008 9522
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10980 8430 11008 9046
rect 12084 9042 12112 9386
rect 12452 9110 12480 9454
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 11306 8732 11602 8752
rect 11362 8730 11386 8732
rect 11442 8730 11466 8732
rect 11522 8730 11546 8732
rect 11384 8678 11386 8730
rect 11448 8678 11460 8730
rect 11522 8678 11524 8730
rect 11362 8676 11386 8678
rect 11442 8676 11466 8678
rect 11522 8676 11546 8678
rect 11306 8656 11602 8676
rect 12084 8430 12112 8978
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 11306 7644 11602 7664
rect 11362 7642 11386 7644
rect 11442 7642 11466 7644
rect 11522 7642 11546 7644
rect 11384 7590 11386 7642
rect 11448 7590 11460 7642
rect 11522 7590 11524 7642
rect 11362 7588 11386 7590
rect 11442 7588 11466 7590
rect 11522 7588 11546 7590
rect 11306 7568 11602 7588
rect 12360 7410 12388 7686
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10612 6866 10640 7210
rect 12544 6914 12572 15438
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12820 12918 12848 13330
rect 12808 12912 12860 12918
rect 12808 12854 12860 12860
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12912 10674 12940 12582
rect 13096 11286 13124 22374
rect 13544 21344 13596 21350
rect 13544 21286 13596 21292
rect 13556 21078 13584 21286
rect 13544 21072 13596 21078
rect 13544 21014 13596 21020
rect 14568 19938 14596 22374
rect 14756 22332 15052 22352
rect 14812 22330 14836 22332
rect 14892 22330 14916 22332
rect 14972 22330 14996 22332
rect 14834 22278 14836 22330
rect 14898 22278 14910 22330
rect 14972 22278 14974 22330
rect 14812 22276 14836 22278
rect 14892 22276 14916 22278
rect 14972 22276 14996 22278
rect 14756 22256 15052 22276
rect 15476 22228 15528 22234
rect 15476 22170 15528 22176
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 15108 21548 15160 21554
rect 15108 21490 15160 21496
rect 14648 21412 14700 21418
rect 14648 21354 14700 21360
rect 14660 21146 14688 21354
rect 14756 21244 15052 21264
rect 14812 21242 14836 21244
rect 14892 21242 14916 21244
rect 14972 21242 14996 21244
rect 14834 21190 14836 21242
rect 14898 21190 14910 21242
rect 14972 21190 14974 21242
rect 14812 21188 14836 21190
rect 14892 21188 14916 21190
rect 14972 21188 14996 21190
rect 14756 21168 15052 21188
rect 14648 21140 14700 21146
rect 14648 21082 14700 21088
rect 15120 21078 15148 21490
rect 15304 21418 15332 21830
rect 15292 21412 15344 21418
rect 15292 21354 15344 21360
rect 15108 21072 15160 21078
rect 15108 21014 15160 21020
rect 15120 20398 15148 21014
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 15212 20466 15240 20946
rect 15384 20936 15436 20942
rect 15384 20878 15436 20884
rect 15396 20806 15424 20878
rect 15384 20800 15436 20806
rect 15384 20742 15436 20748
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15108 20392 15160 20398
rect 15160 20340 15240 20346
rect 15108 20334 15240 20340
rect 15120 20318 15240 20334
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 14756 20156 15052 20176
rect 14812 20154 14836 20156
rect 14892 20154 14916 20156
rect 14972 20154 14996 20156
rect 14834 20102 14836 20154
rect 14898 20102 14910 20154
rect 14972 20102 14974 20154
rect 14812 20100 14836 20102
rect 14892 20100 14916 20102
rect 14972 20100 14996 20102
rect 14756 20080 15052 20100
rect 14464 19916 14516 19922
rect 14568 19910 14780 19938
rect 15120 19922 15148 20198
rect 15212 19922 15240 20318
rect 15396 19990 15424 20742
rect 15384 19984 15436 19990
rect 15384 19926 15436 19932
rect 14464 19858 14516 19864
rect 14476 19310 14504 19858
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14568 19514 14596 19790
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14660 19378 14688 19654
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14752 19310 14780 19910
rect 15108 19916 15160 19922
rect 15108 19858 15160 19864
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 14924 19848 14976 19854
rect 14924 19790 14976 19796
rect 14936 19310 14964 19790
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 15016 19508 15068 19514
rect 15016 19450 15068 19456
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 14464 19304 14516 19310
rect 14740 19304 14792 19310
rect 14464 19246 14516 19252
rect 14660 19252 14740 19258
rect 14660 19246 14792 19252
rect 14924 19304 14976 19310
rect 14924 19246 14976 19252
rect 15028 19258 15056 19450
rect 13924 19174 13952 19246
rect 14660 19230 14780 19246
rect 15028 19242 15148 19258
rect 15212 19242 15240 19654
rect 15016 19236 15148 19242
rect 14660 19174 14688 19230
rect 15068 19230 15148 19236
rect 15016 19178 15068 19184
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14756 19068 15052 19088
rect 14812 19066 14836 19068
rect 14892 19066 14916 19068
rect 14972 19066 14996 19068
rect 14834 19014 14836 19066
rect 14898 19014 14910 19066
rect 14972 19014 14974 19066
rect 14812 19012 14836 19014
rect 14892 19012 14916 19014
rect 14972 19012 14996 19014
rect 14756 18992 15052 19012
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13188 18290 13216 18566
rect 13372 18358 13400 18770
rect 13360 18352 13412 18358
rect 13360 18294 13412 18300
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13280 17338 13308 18158
rect 14756 17980 15052 18000
rect 14812 17978 14836 17980
rect 14892 17978 14916 17980
rect 14972 17978 14996 17980
rect 14834 17926 14836 17978
rect 14898 17926 14910 17978
rect 14972 17926 14974 17978
rect 14812 17924 14836 17926
rect 14892 17924 14916 17926
rect 14972 17924 14996 17926
rect 14756 17904 15052 17924
rect 13912 17740 13964 17746
rect 13912 17682 13964 17688
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13924 14482 13952 17682
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14752 17202 14780 17478
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14756 16892 15052 16912
rect 14812 16890 14836 16892
rect 14892 16890 14916 16892
rect 14972 16890 14996 16892
rect 14834 16838 14836 16890
rect 14898 16838 14910 16890
rect 14972 16838 14974 16890
rect 14812 16836 14836 16838
rect 14892 16836 14916 16838
rect 14972 16836 14996 16838
rect 14756 16816 15052 16836
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 14556 16176 14608 16182
rect 14556 16118 14608 16124
rect 14568 15570 14596 16118
rect 15028 15994 15056 16594
rect 15120 16250 15148 19230
rect 15200 19236 15252 19242
rect 15200 19178 15252 19184
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15212 16658 15240 17682
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15028 15966 15148 15994
rect 14756 15804 15052 15824
rect 14812 15802 14836 15804
rect 14892 15802 14916 15804
rect 14972 15802 14996 15804
rect 14834 15750 14836 15802
rect 14898 15750 14910 15802
rect 14972 15750 14974 15802
rect 14812 15748 14836 15750
rect 14892 15748 14916 15750
rect 14972 15748 14996 15750
rect 14756 15728 15052 15748
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14568 14618 14596 15506
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14660 14618 14688 14894
rect 14756 14716 15052 14736
rect 14812 14714 14836 14716
rect 14892 14714 14916 14716
rect 14972 14714 14996 14716
rect 14834 14662 14836 14714
rect 14898 14662 14910 14714
rect 14972 14662 14974 14714
rect 14812 14660 14836 14662
rect 14892 14660 14916 14662
rect 14972 14660 14996 14662
rect 14756 14640 15052 14660
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13832 14074 13860 14350
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13924 13394 13952 14418
rect 14660 13462 14688 14554
rect 15120 14074 15148 15966
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15212 15570 15240 15846
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 15200 14884 15252 14890
rect 15200 14826 15252 14832
rect 15212 14482 15240 14826
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15108 14068 15160 14074
rect 15108 14010 15160 14016
rect 14756 13628 15052 13648
rect 14812 13626 14836 13628
rect 14892 13626 14916 13628
rect 14972 13626 14996 13628
rect 14834 13574 14836 13626
rect 14898 13574 14910 13626
rect 14972 13574 14974 13626
rect 14812 13572 14836 13574
rect 14892 13572 14916 13574
rect 14972 13572 14996 13574
rect 14756 13552 15052 13572
rect 14372 13456 14424 13462
rect 14372 13398 14424 13404
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 13280 12782 13308 13126
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12912 10130 12940 10610
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13648 10266 13676 10542
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12820 8090 12848 8298
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12452 6886 12572 6914
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11164 5098 11192 6802
rect 11306 6556 11602 6576
rect 11362 6554 11386 6556
rect 11442 6554 11466 6556
rect 11522 6554 11546 6556
rect 11384 6502 11386 6554
rect 11448 6502 11460 6554
rect 11522 6502 11524 6554
rect 11362 6500 11386 6502
rect 11442 6500 11466 6502
rect 11522 6500 11546 6502
rect 11306 6480 11602 6500
rect 11306 5468 11602 5488
rect 11362 5466 11386 5468
rect 11442 5466 11466 5468
rect 11522 5466 11546 5468
rect 11384 5414 11386 5466
rect 11448 5414 11460 5466
rect 11522 5414 11524 5466
rect 11362 5412 11386 5414
rect 11442 5412 11466 5414
rect 11522 5412 11546 5414
rect 11306 5392 11602 5412
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11888 5092 11940 5098
rect 11888 5034 11940 5040
rect 11164 4758 11192 5034
rect 11152 4752 11204 4758
rect 11152 4694 11204 4700
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11306 4380 11602 4400
rect 11362 4378 11386 4380
rect 11442 4378 11466 4380
rect 11522 4378 11546 4380
rect 11384 4326 11386 4378
rect 11448 4326 11460 4378
rect 11522 4326 11524 4378
rect 11362 4324 11386 4326
rect 11442 4324 11466 4326
rect 11522 4324 11546 4326
rect 11306 4304 11602 4324
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10980 2990 11008 3470
rect 11164 3194 11192 3674
rect 11716 3670 11744 4626
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 11900 3602 11928 5034
rect 12360 4826 12388 5102
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11306 3292 11602 3312
rect 11362 3290 11386 3292
rect 11442 3290 11466 3292
rect 11522 3290 11546 3292
rect 11384 3238 11386 3290
rect 11448 3238 11460 3290
rect 11522 3238 11524 3290
rect 11362 3236 11386 3238
rect 11442 3236 11466 3238
rect 11522 3236 11546 3238
rect 11306 3216 11602 3236
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 11808 2922 11836 3334
rect 11900 2990 11928 3538
rect 11992 3398 12020 3878
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 12452 3194 12480 6886
rect 12728 5846 12756 7482
rect 13372 6914 13400 9862
rect 13464 9518 13492 10066
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13556 9382 13584 10066
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13740 7886 13768 13194
rect 14384 12442 14412 13398
rect 15120 13394 15148 14010
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 14756 12540 15052 12560
rect 14812 12538 14836 12540
rect 14892 12538 14916 12540
rect 14972 12538 14996 12540
rect 14834 12486 14836 12538
rect 14898 12486 14910 12538
rect 14972 12486 14974 12538
rect 14812 12484 14836 12486
rect 14892 12484 14916 12486
rect 14972 12484 14996 12486
rect 14756 12464 15052 12484
rect 14372 12436 14424 12442
rect 14372 12378 14424 12384
rect 15120 12374 15148 12582
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 14756 11452 15052 11472
rect 14812 11450 14836 11452
rect 14892 11450 14916 11452
rect 14972 11450 14996 11452
rect 14834 11398 14836 11450
rect 14898 11398 14910 11450
rect 14972 11398 14974 11450
rect 14812 11396 14836 11398
rect 14892 11396 14916 11398
rect 14972 11396 14996 11398
rect 14756 11376 15052 11396
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13832 10198 13860 10746
rect 14844 10606 14872 11018
rect 15028 10810 15056 11154
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14756 10364 15052 10384
rect 14812 10362 14836 10364
rect 14892 10362 14916 10364
rect 14972 10362 14996 10364
rect 14834 10310 14836 10362
rect 14898 10310 14910 10362
rect 14972 10310 14974 10362
rect 14812 10308 14836 10310
rect 14892 10308 14916 10310
rect 14972 10308 14996 10310
rect 14756 10288 15052 10308
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 14756 9276 15052 9296
rect 14812 9274 14836 9276
rect 14892 9274 14916 9276
rect 14972 9274 14996 9276
rect 14834 9222 14836 9274
rect 14898 9222 14910 9274
rect 14972 9222 14974 9274
rect 14812 9220 14836 9222
rect 14892 9220 14916 9222
rect 14972 9220 14996 9222
rect 14756 9200 15052 9220
rect 15304 8974 15332 11086
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15396 10606 15424 11018
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15488 9178 15516 22170
rect 16580 21684 16632 21690
rect 16580 21626 16632 21632
rect 16592 21554 16620 21626
rect 16580 21548 16632 21554
rect 16580 21490 16632 21496
rect 16592 21078 16620 21490
rect 16580 21072 16632 21078
rect 16580 21014 16632 21020
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 15844 20868 15896 20874
rect 15844 20810 15896 20816
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15764 19718 15792 19994
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15764 19174 15792 19654
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15856 18834 15884 20810
rect 16396 20460 16448 20466
rect 16396 20402 16448 20408
rect 16408 19922 16436 20402
rect 15936 19916 15988 19922
rect 15936 19858 15988 19864
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 15948 19802 15976 19858
rect 15948 19774 16068 19802
rect 16040 18834 16068 19774
rect 16132 18834 16160 19858
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 16120 18828 16172 18834
rect 16120 18770 16172 18776
rect 15856 17882 15884 18770
rect 15844 17876 15896 17882
rect 15844 17818 15896 17824
rect 16040 16658 16068 18770
rect 16132 18426 16160 18770
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16120 18420 16172 18426
rect 16120 18362 16172 18368
rect 16224 18154 16252 18702
rect 16212 18148 16264 18154
rect 16212 18090 16264 18096
rect 16212 17808 16264 17814
rect 16212 17750 16264 17756
rect 16224 17338 16252 17750
rect 16408 17746 16436 19858
rect 16500 19786 16528 20878
rect 16488 19780 16540 19786
rect 16488 19722 16540 19728
rect 16486 18864 16542 18873
rect 16542 18808 16620 18816
rect 16486 18799 16488 18808
rect 16540 18788 16620 18808
rect 16488 18770 16540 18776
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 16500 18086 16528 18566
rect 16592 18222 16620 18788
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16592 17678 16620 18158
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 16224 16114 16252 17274
rect 16592 16794 16620 17614
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15580 14482 15608 14758
rect 15764 14482 15792 14758
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15580 14278 15608 14418
rect 15568 14272 15620 14278
rect 15568 14214 15620 14220
rect 15580 13326 15608 14214
rect 16672 13456 16724 13462
rect 16672 13398 16724 13404
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15856 12374 15884 13126
rect 16684 12986 16712 13398
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 16776 12918 16804 22374
rect 17132 22092 17184 22098
rect 17132 22034 17184 22040
rect 17144 21486 17172 22034
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17132 21480 17184 21486
rect 17132 21422 17184 21428
rect 17144 19310 17172 21422
rect 17224 21344 17276 21350
rect 17224 21286 17276 21292
rect 17236 21078 17264 21286
rect 17224 21072 17276 21078
rect 17224 21014 17276 21020
rect 17788 19922 17816 21490
rect 17972 21418 18000 22374
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18206 21788 18502 21808
rect 18262 21786 18286 21788
rect 18342 21786 18366 21788
rect 18422 21786 18446 21788
rect 18284 21734 18286 21786
rect 18348 21734 18360 21786
rect 18422 21734 18424 21786
rect 18262 21732 18286 21734
rect 18342 21732 18366 21734
rect 18422 21732 18446 21734
rect 18206 21712 18502 21732
rect 18708 21418 18736 21830
rect 17960 21412 18012 21418
rect 17960 21354 18012 21360
rect 18696 21412 18748 21418
rect 18696 21354 18748 21360
rect 18206 20700 18502 20720
rect 18262 20698 18286 20700
rect 18342 20698 18366 20700
rect 18422 20698 18446 20700
rect 18284 20646 18286 20698
rect 18348 20646 18360 20698
rect 18422 20646 18424 20698
rect 18262 20644 18286 20646
rect 18342 20644 18366 20646
rect 18422 20644 18446 20646
rect 18206 20624 18502 20644
rect 17776 19916 17828 19922
rect 17776 19858 17828 19864
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 16856 18148 16908 18154
rect 16856 18090 16908 18096
rect 16868 16726 16896 18090
rect 17144 17066 17172 19246
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 17696 18902 17724 19110
rect 17684 18896 17736 18902
rect 17684 18838 17736 18844
rect 17684 18760 17736 18766
rect 17788 18748 17816 19858
rect 18206 19612 18502 19632
rect 18262 19610 18286 19612
rect 18342 19610 18366 19612
rect 18422 19610 18446 19612
rect 18284 19558 18286 19610
rect 18348 19558 18360 19610
rect 18422 19558 18424 19610
rect 18262 19556 18286 19558
rect 18342 19556 18366 19558
rect 18422 19556 18446 19558
rect 18206 19536 18502 19556
rect 18418 18864 18474 18873
rect 19628 18834 19656 22374
rect 20916 22234 20944 22374
rect 20904 22228 20956 22234
rect 20904 22170 20956 22176
rect 21008 22094 21036 22374
rect 20824 22066 21036 22094
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 20180 21418 20208 21830
rect 20168 21412 20220 21418
rect 20168 21354 20220 21360
rect 19708 20324 19760 20330
rect 19708 20266 19760 20272
rect 18418 18799 18474 18808
rect 19156 18828 19208 18834
rect 18432 18766 18460 18799
rect 19156 18770 19208 18776
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19616 18828 19668 18834
rect 19616 18770 19668 18776
rect 17736 18720 17816 18748
rect 18420 18760 18472 18766
rect 17684 18702 17736 18708
rect 18420 18702 18472 18708
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 19064 18760 19116 18766
rect 19064 18702 19116 18708
rect 17316 17876 17368 17882
rect 17316 17818 17368 17824
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 17328 16998 17356 17818
rect 17696 17202 17724 18702
rect 18206 18524 18502 18544
rect 18262 18522 18286 18524
rect 18342 18522 18366 18524
rect 18422 18522 18446 18524
rect 18284 18470 18286 18522
rect 18348 18470 18360 18522
rect 18422 18470 18424 18522
rect 18262 18468 18286 18470
rect 18342 18468 18366 18470
rect 18422 18468 18446 18470
rect 18206 18448 18502 18468
rect 18800 18086 18828 18702
rect 19076 18290 19104 18702
rect 19168 18358 19196 18770
rect 19156 18352 19208 18358
rect 19156 18294 19208 18300
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18206 17436 18502 17456
rect 18262 17434 18286 17436
rect 18342 17434 18366 17436
rect 18422 17434 18446 17436
rect 18284 17382 18286 17434
rect 18348 17382 18360 17434
rect 18422 17382 18424 17434
rect 18262 17380 18286 17382
rect 18342 17380 18366 17382
rect 18422 17380 18446 17382
rect 18206 17360 18502 17380
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 17592 17060 17644 17066
rect 17592 17002 17644 17008
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 16856 16720 16908 16726
rect 16856 16662 16908 16668
rect 16856 16040 16908 16046
rect 16960 16028 16988 16730
rect 17132 16720 17184 16726
rect 17132 16662 17184 16668
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 16908 16000 16988 16028
rect 16856 15982 16908 15988
rect 16960 15638 16988 16000
rect 17052 15638 17080 16594
rect 17144 15706 17172 16662
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17236 16114 17264 16390
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 17328 15706 17356 16934
rect 17604 16658 17632 17002
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17592 16244 17644 16250
rect 17696 16232 17724 17138
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 17644 16204 17724 16232
rect 17592 16186 17644 16192
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 16948 15632 17000 15638
rect 16948 15574 17000 15580
rect 17040 15632 17092 15638
rect 17040 15574 17092 15580
rect 17144 14618 17172 15642
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 17604 13308 17632 16186
rect 17972 15978 18000 16730
rect 18604 16720 18656 16726
rect 18604 16662 18656 16668
rect 18696 16720 18748 16726
rect 18696 16662 18748 16668
rect 18206 16348 18502 16368
rect 18262 16346 18286 16348
rect 18342 16346 18366 16348
rect 18422 16346 18446 16348
rect 18284 16294 18286 16346
rect 18348 16294 18360 16346
rect 18422 16294 18424 16346
rect 18262 16292 18286 16294
rect 18342 16292 18366 16294
rect 18422 16292 18446 16294
rect 18206 16272 18502 16292
rect 18616 15978 18644 16662
rect 18708 16250 18736 16662
rect 19076 16250 19104 18226
rect 19352 18222 19380 18770
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19444 18222 19472 18702
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 18604 15972 18656 15978
rect 18604 15914 18656 15920
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17696 13462 17724 15642
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18206 15260 18502 15280
rect 18262 15258 18286 15260
rect 18342 15258 18366 15260
rect 18422 15258 18446 15260
rect 18284 15206 18286 15258
rect 18348 15206 18360 15258
rect 18422 15206 18424 15258
rect 18262 15204 18286 15206
rect 18342 15204 18366 15206
rect 18422 15204 18446 15206
rect 18206 15184 18502 15204
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 18064 14006 18092 14418
rect 18206 14172 18502 14192
rect 18262 14170 18286 14172
rect 18342 14170 18366 14172
rect 18422 14170 18446 14172
rect 18284 14118 18286 14170
rect 18348 14118 18360 14170
rect 18422 14118 18424 14170
rect 18262 14116 18286 14118
rect 18342 14116 18366 14118
rect 18422 14116 18446 14118
rect 18206 14096 18502 14116
rect 18052 14000 18104 14006
rect 18052 13942 18104 13948
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17684 13456 17736 13462
rect 17684 13398 17736 13404
rect 17684 13320 17736 13326
rect 17604 13280 17684 13308
rect 17684 13262 17736 13268
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 16764 12912 16816 12918
rect 16764 12854 16816 12860
rect 17328 12782 17356 13126
rect 17696 12850 17724 13262
rect 17880 12986 17908 13806
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 17972 13326 18000 13670
rect 18064 13394 18092 13942
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 18616 13326 18644 15302
rect 18708 14482 18736 16186
rect 18972 15972 19024 15978
rect 18972 15914 19024 15920
rect 18984 14618 19012 15914
rect 19444 15706 19472 18158
rect 19720 16998 19748 20266
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 20640 19514 20668 19926
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20444 19304 20496 19310
rect 20444 19246 20496 19252
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 19812 18222 19840 18566
rect 19800 18216 19852 18222
rect 19800 18158 19852 18164
rect 20456 17746 20484 19246
rect 20444 17740 20496 17746
rect 20444 17682 20496 17688
rect 19984 17060 20036 17066
rect 19984 17002 20036 17008
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19720 16658 19748 16934
rect 19996 16794 20024 17002
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19708 16652 19760 16658
rect 19708 16594 19760 16600
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 19536 16046 19564 16390
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 18972 14612 19024 14618
rect 18972 14554 19024 14560
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18984 14074 19012 14554
rect 19156 14476 19208 14482
rect 19156 14418 19208 14424
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 18696 13796 18748 13802
rect 18696 13738 18748 13744
rect 18708 13394 18736 13738
rect 18984 13462 19012 14010
rect 18972 13456 19024 13462
rect 18972 13398 19024 13404
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 19168 13326 19196 14418
rect 19352 13870 19380 14418
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19352 13462 19380 13806
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 19628 13394 19656 16594
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19904 16046 19932 16390
rect 19892 16040 19944 16046
rect 19892 15982 19944 15988
rect 19984 15972 20036 15978
rect 19984 15914 20036 15920
rect 19996 15502 20024 15914
rect 20168 15700 20220 15706
rect 20168 15642 20220 15648
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19996 14958 20024 15438
rect 20180 14958 20208 15642
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 19892 14884 19944 14890
rect 19892 14826 19944 14832
rect 19904 14482 19932 14826
rect 20180 14618 20208 14894
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20364 14618 20392 14758
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20352 14612 20404 14618
rect 20352 14554 20404 14560
rect 19892 14476 19944 14482
rect 19892 14418 19944 14424
rect 20364 14278 20392 14554
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 20088 13462 20116 14214
rect 20076 13456 20128 13462
rect 20076 13398 20128 13404
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19800 13388 19852 13394
rect 19800 13330 19852 13336
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 19156 13320 19208 13326
rect 19156 13262 19208 13268
rect 18206 13084 18502 13104
rect 18262 13082 18286 13084
rect 18342 13082 18366 13084
rect 18422 13082 18446 13084
rect 18284 13030 18286 13082
rect 18348 13030 18360 13082
rect 18422 13030 18424 13082
rect 18262 13028 18286 13030
rect 18342 13028 18366 13030
rect 18422 13028 18446 13030
rect 18206 13008 18502 13028
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 15844 12368 15896 12374
rect 15844 12310 15896 12316
rect 17696 12306 17724 12786
rect 18616 12714 18644 13262
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18892 12782 18920 13126
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 18604 12708 18656 12714
rect 18604 12650 18656 12656
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17236 10810 17264 10950
rect 17696 10810 17724 11154
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17880 10742 17908 11222
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17972 10538 18000 12650
rect 18206 11996 18502 12016
rect 18262 11994 18286 11996
rect 18342 11994 18366 11996
rect 18422 11994 18446 11996
rect 18284 11942 18286 11994
rect 18348 11942 18360 11994
rect 18422 11942 18424 11994
rect 18262 11940 18286 11942
rect 18342 11940 18366 11942
rect 18422 11940 18446 11942
rect 18206 11920 18502 11940
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18432 11354 18460 11494
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18064 10674 18092 11086
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 18206 10908 18502 10928
rect 18262 10906 18286 10908
rect 18342 10906 18366 10908
rect 18422 10906 18446 10908
rect 18284 10854 18286 10906
rect 18348 10854 18360 10906
rect 18422 10854 18424 10906
rect 18262 10852 18286 10854
rect 18342 10852 18366 10854
rect 18422 10852 18446 10854
rect 18206 10832 18502 10852
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 17960 10532 18012 10538
rect 17960 10474 18012 10480
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 16776 9110 16804 10406
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 14756 8188 15052 8208
rect 14812 8186 14836 8188
rect 14892 8186 14916 8188
rect 14972 8186 14996 8188
rect 14834 8134 14836 8186
rect 14898 8134 14910 8186
rect 14972 8134 14974 8186
rect 14812 8132 14836 8134
rect 14892 8132 14916 8134
rect 14972 8132 14996 8134
rect 14756 8112 15052 8132
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 14384 7818 14412 7890
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 14384 7410 14412 7754
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14476 7342 14504 7890
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14756 7100 15052 7120
rect 14812 7098 14836 7100
rect 14892 7098 14916 7100
rect 14972 7098 14996 7100
rect 14834 7046 14836 7098
rect 14898 7046 14910 7098
rect 14972 7046 14974 7098
rect 14812 7044 14836 7046
rect 14892 7044 14916 7046
rect 14972 7044 14996 7046
rect 14756 7024 15052 7044
rect 13372 6886 13492 6914
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12992 5160 13044 5166
rect 13044 5108 13216 5114
rect 12992 5102 13216 5108
rect 13004 5098 13216 5102
rect 13004 5092 13228 5098
rect 13004 5086 13176 5092
rect 13176 5034 13228 5040
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 13464 2990 13492 6886
rect 14756 6012 15052 6032
rect 14812 6010 14836 6012
rect 14892 6010 14916 6012
rect 14972 6010 14996 6012
rect 14834 5958 14836 6010
rect 14898 5958 14910 6010
rect 14972 5958 14974 6010
rect 14812 5956 14836 5958
rect 14892 5956 14916 5958
rect 14972 5956 14996 5958
rect 14756 5936 15052 5956
rect 15120 5778 15148 8774
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16776 8022 16804 8570
rect 16868 8430 16896 8774
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16764 8016 16816 8022
rect 16764 7958 16816 7964
rect 17236 6866 17264 10202
rect 18206 9820 18502 9840
rect 18262 9818 18286 9820
rect 18342 9818 18366 9820
rect 18422 9818 18446 9820
rect 18284 9766 18286 9818
rect 18348 9766 18360 9818
rect 18422 9766 18424 9818
rect 18262 9764 18286 9766
rect 18342 9764 18366 9766
rect 18422 9764 18446 9766
rect 18206 9744 18502 9764
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 17328 8498 17356 8774
rect 18206 8732 18502 8752
rect 18262 8730 18286 8732
rect 18342 8730 18366 8732
rect 18422 8730 18446 8732
rect 18284 8678 18286 8730
rect 18348 8678 18360 8730
rect 18422 8678 18424 8730
rect 18262 8676 18286 8678
rect 18342 8676 18366 8678
rect 18422 8676 18446 8678
rect 18206 8656 18502 8676
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 18616 8362 18644 8978
rect 18800 8498 18828 11018
rect 19168 10674 19196 12786
rect 19352 12646 19380 12854
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19260 10810 19288 12582
rect 19352 11218 19380 12582
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19812 10810 19840 13330
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19996 12850 20024 13126
rect 20088 12986 20116 13398
rect 20456 13394 20484 17682
rect 20444 13388 20496 13394
rect 20444 13330 20496 13336
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 19984 12844 20036 12850
rect 19984 12786 20036 12792
rect 20456 12730 20484 13330
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20364 12702 20484 12730
rect 20732 12714 20760 13126
rect 20720 12708 20772 12714
rect 20364 12646 20392 12702
rect 20720 12650 20772 12656
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19800 10804 19852 10810
rect 19800 10746 19852 10752
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18206 7644 18502 7664
rect 18262 7642 18286 7644
rect 18342 7642 18366 7644
rect 18422 7642 18446 7644
rect 18284 7590 18286 7642
rect 18348 7590 18360 7642
rect 18422 7590 18424 7642
rect 18262 7588 18286 7590
rect 18342 7588 18366 7590
rect 18422 7588 18446 7590
rect 18206 7568 18502 7588
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 15948 5914 15976 6802
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16224 6322 16252 6734
rect 18206 6556 18502 6576
rect 18262 6554 18286 6556
rect 18342 6554 18366 6556
rect 18422 6554 18446 6556
rect 18284 6502 18286 6554
rect 18348 6502 18360 6554
rect 18422 6502 18424 6554
rect 18262 6500 18286 6502
rect 18342 6500 18366 6502
rect 18422 6500 18446 6502
rect 18206 6480 18502 6500
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 17420 5778 17448 6054
rect 17604 5846 17632 6190
rect 17592 5840 17644 5846
rect 17592 5782 17644 5788
rect 18064 5778 18092 6190
rect 14832 5772 14884 5778
rect 14832 5714 14884 5720
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14752 5166 14780 5510
rect 14844 5166 14872 5714
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15212 5370 15240 5646
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 15304 5030 15332 5646
rect 16960 5370 16988 5714
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 17420 5250 17448 5714
rect 17960 5704 18012 5710
rect 17960 5646 18012 5652
rect 17420 5222 17540 5250
rect 17972 5234 18000 5646
rect 18064 5370 18092 5714
rect 18248 5710 18276 6258
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18432 5778 18460 6190
rect 18696 6180 18748 6186
rect 18696 6122 18748 6128
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18420 5772 18472 5778
rect 18420 5714 18472 5720
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18206 5468 18502 5488
rect 18262 5466 18286 5468
rect 18342 5466 18366 5468
rect 18422 5466 18446 5468
rect 18284 5414 18286 5466
rect 18348 5414 18360 5466
rect 18422 5414 18424 5466
rect 18262 5412 18286 5414
rect 18342 5412 18366 5414
rect 18422 5412 18446 5414
rect 18206 5392 18502 5412
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 14756 4924 15052 4944
rect 14812 4922 14836 4924
rect 14892 4922 14916 4924
rect 14972 4922 14996 4924
rect 14834 4870 14836 4922
rect 14898 4870 14910 4922
rect 14972 4870 14974 4922
rect 14812 4868 14836 4870
rect 14892 4868 14916 4870
rect 14972 4868 14996 4870
rect 14756 4848 15052 4868
rect 15396 4214 15424 5102
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17328 4826 17356 4966
rect 17316 4820 17368 4826
rect 17316 4762 17368 4768
rect 17420 4282 17448 4966
rect 16948 4276 17000 4282
rect 16948 4218 17000 4224
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 15384 4208 15436 4214
rect 15384 4150 15436 4156
rect 15108 4004 15160 4010
rect 15108 3946 15160 3952
rect 14756 3836 15052 3856
rect 14812 3834 14836 3836
rect 14892 3834 14916 3836
rect 14972 3834 14996 3836
rect 14834 3782 14836 3834
rect 14898 3782 14910 3834
rect 14972 3782 14974 3834
rect 14812 3780 14836 3782
rect 14892 3780 14916 3782
rect 14972 3780 14996 3782
rect 14756 3760 15052 3780
rect 15120 3738 15148 3946
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13832 3194 13860 3470
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13832 2990 13860 3130
rect 14476 3126 14504 3674
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 14568 3194 14596 3402
rect 15120 3194 15148 3674
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15580 3194 15608 3470
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 15948 2990 15976 3334
rect 16960 3058 16988 4218
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 11796 2916 11848 2922
rect 11796 2858 11848 2864
rect 12164 2848 12216 2854
rect 12164 2790 12216 2796
rect 12176 2650 12204 2790
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 2044 2576 2096 2582
rect 2044 2518 2096 2524
rect 8208 2576 8260 2582
rect 8208 2518 8260 2524
rect 480 2508 532 2514
rect 480 2450 532 2456
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 492 800 520 2450
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 1872 800 1900 2314
rect 3712 800 3740 2450
rect 4406 2204 4702 2224
rect 4462 2202 4486 2204
rect 4542 2202 4566 2204
rect 4622 2202 4646 2204
rect 4484 2150 4486 2202
rect 4548 2150 4560 2202
rect 4622 2150 4624 2202
rect 4462 2148 4486 2150
rect 4542 2148 4566 2150
rect 4622 2148 4646 2150
rect 4406 2128 4702 2148
rect 5552 800 5580 2450
rect 6932 800 6960 2450
rect 8772 800 8800 2450
rect 10612 800 10640 2450
rect 11306 2204 11602 2224
rect 11362 2202 11386 2204
rect 11442 2202 11466 2204
rect 11522 2202 11546 2204
rect 11384 2150 11386 2202
rect 11448 2150 11460 2202
rect 11522 2150 11524 2202
rect 11362 2148 11386 2150
rect 11442 2148 11466 2150
rect 11522 2148 11546 2150
rect 11306 2128 11602 2148
rect 11992 800 12020 2450
rect 12544 2446 12572 2926
rect 16132 2922 16160 2994
rect 16120 2916 16172 2922
rect 16120 2858 16172 2864
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13832 2650 13860 2790
rect 14756 2748 15052 2768
rect 14812 2746 14836 2748
rect 14892 2746 14916 2748
rect 14972 2746 14996 2748
rect 14834 2694 14836 2746
rect 14898 2694 14910 2746
rect 14972 2694 14974 2746
rect 14812 2692 14836 2694
rect 14892 2692 14916 2694
rect 14972 2692 14996 2694
rect 14756 2672 15052 2692
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 15660 2508 15712 2514
rect 15660 2450 15712 2456
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 13832 800 13860 2450
rect 15672 800 15700 2450
rect 16132 2446 16160 2858
rect 17512 2650 17540 5222
rect 17960 5228 18012 5234
rect 17960 5170 18012 5176
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 17960 3664 18012 3670
rect 17960 3606 18012 3612
rect 17972 3058 18000 3606
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 17052 800 17080 2450
rect 18064 2378 18092 5102
rect 18616 4622 18644 6054
rect 18708 5778 18736 6122
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 18696 5636 18748 5642
rect 18696 5578 18748 5584
rect 18708 5166 18736 5578
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18206 4380 18502 4400
rect 18262 4378 18286 4380
rect 18342 4378 18366 4380
rect 18422 4378 18446 4380
rect 18284 4326 18286 4378
rect 18348 4326 18360 4378
rect 18422 4326 18424 4378
rect 18262 4324 18286 4326
rect 18342 4324 18366 4326
rect 18422 4324 18446 4326
rect 18206 4304 18502 4324
rect 18206 3292 18502 3312
rect 18262 3290 18286 3292
rect 18342 3290 18366 3292
rect 18422 3290 18446 3292
rect 18284 3238 18286 3290
rect 18348 3238 18360 3290
rect 18422 3238 18424 3290
rect 18262 3236 18286 3238
rect 18342 3236 18366 3238
rect 18422 3236 18446 3238
rect 18206 3216 18502 3236
rect 18892 2650 18920 10406
rect 19168 10266 19196 10610
rect 20180 10538 20208 11018
rect 20168 10532 20220 10538
rect 20168 10474 20220 10480
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 20824 5778 20852 22066
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20916 20398 20944 21286
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20916 19854 20944 20334
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 21008 17066 21036 17478
rect 20996 17060 21048 17066
rect 20996 17002 21048 17008
rect 20812 5772 20864 5778
rect 20812 5714 20864 5720
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 18984 4214 19012 4694
rect 19156 4684 19208 4690
rect 19156 4626 19208 4632
rect 18972 4208 19024 4214
rect 18972 4150 19024 4156
rect 18984 3194 19012 4150
rect 19168 3194 19196 4626
rect 21100 4214 21128 20946
rect 21364 20800 21416 20806
rect 21364 20742 21416 20748
rect 21376 20505 21404 20742
rect 21362 20496 21418 20505
rect 21362 20431 21418 20440
rect 21364 20324 21416 20330
rect 21364 20266 21416 20272
rect 21376 20058 21404 20266
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 21192 11150 21220 17478
rect 21284 15706 21312 18226
rect 21454 17776 21510 17785
rect 21454 17711 21456 17720
rect 21508 17711 21510 17720
rect 21456 17682 21508 17688
rect 21454 15736 21510 15745
rect 21272 15700 21324 15706
rect 21454 15671 21510 15680
rect 21272 15642 21324 15648
rect 21468 15570 21496 15671
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21468 13025 21496 13330
rect 21454 13016 21510 13025
rect 21454 12951 21510 12960
rect 21272 11280 21324 11286
rect 21272 11222 21324 11228
rect 21180 11144 21232 11150
rect 21180 11086 21232 11092
rect 21284 10266 21312 11222
rect 21454 10296 21510 10305
rect 21272 10260 21324 10266
rect 21454 10231 21510 10240
rect 21272 10202 21324 10208
rect 21468 10130 21496 10231
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21272 8288 21324 8294
rect 21468 8265 21496 8366
rect 21272 8230 21324 8236
rect 21454 8256 21510 8265
rect 21284 7886 21312 8230
rect 21454 8191 21510 8200
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21456 5772 21508 5778
rect 21456 5714 21508 5720
rect 21468 5545 21496 5714
rect 21454 5536 21510 5545
rect 21454 5471 21510 5480
rect 21088 4208 21140 4214
rect 21088 4150 21140 4156
rect 18972 3188 19024 3194
rect 18972 3130 19024 3136
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 18984 2990 19012 3130
rect 20904 3052 20956 3058
rect 21100 3040 21128 4150
rect 21180 3052 21232 3058
rect 21100 3012 21180 3040
rect 20904 2994 20956 3000
rect 21180 2994 21232 3000
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 20916 2514 20944 2994
rect 21456 2984 21508 2990
rect 21456 2926 21508 2932
rect 21468 2825 21496 2926
rect 21454 2816 21510 2825
rect 21454 2751 21510 2760
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 20904 2508 20956 2514
rect 20904 2450 20956 2456
rect 22100 2508 22152 2514
rect 22100 2450 22152 2456
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 18206 2204 18502 2224
rect 18262 2202 18286 2204
rect 18342 2202 18366 2204
rect 18422 2202 18446 2204
rect 18284 2150 18286 2202
rect 18348 2150 18360 2202
rect 18422 2150 18424 2202
rect 18262 2148 18286 2150
rect 18342 2148 18366 2150
rect 18422 2148 18446 2150
rect 18206 2128 18502 2148
rect 18892 800 18920 2450
rect 20720 2372 20772 2378
rect 20720 2314 20772 2320
rect 20732 800 20760 2314
rect 22112 800 22140 2450
rect 478 0 534 800
rect 1858 0 1914 800
rect 3698 0 3754 800
rect 5538 0 5594 800
rect 6918 0 6974 800
rect 8758 0 8814 800
rect 10598 0 10654 800
rect 11978 0 12034 800
rect 13818 0 13874 800
rect 15658 0 15714 800
rect 17038 0 17094 800
rect 18878 0 18934 800
rect 20718 0 20774 800
rect 22098 0 22154 800
<< via2 >>
rect 1490 23160 1546 23216
rect 4406 22874 4462 22876
rect 4486 22874 4542 22876
rect 4566 22874 4622 22876
rect 4646 22874 4702 22876
rect 4406 22822 4432 22874
rect 4432 22822 4462 22874
rect 4486 22822 4496 22874
rect 4496 22822 4542 22874
rect 4566 22822 4612 22874
rect 4612 22822 4622 22874
rect 4646 22822 4676 22874
rect 4676 22822 4702 22874
rect 4406 22820 4462 22822
rect 4486 22820 4542 22822
rect 4566 22820 4622 22822
rect 4646 22820 4702 22822
rect 1398 20440 1454 20496
rect 1398 17740 1454 17776
rect 1398 17720 1400 17740
rect 1400 17720 1452 17740
rect 1452 17720 1454 17740
rect 1398 15680 1454 15736
rect 1490 12980 1546 13016
rect 1490 12960 1492 12980
rect 1492 12960 1544 12980
rect 1544 12960 1546 12980
rect 1490 10260 1546 10296
rect 1490 10240 1492 10260
rect 1492 10240 1544 10260
rect 1544 10240 1546 10260
rect 4406 21786 4462 21788
rect 4486 21786 4542 21788
rect 4566 21786 4622 21788
rect 4646 21786 4702 21788
rect 4406 21734 4432 21786
rect 4432 21734 4462 21786
rect 4486 21734 4496 21786
rect 4496 21734 4542 21786
rect 4566 21734 4612 21786
rect 4612 21734 4622 21786
rect 4646 21734 4676 21786
rect 4676 21734 4702 21786
rect 4406 21732 4462 21734
rect 4486 21732 4542 21734
rect 4566 21732 4622 21734
rect 4646 21732 4702 21734
rect 4406 20698 4462 20700
rect 4486 20698 4542 20700
rect 4566 20698 4622 20700
rect 4646 20698 4702 20700
rect 4406 20646 4432 20698
rect 4432 20646 4462 20698
rect 4486 20646 4496 20698
rect 4496 20646 4542 20698
rect 4566 20646 4612 20698
rect 4612 20646 4622 20698
rect 4646 20646 4676 20698
rect 4676 20646 4702 20698
rect 4406 20644 4462 20646
rect 4486 20644 4542 20646
rect 4566 20644 4622 20646
rect 4646 20644 4702 20646
rect 4406 19610 4462 19612
rect 4486 19610 4542 19612
rect 4566 19610 4622 19612
rect 4646 19610 4702 19612
rect 4406 19558 4432 19610
rect 4432 19558 4462 19610
rect 4486 19558 4496 19610
rect 4496 19558 4542 19610
rect 4566 19558 4612 19610
rect 4612 19558 4622 19610
rect 4646 19558 4676 19610
rect 4676 19558 4702 19610
rect 4406 19556 4462 19558
rect 4486 19556 4542 19558
rect 4566 19556 4622 19558
rect 4646 19556 4702 19558
rect 4406 18522 4462 18524
rect 4486 18522 4542 18524
rect 4566 18522 4622 18524
rect 4646 18522 4702 18524
rect 4406 18470 4432 18522
rect 4432 18470 4462 18522
rect 4486 18470 4496 18522
rect 4496 18470 4542 18522
rect 4566 18470 4612 18522
rect 4612 18470 4622 18522
rect 4646 18470 4676 18522
rect 4676 18470 4702 18522
rect 4406 18468 4462 18470
rect 4486 18468 4542 18470
rect 4566 18468 4622 18470
rect 4646 18468 4702 18470
rect 4406 17434 4462 17436
rect 4486 17434 4542 17436
rect 4566 17434 4622 17436
rect 4646 17434 4702 17436
rect 4406 17382 4432 17434
rect 4432 17382 4462 17434
rect 4486 17382 4496 17434
rect 4496 17382 4542 17434
rect 4566 17382 4612 17434
rect 4612 17382 4622 17434
rect 4646 17382 4676 17434
rect 4676 17382 4702 17434
rect 4406 17380 4462 17382
rect 4486 17380 4542 17382
rect 4566 17380 4622 17382
rect 4646 17380 4702 17382
rect 4406 16346 4462 16348
rect 4486 16346 4542 16348
rect 4566 16346 4622 16348
rect 4646 16346 4702 16348
rect 4406 16294 4432 16346
rect 4432 16294 4462 16346
rect 4486 16294 4496 16346
rect 4496 16294 4542 16346
rect 4566 16294 4612 16346
rect 4612 16294 4622 16346
rect 4646 16294 4676 16346
rect 4676 16294 4702 16346
rect 4406 16292 4462 16294
rect 4486 16292 4542 16294
rect 4566 16292 4622 16294
rect 4646 16292 4702 16294
rect 1398 8200 1454 8256
rect 4406 15258 4462 15260
rect 4486 15258 4542 15260
rect 4566 15258 4622 15260
rect 4646 15258 4702 15260
rect 4406 15206 4432 15258
rect 4432 15206 4462 15258
rect 4486 15206 4496 15258
rect 4496 15206 4542 15258
rect 4566 15206 4612 15258
rect 4612 15206 4622 15258
rect 4646 15206 4676 15258
rect 4676 15206 4702 15258
rect 4406 15204 4462 15206
rect 4486 15204 4542 15206
rect 4566 15204 4622 15206
rect 4646 15204 4702 15206
rect 4406 14170 4462 14172
rect 4486 14170 4542 14172
rect 4566 14170 4622 14172
rect 4646 14170 4702 14172
rect 4406 14118 4432 14170
rect 4432 14118 4462 14170
rect 4486 14118 4496 14170
rect 4496 14118 4542 14170
rect 4566 14118 4612 14170
rect 4612 14118 4622 14170
rect 4646 14118 4676 14170
rect 4676 14118 4702 14170
rect 4406 14116 4462 14118
rect 4486 14116 4542 14118
rect 4566 14116 4622 14118
rect 4646 14116 4702 14118
rect 11306 22874 11362 22876
rect 11386 22874 11442 22876
rect 11466 22874 11522 22876
rect 11546 22874 11602 22876
rect 11306 22822 11332 22874
rect 11332 22822 11362 22874
rect 11386 22822 11396 22874
rect 11396 22822 11442 22874
rect 11466 22822 11512 22874
rect 11512 22822 11522 22874
rect 11546 22822 11576 22874
rect 11576 22822 11602 22874
rect 11306 22820 11362 22822
rect 11386 22820 11442 22822
rect 11466 22820 11522 22822
rect 11546 22820 11602 22822
rect 4406 13082 4462 13084
rect 4486 13082 4542 13084
rect 4566 13082 4622 13084
rect 4646 13082 4702 13084
rect 4406 13030 4432 13082
rect 4432 13030 4462 13082
rect 4486 13030 4496 13082
rect 4496 13030 4542 13082
rect 4566 13030 4612 13082
rect 4612 13030 4622 13082
rect 4646 13030 4676 13082
rect 4676 13030 4702 13082
rect 4406 13028 4462 13030
rect 4486 13028 4542 13030
rect 4566 13028 4622 13030
rect 4646 13028 4702 13030
rect 1490 5516 1492 5536
rect 1492 5516 1544 5536
rect 1544 5516 1546 5536
rect 1490 5480 1546 5516
rect 4406 11994 4462 11996
rect 4486 11994 4542 11996
rect 4566 11994 4622 11996
rect 4646 11994 4702 11996
rect 4406 11942 4432 11994
rect 4432 11942 4462 11994
rect 4486 11942 4496 11994
rect 4496 11942 4542 11994
rect 4566 11942 4612 11994
rect 4612 11942 4622 11994
rect 4646 11942 4676 11994
rect 4676 11942 4702 11994
rect 4406 11940 4462 11942
rect 4486 11940 4542 11942
rect 4566 11940 4622 11942
rect 4646 11940 4702 11942
rect 4406 10906 4462 10908
rect 4486 10906 4542 10908
rect 4566 10906 4622 10908
rect 4646 10906 4702 10908
rect 4406 10854 4432 10906
rect 4432 10854 4462 10906
rect 4486 10854 4496 10906
rect 4496 10854 4542 10906
rect 4566 10854 4612 10906
rect 4612 10854 4622 10906
rect 4646 10854 4676 10906
rect 4676 10854 4702 10906
rect 4406 10852 4462 10854
rect 4486 10852 4542 10854
rect 4566 10852 4622 10854
rect 4646 10852 4702 10854
rect 4406 9818 4462 9820
rect 4486 9818 4542 9820
rect 4566 9818 4622 9820
rect 4646 9818 4702 9820
rect 4406 9766 4432 9818
rect 4432 9766 4462 9818
rect 4486 9766 4496 9818
rect 4496 9766 4542 9818
rect 4566 9766 4612 9818
rect 4612 9766 4622 9818
rect 4646 9766 4676 9818
rect 4676 9766 4702 9818
rect 4406 9764 4462 9766
rect 4486 9764 4542 9766
rect 4566 9764 4622 9766
rect 4646 9764 4702 9766
rect 4406 8730 4462 8732
rect 4486 8730 4542 8732
rect 4566 8730 4622 8732
rect 4646 8730 4702 8732
rect 4406 8678 4432 8730
rect 4432 8678 4462 8730
rect 4486 8678 4496 8730
rect 4496 8678 4542 8730
rect 4566 8678 4612 8730
rect 4612 8678 4622 8730
rect 4646 8678 4676 8730
rect 4676 8678 4702 8730
rect 4406 8676 4462 8678
rect 4486 8676 4542 8678
rect 4566 8676 4622 8678
rect 4646 8676 4702 8678
rect 1398 2760 1454 2816
rect 4406 7642 4462 7644
rect 4486 7642 4542 7644
rect 4566 7642 4622 7644
rect 4646 7642 4702 7644
rect 4406 7590 4432 7642
rect 4432 7590 4462 7642
rect 4486 7590 4496 7642
rect 4496 7590 4542 7642
rect 4566 7590 4612 7642
rect 4612 7590 4622 7642
rect 4646 7590 4676 7642
rect 4676 7590 4702 7642
rect 4406 7588 4462 7590
rect 4486 7588 4542 7590
rect 4566 7588 4622 7590
rect 4646 7588 4702 7590
rect 4406 6554 4462 6556
rect 4486 6554 4542 6556
rect 4566 6554 4622 6556
rect 4646 6554 4702 6556
rect 4406 6502 4432 6554
rect 4432 6502 4462 6554
rect 4486 6502 4496 6554
rect 4496 6502 4542 6554
rect 4566 6502 4612 6554
rect 4612 6502 4622 6554
rect 4646 6502 4676 6554
rect 4676 6502 4702 6554
rect 4406 6500 4462 6502
rect 4486 6500 4542 6502
rect 4566 6500 4622 6502
rect 4646 6500 4702 6502
rect 4406 5466 4462 5468
rect 4486 5466 4542 5468
rect 4566 5466 4622 5468
rect 4646 5466 4702 5468
rect 4406 5414 4432 5466
rect 4432 5414 4462 5466
rect 4486 5414 4496 5466
rect 4496 5414 4542 5466
rect 4566 5414 4612 5466
rect 4612 5414 4622 5466
rect 4646 5414 4676 5466
rect 4676 5414 4702 5466
rect 4406 5412 4462 5414
rect 4486 5412 4542 5414
rect 4566 5412 4622 5414
rect 4646 5412 4702 5414
rect 4406 4378 4462 4380
rect 4486 4378 4542 4380
rect 4566 4378 4622 4380
rect 4646 4378 4702 4380
rect 4406 4326 4432 4378
rect 4432 4326 4462 4378
rect 4486 4326 4496 4378
rect 4496 4326 4542 4378
rect 4566 4326 4612 4378
rect 4612 4326 4622 4378
rect 4646 4326 4676 4378
rect 4676 4326 4702 4378
rect 4406 4324 4462 4326
rect 4486 4324 4542 4326
rect 4566 4324 4622 4326
rect 4646 4324 4702 4326
rect 4406 3290 4462 3292
rect 4486 3290 4542 3292
rect 4566 3290 4622 3292
rect 4646 3290 4702 3292
rect 4406 3238 4432 3290
rect 4432 3238 4462 3290
rect 4486 3238 4496 3290
rect 4496 3238 4542 3290
rect 4566 3238 4612 3290
rect 4612 3238 4622 3290
rect 4646 3238 4676 3290
rect 4676 3238 4702 3290
rect 4406 3236 4462 3238
rect 4486 3236 4542 3238
rect 4566 3236 4622 3238
rect 4646 3236 4702 3238
rect 7856 22330 7912 22332
rect 7936 22330 7992 22332
rect 8016 22330 8072 22332
rect 8096 22330 8152 22332
rect 7856 22278 7882 22330
rect 7882 22278 7912 22330
rect 7936 22278 7946 22330
rect 7946 22278 7992 22330
rect 8016 22278 8062 22330
rect 8062 22278 8072 22330
rect 8096 22278 8126 22330
rect 8126 22278 8152 22330
rect 7856 22276 7912 22278
rect 7936 22276 7992 22278
rect 8016 22276 8072 22278
rect 8096 22276 8152 22278
rect 7856 21242 7912 21244
rect 7936 21242 7992 21244
rect 8016 21242 8072 21244
rect 8096 21242 8152 21244
rect 7856 21190 7882 21242
rect 7882 21190 7912 21242
rect 7936 21190 7946 21242
rect 7946 21190 7992 21242
rect 8016 21190 8062 21242
rect 8062 21190 8072 21242
rect 8096 21190 8126 21242
rect 8126 21190 8152 21242
rect 7856 21188 7912 21190
rect 7936 21188 7992 21190
rect 8016 21188 8072 21190
rect 8096 21188 8152 21190
rect 7562 19252 7564 19272
rect 7564 19252 7616 19272
rect 7616 19252 7618 19272
rect 7562 19216 7618 19252
rect 7856 20154 7912 20156
rect 7936 20154 7992 20156
rect 8016 20154 8072 20156
rect 8096 20154 8152 20156
rect 7856 20102 7882 20154
rect 7882 20102 7912 20154
rect 7936 20102 7946 20154
rect 7946 20102 7992 20154
rect 8016 20102 8062 20154
rect 8062 20102 8072 20154
rect 8096 20102 8126 20154
rect 8126 20102 8152 20154
rect 7856 20100 7912 20102
rect 7936 20100 7992 20102
rect 8016 20100 8072 20102
rect 8096 20100 8152 20102
rect 7856 19066 7912 19068
rect 7936 19066 7992 19068
rect 8016 19066 8072 19068
rect 8096 19066 8152 19068
rect 7856 19014 7882 19066
rect 7882 19014 7912 19066
rect 7936 19014 7946 19066
rect 7946 19014 7992 19066
rect 8016 19014 8062 19066
rect 8062 19014 8072 19066
rect 8096 19014 8126 19066
rect 8126 19014 8152 19066
rect 7856 19012 7912 19014
rect 7936 19012 7992 19014
rect 8016 19012 8072 19014
rect 8096 19012 8152 19014
rect 7856 17978 7912 17980
rect 7936 17978 7992 17980
rect 8016 17978 8072 17980
rect 8096 17978 8152 17980
rect 7856 17926 7882 17978
rect 7882 17926 7912 17978
rect 7936 17926 7946 17978
rect 7946 17926 7992 17978
rect 8016 17926 8062 17978
rect 8062 17926 8072 17978
rect 8096 17926 8126 17978
rect 8126 17926 8152 17978
rect 7856 17924 7912 17926
rect 7936 17924 7992 17926
rect 8016 17924 8072 17926
rect 8096 17924 8152 17926
rect 8298 19252 8300 19272
rect 8300 19252 8352 19272
rect 8352 19252 8354 19272
rect 8298 19216 8354 19252
rect 8574 19216 8630 19272
rect 7856 16890 7912 16892
rect 7936 16890 7992 16892
rect 8016 16890 8072 16892
rect 8096 16890 8152 16892
rect 7856 16838 7882 16890
rect 7882 16838 7912 16890
rect 7936 16838 7946 16890
rect 7946 16838 7992 16890
rect 8016 16838 8062 16890
rect 8062 16838 8072 16890
rect 8096 16838 8126 16890
rect 8126 16838 8152 16890
rect 7856 16836 7912 16838
rect 7936 16836 7992 16838
rect 8016 16836 8072 16838
rect 8096 16836 8152 16838
rect 7856 15802 7912 15804
rect 7936 15802 7992 15804
rect 8016 15802 8072 15804
rect 8096 15802 8152 15804
rect 7856 15750 7882 15802
rect 7882 15750 7912 15802
rect 7936 15750 7946 15802
rect 7946 15750 7992 15802
rect 8016 15750 8062 15802
rect 8062 15750 8072 15802
rect 8096 15750 8126 15802
rect 8126 15750 8152 15802
rect 7856 15748 7912 15750
rect 7936 15748 7992 15750
rect 8016 15748 8072 15750
rect 8096 15748 8152 15750
rect 7856 14714 7912 14716
rect 7936 14714 7992 14716
rect 8016 14714 8072 14716
rect 8096 14714 8152 14716
rect 7856 14662 7882 14714
rect 7882 14662 7912 14714
rect 7936 14662 7946 14714
rect 7946 14662 7992 14714
rect 8016 14662 8062 14714
rect 8062 14662 8072 14714
rect 8096 14662 8126 14714
rect 8126 14662 8152 14714
rect 7856 14660 7912 14662
rect 7936 14660 7992 14662
rect 8016 14660 8072 14662
rect 8096 14660 8152 14662
rect 7856 13626 7912 13628
rect 7936 13626 7992 13628
rect 8016 13626 8072 13628
rect 8096 13626 8152 13628
rect 7856 13574 7882 13626
rect 7882 13574 7912 13626
rect 7936 13574 7946 13626
rect 7946 13574 7992 13626
rect 8016 13574 8062 13626
rect 8062 13574 8072 13626
rect 8096 13574 8126 13626
rect 8126 13574 8152 13626
rect 7856 13572 7912 13574
rect 7936 13572 7992 13574
rect 8016 13572 8072 13574
rect 8096 13572 8152 13574
rect 7856 12538 7912 12540
rect 7936 12538 7992 12540
rect 8016 12538 8072 12540
rect 8096 12538 8152 12540
rect 7856 12486 7882 12538
rect 7882 12486 7912 12538
rect 7936 12486 7946 12538
rect 7946 12486 7992 12538
rect 8016 12486 8062 12538
rect 8062 12486 8072 12538
rect 8096 12486 8126 12538
rect 8126 12486 8152 12538
rect 7856 12484 7912 12486
rect 7936 12484 7992 12486
rect 8016 12484 8072 12486
rect 8096 12484 8152 12486
rect 7856 11450 7912 11452
rect 7936 11450 7992 11452
rect 8016 11450 8072 11452
rect 8096 11450 8152 11452
rect 7856 11398 7882 11450
rect 7882 11398 7912 11450
rect 7936 11398 7946 11450
rect 7946 11398 7992 11450
rect 8016 11398 8062 11450
rect 8062 11398 8072 11450
rect 8096 11398 8126 11450
rect 8126 11398 8152 11450
rect 7856 11396 7912 11398
rect 7936 11396 7992 11398
rect 8016 11396 8072 11398
rect 8096 11396 8152 11398
rect 7856 10362 7912 10364
rect 7936 10362 7992 10364
rect 8016 10362 8072 10364
rect 8096 10362 8152 10364
rect 7856 10310 7882 10362
rect 7882 10310 7912 10362
rect 7936 10310 7946 10362
rect 7946 10310 7992 10362
rect 8016 10310 8062 10362
rect 8062 10310 8072 10362
rect 8096 10310 8126 10362
rect 8126 10310 8152 10362
rect 7856 10308 7912 10310
rect 7936 10308 7992 10310
rect 8016 10308 8072 10310
rect 8096 10308 8152 10310
rect 7856 9274 7912 9276
rect 7936 9274 7992 9276
rect 8016 9274 8072 9276
rect 8096 9274 8152 9276
rect 7856 9222 7882 9274
rect 7882 9222 7912 9274
rect 7936 9222 7946 9274
rect 7946 9222 7992 9274
rect 8016 9222 8062 9274
rect 8062 9222 8072 9274
rect 8096 9222 8126 9274
rect 8126 9222 8152 9274
rect 7856 9220 7912 9222
rect 7936 9220 7992 9222
rect 8016 9220 8072 9222
rect 8096 9220 8152 9222
rect 7856 8186 7912 8188
rect 7936 8186 7992 8188
rect 8016 8186 8072 8188
rect 8096 8186 8152 8188
rect 7856 8134 7882 8186
rect 7882 8134 7912 8186
rect 7936 8134 7946 8186
rect 7946 8134 7992 8186
rect 8016 8134 8062 8186
rect 8062 8134 8072 8186
rect 8096 8134 8126 8186
rect 8126 8134 8152 8186
rect 7856 8132 7912 8134
rect 7936 8132 7992 8134
rect 8016 8132 8072 8134
rect 8096 8132 8152 8134
rect 7856 7098 7912 7100
rect 7936 7098 7992 7100
rect 8016 7098 8072 7100
rect 8096 7098 8152 7100
rect 7856 7046 7882 7098
rect 7882 7046 7912 7098
rect 7936 7046 7946 7098
rect 7946 7046 7992 7098
rect 8016 7046 8062 7098
rect 8062 7046 8072 7098
rect 8096 7046 8126 7098
rect 8126 7046 8152 7098
rect 7856 7044 7912 7046
rect 7936 7044 7992 7046
rect 8016 7044 8072 7046
rect 8096 7044 8152 7046
rect 7856 6010 7912 6012
rect 7936 6010 7992 6012
rect 8016 6010 8072 6012
rect 8096 6010 8152 6012
rect 7856 5958 7882 6010
rect 7882 5958 7912 6010
rect 7936 5958 7946 6010
rect 7946 5958 7992 6010
rect 8016 5958 8062 6010
rect 8062 5958 8072 6010
rect 8096 5958 8126 6010
rect 8126 5958 8152 6010
rect 7856 5956 7912 5958
rect 7936 5956 7992 5958
rect 8016 5956 8072 5958
rect 8096 5956 8152 5958
rect 7856 4922 7912 4924
rect 7936 4922 7992 4924
rect 8016 4922 8072 4924
rect 8096 4922 8152 4924
rect 7856 4870 7882 4922
rect 7882 4870 7912 4922
rect 7936 4870 7946 4922
rect 7946 4870 7992 4922
rect 8016 4870 8062 4922
rect 8062 4870 8072 4922
rect 8096 4870 8126 4922
rect 8126 4870 8152 4922
rect 7856 4868 7912 4870
rect 7936 4868 7992 4870
rect 8016 4868 8072 4870
rect 8096 4868 8152 4870
rect 7856 3834 7912 3836
rect 7936 3834 7992 3836
rect 8016 3834 8072 3836
rect 8096 3834 8152 3836
rect 7856 3782 7882 3834
rect 7882 3782 7912 3834
rect 7936 3782 7946 3834
rect 7946 3782 7992 3834
rect 8016 3782 8062 3834
rect 8062 3782 8072 3834
rect 8096 3782 8126 3834
rect 8126 3782 8152 3834
rect 7856 3780 7912 3782
rect 7936 3780 7992 3782
rect 8016 3780 8072 3782
rect 8096 3780 8152 3782
rect 7856 2746 7912 2748
rect 7936 2746 7992 2748
rect 8016 2746 8072 2748
rect 8096 2746 8152 2748
rect 7856 2694 7882 2746
rect 7882 2694 7912 2746
rect 7936 2694 7946 2746
rect 7946 2694 7992 2746
rect 8016 2694 8062 2746
rect 8062 2694 8072 2746
rect 8096 2694 8126 2746
rect 8126 2694 8152 2746
rect 7856 2692 7912 2694
rect 7936 2692 7992 2694
rect 8016 2692 8072 2694
rect 8096 2692 8152 2694
rect 11306 21786 11362 21788
rect 11386 21786 11442 21788
rect 11466 21786 11522 21788
rect 11546 21786 11602 21788
rect 11306 21734 11332 21786
rect 11332 21734 11362 21786
rect 11386 21734 11396 21786
rect 11396 21734 11442 21786
rect 11466 21734 11512 21786
rect 11512 21734 11522 21786
rect 11546 21734 11576 21786
rect 11576 21734 11602 21786
rect 11306 21732 11362 21734
rect 11386 21732 11442 21734
rect 11466 21732 11522 21734
rect 11546 21732 11602 21734
rect 11306 20698 11362 20700
rect 11386 20698 11442 20700
rect 11466 20698 11522 20700
rect 11546 20698 11602 20700
rect 11306 20646 11332 20698
rect 11332 20646 11362 20698
rect 11386 20646 11396 20698
rect 11396 20646 11442 20698
rect 11466 20646 11512 20698
rect 11512 20646 11522 20698
rect 11546 20646 11576 20698
rect 11576 20646 11602 20698
rect 11306 20644 11362 20646
rect 11386 20644 11442 20646
rect 11466 20644 11522 20646
rect 11546 20644 11602 20646
rect 11306 19610 11362 19612
rect 11386 19610 11442 19612
rect 11466 19610 11522 19612
rect 11546 19610 11602 19612
rect 11306 19558 11332 19610
rect 11332 19558 11362 19610
rect 11386 19558 11396 19610
rect 11396 19558 11442 19610
rect 11466 19558 11512 19610
rect 11512 19558 11522 19610
rect 11546 19558 11576 19610
rect 11576 19558 11602 19610
rect 11306 19556 11362 19558
rect 11386 19556 11442 19558
rect 11466 19556 11522 19558
rect 11546 19556 11602 19558
rect 11306 18522 11362 18524
rect 11386 18522 11442 18524
rect 11466 18522 11522 18524
rect 11546 18522 11602 18524
rect 11306 18470 11332 18522
rect 11332 18470 11362 18522
rect 11386 18470 11396 18522
rect 11396 18470 11442 18522
rect 11466 18470 11512 18522
rect 11512 18470 11522 18522
rect 11546 18470 11576 18522
rect 11576 18470 11602 18522
rect 11306 18468 11362 18470
rect 11386 18468 11442 18470
rect 11466 18468 11522 18470
rect 11546 18468 11602 18470
rect 18206 22874 18262 22876
rect 18286 22874 18342 22876
rect 18366 22874 18422 22876
rect 18446 22874 18502 22876
rect 18206 22822 18232 22874
rect 18232 22822 18262 22874
rect 18286 22822 18296 22874
rect 18296 22822 18342 22874
rect 18366 22822 18412 22874
rect 18412 22822 18422 22874
rect 18446 22822 18476 22874
rect 18476 22822 18502 22874
rect 18206 22820 18262 22822
rect 18286 22820 18342 22822
rect 18366 22820 18422 22822
rect 18446 22820 18502 22822
rect 21086 23160 21142 23216
rect 11306 17434 11362 17436
rect 11386 17434 11442 17436
rect 11466 17434 11522 17436
rect 11546 17434 11602 17436
rect 11306 17382 11332 17434
rect 11332 17382 11362 17434
rect 11386 17382 11396 17434
rect 11396 17382 11442 17434
rect 11466 17382 11512 17434
rect 11512 17382 11522 17434
rect 11546 17382 11576 17434
rect 11576 17382 11602 17434
rect 11306 17380 11362 17382
rect 11386 17380 11442 17382
rect 11466 17380 11522 17382
rect 11546 17380 11602 17382
rect 11306 16346 11362 16348
rect 11386 16346 11442 16348
rect 11466 16346 11522 16348
rect 11546 16346 11602 16348
rect 11306 16294 11332 16346
rect 11332 16294 11362 16346
rect 11386 16294 11396 16346
rect 11396 16294 11442 16346
rect 11466 16294 11512 16346
rect 11512 16294 11522 16346
rect 11546 16294 11576 16346
rect 11576 16294 11602 16346
rect 11306 16292 11362 16294
rect 11386 16292 11442 16294
rect 11466 16292 11522 16294
rect 11546 16292 11602 16294
rect 11306 15258 11362 15260
rect 11386 15258 11442 15260
rect 11466 15258 11522 15260
rect 11546 15258 11602 15260
rect 11306 15206 11332 15258
rect 11332 15206 11362 15258
rect 11386 15206 11396 15258
rect 11396 15206 11442 15258
rect 11466 15206 11512 15258
rect 11512 15206 11522 15258
rect 11546 15206 11576 15258
rect 11576 15206 11602 15258
rect 11306 15204 11362 15206
rect 11386 15204 11442 15206
rect 11466 15204 11522 15206
rect 11546 15204 11602 15206
rect 11306 14170 11362 14172
rect 11386 14170 11442 14172
rect 11466 14170 11522 14172
rect 11546 14170 11602 14172
rect 11306 14118 11332 14170
rect 11332 14118 11362 14170
rect 11386 14118 11396 14170
rect 11396 14118 11442 14170
rect 11466 14118 11512 14170
rect 11512 14118 11522 14170
rect 11546 14118 11576 14170
rect 11576 14118 11602 14170
rect 11306 14116 11362 14118
rect 11386 14116 11442 14118
rect 11466 14116 11522 14118
rect 11546 14116 11602 14118
rect 11306 13082 11362 13084
rect 11386 13082 11442 13084
rect 11466 13082 11522 13084
rect 11546 13082 11602 13084
rect 11306 13030 11332 13082
rect 11332 13030 11362 13082
rect 11386 13030 11396 13082
rect 11396 13030 11442 13082
rect 11466 13030 11512 13082
rect 11512 13030 11522 13082
rect 11546 13030 11576 13082
rect 11576 13030 11602 13082
rect 11306 13028 11362 13030
rect 11386 13028 11442 13030
rect 11466 13028 11522 13030
rect 11546 13028 11602 13030
rect 11306 11994 11362 11996
rect 11386 11994 11442 11996
rect 11466 11994 11522 11996
rect 11546 11994 11602 11996
rect 11306 11942 11332 11994
rect 11332 11942 11362 11994
rect 11386 11942 11396 11994
rect 11396 11942 11442 11994
rect 11466 11942 11512 11994
rect 11512 11942 11522 11994
rect 11546 11942 11576 11994
rect 11576 11942 11602 11994
rect 11306 11940 11362 11942
rect 11386 11940 11442 11942
rect 11466 11940 11522 11942
rect 11546 11940 11602 11942
rect 11306 10906 11362 10908
rect 11386 10906 11442 10908
rect 11466 10906 11522 10908
rect 11546 10906 11602 10908
rect 11306 10854 11332 10906
rect 11332 10854 11362 10906
rect 11386 10854 11396 10906
rect 11396 10854 11442 10906
rect 11466 10854 11512 10906
rect 11512 10854 11522 10906
rect 11546 10854 11576 10906
rect 11576 10854 11602 10906
rect 11306 10852 11362 10854
rect 11386 10852 11442 10854
rect 11466 10852 11522 10854
rect 11546 10852 11602 10854
rect 11306 9818 11362 9820
rect 11386 9818 11442 9820
rect 11466 9818 11522 9820
rect 11546 9818 11602 9820
rect 11306 9766 11332 9818
rect 11332 9766 11362 9818
rect 11386 9766 11396 9818
rect 11396 9766 11442 9818
rect 11466 9766 11512 9818
rect 11512 9766 11522 9818
rect 11546 9766 11576 9818
rect 11576 9766 11602 9818
rect 11306 9764 11362 9766
rect 11386 9764 11442 9766
rect 11466 9764 11522 9766
rect 11546 9764 11602 9766
rect 11306 8730 11362 8732
rect 11386 8730 11442 8732
rect 11466 8730 11522 8732
rect 11546 8730 11602 8732
rect 11306 8678 11332 8730
rect 11332 8678 11362 8730
rect 11386 8678 11396 8730
rect 11396 8678 11442 8730
rect 11466 8678 11512 8730
rect 11512 8678 11522 8730
rect 11546 8678 11576 8730
rect 11576 8678 11602 8730
rect 11306 8676 11362 8678
rect 11386 8676 11442 8678
rect 11466 8676 11522 8678
rect 11546 8676 11602 8678
rect 11306 7642 11362 7644
rect 11386 7642 11442 7644
rect 11466 7642 11522 7644
rect 11546 7642 11602 7644
rect 11306 7590 11332 7642
rect 11332 7590 11362 7642
rect 11386 7590 11396 7642
rect 11396 7590 11442 7642
rect 11466 7590 11512 7642
rect 11512 7590 11522 7642
rect 11546 7590 11576 7642
rect 11576 7590 11602 7642
rect 11306 7588 11362 7590
rect 11386 7588 11442 7590
rect 11466 7588 11522 7590
rect 11546 7588 11602 7590
rect 14756 22330 14812 22332
rect 14836 22330 14892 22332
rect 14916 22330 14972 22332
rect 14996 22330 15052 22332
rect 14756 22278 14782 22330
rect 14782 22278 14812 22330
rect 14836 22278 14846 22330
rect 14846 22278 14892 22330
rect 14916 22278 14962 22330
rect 14962 22278 14972 22330
rect 14996 22278 15026 22330
rect 15026 22278 15052 22330
rect 14756 22276 14812 22278
rect 14836 22276 14892 22278
rect 14916 22276 14972 22278
rect 14996 22276 15052 22278
rect 14756 21242 14812 21244
rect 14836 21242 14892 21244
rect 14916 21242 14972 21244
rect 14996 21242 15052 21244
rect 14756 21190 14782 21242
rect 14782 21190 14812 21242
rect 14836 21190 14846 21242
rect 14846 21190 14892 21242
rect 14916 21190 14962 21242
rect 14962 21190 14972 21242
rect 14996 21190 15026 21242
rect 15026 21190 15052 21242
rect 14756 21188 14812 21190
rect 14836 21188 14892 21190
rect 14916 21188 14972 21190
rect 14996 21188 15052 21190
rect 14756 20154 14812 20156
rect 14836 20154 14892 20156
rect 14916 20154 14972 20156
rect 14996 20154 15052 20156
rect 14756 20102 14782 20154
rect 14782 20102 14812 20154
rect 14836 20102 14846 20154
rect 14846 20102 14892 20154
rect 14916 20102 14962 20154
rect 14962 20102 14972 20154
rect 14996 20102 15026 20154
rect 15026 20102 15052 20154
rect 14756 20100 14812 20102
rect 14836 20100 14892 20102
rect 14916 20100 14972 20102
rect 14996 20100 15052 20102
rect 14756 19066 14812 19068
rect 14836 19066 14892 19068
rect 14916 19066 14972 19068
rect 14996 19066 15052 19068
rect 14756 19014 14782 19066
rect 14782 19014 14812 19066
rect 14836 19014 14846 19066
rect 14846 19014 14892 19066
rect 14916 19014 14962 19066
rect 14962 19014 14972 19066
rect 14996 19014 15026 19066
rect 15026 19014 15052 19066
rect 14756 19012 14812 19014
rect 14836 19012 14892 19014
rect 14916 19012 14972 19014
rect 14996 19012 15052 19014
rect 14756 17978 14812 17980
rect 14836 17978 14892 17980
rect 14916 17978 14972 17980
rect 14996 17978 15052 17980
rect 14756 17926 14782 17978
rect 14782 17926 14812 17978
rect 14836 17926 14846 17978
rect 14846 17926 14892 17978
rect 14916 17926 14962 17978
rect 14962 17926 14972 17978
rect 14996 17926 15026 17978
rect 15026 17926 15052 17978
rect 14756 17924 14812 17926
rect 14836 17924 14892 17926
rect 14916 17924 14972 17926
rect 14996 17924 15052 17926
rect 14756 16890 14812 16892
rect 14836 16890 14892 16892
rect 14916 16890 14972 16892
rect 14996 16890 15052 16892
rect 14756 16838 14782 16890
rect 14782 16838 14812 16890
rect 14836 16838 14846 16890
rect 14846 16838 14892 16890
rect 14916 16838 14962 16890
rect 14962 16838 14972 16890
rect 14996 16838 15026 16890
rect 15026 16838 15052 16890
rect 14756 16836 14812 16838
rect 14836 16836 14892 16838
rect 14916 16836 14972 16838
rect 14996 16836 15052 16838
rect 14756 15802 14812 15804
rect 14836 15802 14892 15804
rect 14916 15802 14972 15804
rect 14996 15802 15052 15804
rect 14756 15750 14782 15802
rect 14782 15750 14812 15802
rect 14836 15750 14846 15802
rect 14846 15750 14892 15802
rect 14916 15750 14962 15802
rect 14962 15750 14972 15802
rect 14996 15750 15026 15802
rect 15026 15750 15052 15802
rect 14756 15748 14812 15750
rect 14836 15748 14892 15750
rect 14916 15748 14972 15750
rect 14996 15748 15052 15750
rect 14756 14714 14812 14716
rect 14836 14714 14892 14716
rect 14916 14714 14972 14716
rect 14996 14714 15052 14716
rect 14756 14662 14782 14714
rect 14782 14662 14812 14714
rect 14836 14662 14846 14714
rect 14846 14662 14892 14714
rect 14916 14662 14962 14714
rect 14962 14662 14972 14714
rect 14996 14662 15026 14714
rect 15026 14662 15052 14714
rect 14756 14660 14812 14662
rect 14836 14660 14892 14662
rect 14916 14660 14972 14662
rect 14996 14660 15052 14662
rect 14756 13626 14812 13628
rect 14836 13626 14892 13628
rect 14916 13626 14972 13628
rect 14996 13626 15052 13628
rect 14756 13574 14782 13626
rect 14782 13574 14812 13626
rect 14836 13574 14846 13626
rect 14846 13574 14892 13626
rect 14916 13574 14962 13626
rect 14962 13574 14972 13626
rect 14996 13574 15026 13626
rect 15026 13574 15052 13626
rect 14756 13572 14812 13574
rect 14836 13572 14892 13574
rect 14916 13572 14972 13574
rect 14996 13572 15052 13574
rect 11306 6554 11362 6556
rect 11386 6554 11442 6556
rect 11466 6554 11522 6556
rect 11546 6554 11602 6556
rect 11306 6502 11332 6554
rect 11332 6502 11362 6554
rect 11386 6502 11396 6554
rect 11396 6502 11442 6554
rect 11466 6502 11512 6554
rect 11512 6502 11522 6554
rect 11546 6502 11576 6554
rect 11576 6502 11602 6554
rect 11306 6500 11362 6502
rect 11386 6500 11442 6502
rect 11466 6500 11522 6502
rect 11546 6500 11602 6502
rect 11306 5466 11362 5468
rect 11386 5466 11442 5468
rect 11466 5466 11522 5468
rect 11546 5466 11602 5468
rect 11306 5414 11332 5466
rect 11332 5414 11362 5466
rect 11386 5414 11396 5466
rect 11396 5414 11442 5466
rect 11466 5414 11512 5466
rect 11512 5414 11522 5466
rect 11546 5414 11576 5466
rect 11576 5414 11602 5466
rect 11306 5412 11362 5414
rect 11386 5412 11442 5414
rect 11466 5412 11522 5414
rect 11546 5412 11602 5414
rect 11306 4378 11362 4380
rect 11386 4378 11442 4380
rect 11466 4378 11522 4380
rect 11546 4378 11602 4380
rect 11306 4326 11332 4378
rect 11332 4326 11362 4378
rect 11386 4326 11396 4378
rect 11396 4326 11442 4378
rect 11466 4326 11512 4378
rect 11512 4326 11522 4378
rect 11546 4326 11576 4378
rect 11576 4326 11602 4378
rect 11306 4324 11362 4326
rect 11386 4324 11442 4326
rect 11466 4324 11522 4326
rect 11546 4324 11602 4326
rect 11306 3290 11362 3292
rect 11386 3290 11442 3292
rect 11466 3290 11522 3292
rect 11546 3290 11602 3292
rect 11306 3238 11332 3290
rect 11332 3238 11362 3290
rect 11386 3238 11396 3290
rect 11396 3238 11442 3290
rect 11466 3238 11512 3290
rect 11512 3238 11522 3290
rect 11546 3238 11576 3290
rect 11576 3238 11602 3290
rect 11306 3236 11362 3238
rect 11386 3236 11442 3238
rect 11466 3236 11522 3238
rect 11546 3236 11602 3238
rect 14756 12538 14812 12540
rect 14836 12538 14892 12540
rect 14916 12538 14972 12540
rect 14996 12538 15052 12540
rect 14756 12486 14782 12538
rect 14782 12486 14812 12538
rect 14836 12486 14846 12538
rect 14846 12486 14892 12538
rect 14916 12486 14962 12538
rect 14962 12486 14972 12538
rect 14996 12486 15026 12538
rect 15026 12486 15052 12538
rect 14756 12484 14812 12486
rect 14836 12484 14892 12486
rect 14916 12484 14972 12486
rect 14996 12484 15052 12486
rect 14756 11450 14812 11452
rect 14836 11450 14892 11452
rect 14916 11450 14972 11452
rect 14996 11450 15052 11452
rect 14756 11398 14782 11450
rect 14782 11398 14812 11450
rect 14836 11398 14846 11450
rect 14846 11398 14892 11450
rect 14916 11398 14962 11450
rect 14962 11398 14972 11450
rect 14996 11398 15026 11450
rect 15026 11398 15052 11450
rect 14756 11396 14812 11398
rect 14836 11396 14892 11398
rect 14916 11396 14972 11398
rect 14996 11396 15052 11398
rect 14756 10362 14812 10364
rect 14836 10362 14892 10364
rect 14916 10362 14972 10364
rect 14996 10362 15052 10364
rect 14756 10310 14782 10362
rect 14782 10310 14812 10362
rect 14836 10310 14846 10362
rect 14846 10310 14892 10362
rect 14916 10310 14962 10362
rect 14962 10310 14972 10362
rect 14996 10310 15026 10362
rect 15026 10310 15052 10362
rect 14756 10308 14812 10310
rect 14836 10308 14892 10310
rect 14916 10308 14972 10310
rect 14996 10308 15052 10310
rect 14756 9274 14812 9276
rect 14836 9274 14892 9276
rect 14916 9274 14972 9276
rect 14996 9274 15052 9276
rect 14756 9222 14782 9274
rect 14782 9222 14812 9274
rect 14836 9222 14846 9274
rect 14846 9222 14892 9274
rect 14916 9222 14962 9274
rect 14962 9222 14972 9274
rect 14996 9222 15026 9274
rect 15026 9222 15052 9274
rect 14756 9220 14812 9222
rect 14836 9220 14892 9222
rect 14916 9220 14972 9222
rect 14996 9220 15052 9222
rect 16486 18828 16542 18864
rect 16486 18808 16488 18828
rect 16488 18808 16540 18828
rect 16540 18808 16542 18828
rect 18206 21786 18262 21788
rect 18286 21786 18342 21788
rect 18366 21786 18422 21788
rect 18446 21786 18502 21788
rect 18206 21734 18232 21786
rect 18232 21734 18262 21786
rect 18286 21734 18296 21786
rect 18296 21734 18342 21786
rect 18366 21734 18412 21786
rect 18412 21734 18422 21786
rect 18446 21734 18476 21786
rect 18476 21734 18502 21786
rect 18206 21732 18262 21734
rect 18286 21732 18342 21734
rect 18366 21732 18422 21734
rect 18446 21732 18502 21734
rect 18206 20698 18262 20700
rect 18286 20698 18342 20700
rect 18366 20698 18422 20700
rect 18446 20698 18502 20700
rect 18206 20646 18232 20698
rect 18232 20646 18262 20698
rect 18286 20646 18296 20698
rect 18296 20646 18342 20698
rect 18366 20646 18412 20698
rect 18412 20646 18422 20698
rect 18446 20646 18476 20698
rect 18476 20646 18502 20698
rect 18206 20644 18262 20646
rect 18286 20644 18342 20646
rect 18366 20644 18422 20646
rect 18446 20644 18502 20646
rect 18206 19610 18262 19612
rect 18286 19610 18342 19612
rect 18366 19610 18422 19612
rect 18446 19610 18502 19612
rect 18206 19558 18232 19610
rect 18232 19558 18262 19610
rect 18286 19558 18296 19610
rect 18296 19558 18342 19610
rect 18366 19558 18412 19610
rect 18412 19558 18422 19610
rect 18446 19558 18476 19610
rect 18476 19558 18502 19610
rect 18206 19556 18262 19558
rect 18286 19556 18342 19558
rect 18366 19556 18422 19558
rect 18446 19556 18502 19558
rect 18418 18808 18474 18864
rect 18206 18522 18262 18524
rect 18286 18522 18342 18524
rect 18366 18522 18422 18524
rect 18446 18522 18502 18524
rect 18206 18470 18232 18522
rect 18232 18470 18262 18522
rect 18286 18470 18296 18522
rect 18296 18470 18342 18522
rect 18366 18470 18412 18522
rect 18412 18470 18422 18522
rect 18446 18470 18476 18522
rect 18476 18470 18502 18522
rect 18206 18468 18262 18470
rect 18286 18468 18342 18470
rect 18366 18468 18422 18470
rect 18446 18468 18502 18470
rect 18206 17434 18262 17436
rect 18286 17434 18342 17436
rect 18366 17434 18422 17436
rect 18446 17434 18502 17436
rect 18206 17382 18232 17434
rect 18232 17382 18262 17434
rect 18286 17382 18296 17434
rect 18296 17382 18342 17434
rect 18366 17382 18412 17434
rect 18412 17382 18422 17434
rect 18446 17382 18476 17434
rect 18476 17382 18502 17434
rect 18206 17380 18262 17382
rect 18286 17380 18342 17382
rect 18366 17380 18422 17382
rect 18446 17380 18502 17382
rect 18206 16346 18262 16348
rect 18286 16346 18342 16348
rect 18366 16346 18422 16348
rect 18446 16346 18502 16348
rect 18206 16294 18232 16346
rect 18232 16294 18262 16346
rect 18286 16294 18296 16346
rect 18296 16294 18342 16346
rect 18366 16294 18412 16346
rect 18412 16294 18422 16346
rect 18446 16294 18476 16346
rect 18476 16294 18502 16346
rect 18206 16292 18262 16294
rect 18286 16292 18342 16294
rect 18366 16292 18422 16294
rect 18446 16292 18502 16294
rect 18206 15258 18262 15260
rect 18286 15258 18342 15260
rect 18366 15258 18422 15260
rect 18446 15258 18502 15260
rect 18206 15206 18232 15258
rect 18232 15206 18262 15258
rect 18286 15206 18296 15258
rect 18296 15206 18342 15258
rect 18366 15206 18412 15258
rect 18412 15206 18422 15258
rect 18446 15206 18476 15258
rect 18476 15206 18502 15258
rect 18206 15204 18262 15206
rect 18286 15204 18342 15206
rect 18366 15204 18422 15206
rect 18446 15204 18502 15206
rect 18206 14170 18262 14172
rect 18286 14170 18342 14172
rect 18366 14170 18422 14172
rect 18446 14170 18502 14172
rect 18206 14118 18232 14170
rect 18232 14118 18262 14170
rect 18286 14118 18296 14170
rect 18296 14118 18342 14170
rect 18366 14118 18412 14170
rect 18412 14118 18422 14170
rect 18446 14118 18476 14170
rect 18476 14118 18502 14170
rect 18206 14116 18262 14118
rect 18286 14116 18342 14118
rect 18366 14116 18422 14118
rect 18446 14116 18502 14118
rect 18206 13082 18262 13084
rect 18286 13082 18342 13084
rect 18366 13082 18422 13084
rect 18446 13082 18502 13084
rect 18206 13030 18232 13082
rect 18232 13030 18262 13082
rect 18286 13030 18296 13082
rect 18296 13030 18342 13082
rect 18366 13030 18412 13082
rect 18412 13030 18422 13082
rect 18446 13030 18476 13082
rect 18476 13030 18502 13082
rect 18206 13028 18262 13030
rect 18286 13028 18342 13030
rect 18366 13028 18422 13030
rect 18446 13028 18502 13030
rect 18206 11994 18262 11996
rect 18286 11994 18342 11996
rect 18366 11994 18422 11996
rect 18446 11994 18502 11996
rect 18206 11942 18232 11994
rect 18232 11942 18262 11994
rect 18286 11942 18296 11994
rect 18296 11942 18342 11994
rect 18366 11942 18412 11994
rect 18412 11942 18422 11994
rect 18446 11942 18476 11994
rect 18476 11942 18502 11994
rect 18206 11940 18262 11942
rect 18286 11940 18342 11942
rect 18366 11940 18422 11942
rect 18446 11940 18502 11942
rect 18206 10906 18262 10908
rect 18286 10906 18342 10908
rect 18366 10906 18422 10908
rect 18446 10906 18502 10908
rect 18206 10854 18232 10906
rect 18232 10854 18262 10906
rect 18286 10854 18296 10906
rect 18296 10854 18342 10906
rect 18366 10854 18412 10906
rect 18412 10854 18422 10906
rect 18446 10854 18476 10906
rect 18476 10854 18502 10906
rect 18206 10852 18262 10854
rect 18286 10852 18342 10854
rect 18366 10852 18422 10854
rect 18446 10852 18502 10854
rect 14756 8186 14812 8188
rect 14836 8186 14892 8188
rect 14916 8186 14972 8188
rect 14996 8186 15052 8188
rect 14756 8134 14782 8186
rect 14782 8134 14812 8186
rect 14836 8134 14846 8186
rect 14846 8134 14892 8186
rect 14916 8134 14962 8186
rect 14962 8134 14972 8186
rect 14996 8134 15026 8186
rect 15026 8134 15052 8186
rect 14756 8132 14812 8134
rect 14836 8132 14892 8134
rect 14916 8132 14972 8134
rect 14996 8132 15052 8134
rect 14756 7098 14812 7100
rect 14836 7098 14892 7100
rect 14916 7098 14972 7100
rect 14996 7098 15052 7100
rect 14756 7046 14782 7098
rect 14782 7046 14812 7098
rect 14836 7046 14846 7098
rect 14846 7046 14892 7098
rect 14916 7046 14962 7098
rect 14962 7046 14972 7098
rect 14996 7046 15026 7098
rect 15026 7046 15052 7098
rect 14756 7044 14812 7046
rect 14836 7044 14892 7046
rect 14916 7044 14972 7046
rect 14996 7044 15052 7046
rect 14756 6010 14812 6012
rect 14836 6010 14892 6012
rect 14916 6010 14972 6012
rect 14996 6010 15052 6012
rect 14756 5958 14782 6010
rect 14782 5958 14812 6010
rect 14836 5958 14846 6010
rect 14846 5958 14892 6010
rect 14916 5958 14962 6010
rect 14962 5958 14972 6010
rect 14996 5958 15026 6010
rect 15026 5958 15052 6010
rect 14756 5956 14812 5958
rect 14836 5956 14892 5958
rect 14916 5956 14972 5958
rect 14996 5956 15052 5958
rect 18206 9818 18262 9820
rect 18286 9818 18342 9820
rect 18366 9818 18422 9820
rect 18446 9818 18502 9820
rect 18206 9766 18232 9818
rect 18232 9766 18262 9818
rect 18286 9766 18296 9818
rect 18296 9766 18342 9818
rect 18366 9766 18412 9818
rect 18412 9766 18422 9818
rect 18446 9766 18476 9818
rect 18476 9766 18502 9818
rect 18206 9764 18262 9766
rect 18286 9764 18342 9766
rect 18366 9764 18422 9766
rect 18446 9764 18502 9766
rect 18206 8730 18262 8732
rect 18286 8730 18342 8732
rect 18366 8730 18422 8732
rect 18446 8730 18502 8732
rect 18206 8678 18232 8730
rect 18232 8678 18262 8730
rect 18286 8678 18296 8730
rect 18296 8678 18342 8730
rect 18366 8678 18412 8730
rect 18412 8678 18422 8730
rect 18446 8678 18476 8730
rect 18476 8678 18502 8730
rect 18206 8676 18262 8678
rect 18286 8676 18342 8678
rect 18366 8676 18422 8678
rect 18446 8676 18502 8678
rect 18206 7642 18262 7644
rect 18286 7642 18342 7644
rect 18366 7642 18422 7644
rect 18446 7642 18502 7644
rect 18206 7590 18232 7642
rect 18232 7590 18262 7642
rect 18286 7590 18296 7642
rect 18296 7590 18342 7642
rect 18366 7590 18412 7642
rect 18412 7590 18422 7642
rect 18446 7590 18476 7642
rect 18476 7590 18502 7642
rect 18206 7588 18262 7590
rect 18286 7588 18342 7590
rect 18366 7588 18422 7590
rect 18446 7588 18502 7590
rect 18206 6554 18262 6556
rect 18286 6554 18342 6556
rect 18366 6554 18422 6556
rect 18446 6554 18502 6556
rect 18206 6502 18232 6554
rect 18232 6502 18262 6554
rect 18286 6502 18296 6554
rect 18296 6502 18342 6554
rect 18366 6502 18412 6554
rect 18412 6502 18422 6554
rect 18446 6502 18476 6554
rect 18476 6502 18502 6554
rect 18206 6500 18262 6502
rect 18286 6500 18342 6502
rect 18366 6500 18422 6502
rect 18446 6500 18502 6502
rect 18206 5466 18262 5468
rect 18286 5466 18342 5468
rect 18366 5466 18422 5468
rect 18446 5466 18502 5468
rect 18206 5414 18232 5466
rect 18232 5414 18262 5466
rect 18286 5414 18296 5466
rect 18296 5414 18342 5466
rect 18366 5414 18412 5466
rect 18412 5414 18422 5466
rect 18446 5414 18476 5466
rect 18476 5414 18502 5466
rect 18206 5412 18262 5414
rect 18286 5412 18342 5414
rect 18366 5412 18422 5414
rect 18446 5412 18502 5414
rect 14756 4922 14812 4924
rect 14836 4922 14892 4924
rect 14916 4922 14972 4924
rect 14996 4922 15052 4924
rect 14756 4870 14782 4922
rect 14782 4870 14812 4922
rect 14836 4870 14846 4922
rect 14846 4870 14892 4922
rect 14916 4870 14962 4922
rect 14962 4870 14972 4922
rect 14996 4870 15026 4922
rect 15026 4870 15052 4922
rect 14756 4868 14812 4870
rect 14836 4868 14892 4870
rect 14916 4868 14972 4870
rect 14996 4868 15052 4870
rect 14756 3834 14812 3836
rect 14836 3834 14892 3836
rect 14916 3834 14972 3836
rect 14996 3834 15052 3836
rect 14756 3782 14782 3834
rect 14782 3782 14812 3834
rect 14836 3782 14846 3834
rect 14846 3782 14892 3834
rect 14916 3782 14962 3834
rect 14962 3782 14972 3834
rect 14996 3782 15026 3834
rect 15026 3782 15052 3834
rect 14756 3780 14812 3782
rect 14836 3780 14892 3782
rect 14916 3780 14972 3782
rect 14996 3780 15052 3782
rect 4406 2202 4462 2204
rect 4486 2202 4542 2204
rect 4566 2202 4622 2204
rect 4646 2202 4702 2204
rect 4406 2150 4432 2202
rect 4432 2150 4462 2202
rect 4486 2150 4496 2202
rect 4496 2150 4542 2202
rect 4566 2150 4612 2202
rect 4612 2150 4622 2202
rect 4646 2150 4676 2202
rect 4676 2150 4702 2202
rect 4406 2148 4462 2150
rect 4486 2148 4542 2150
rect 4566 2148 4622 2150
rect 4646 2148 4702 2150
rect 11306 2202 11362 2204
rect 11386 2202 11442 2204
rect 11466 2202 11522 2204
rect 11546 2202 11602 2204
rect 11306 2150 11332 2202
rect 11332 2150 11362 2202
rect 11386 2150 11396 2202
rect 11396 2150 11442 2202
rect 11466 2150 11512 2202
rect 11512 2150 11522 2202
rect 11546 2150 11576 2202
rect 11576 2150 11602 2202
rect 11306 2148 11362 2150
rect 11386 2148 11442 2150
rect 11466 2148 11522 2150
rect 11546 2148 11602 2150
rect 14756 2746 14812 2748
rect 14836 2746 14892 2748
rect 14916 2746 14972 2748
rect 14996 2746 15052 2748
rect 14756 2694 14782 2746
rect 14782 2694 14812 2746
rect 14836 2694 14846 2746
rect 14846 2694 14892 2746
rect 14916 2694 14962 2746
rect 14962 2694 14972 2746
rect 14996 2694 15026 2746
rect 15026 2694 15052 2746
rect 14756 2692 14812 2694
rect 14836 2692 14892 2694
rect 14916 2692 14972 2694
rect 14996 2692 15052 2694
rect 18206 4378 18262 4380
rect 18286 4378 18342 4380
rect 18366 4378 18422 4380
rect 18446 4378 18502 4380
rect 18206 4326 18232 4378
rect 18232 4326 18262 4378
rect 18286 4326 18296 4378
rect 18296 4326 18342 4378
rect 18366 4326 18412 4378
rect 18412 4326 18422 4378
rect 18446 4326 18476 4378
rect 18476 4326 18502 4378
rect 18206 4324 18262 4326
rect 18286 4324 18342 4326
rect 18366 4324 18422 4326
rect 18446 4324 18502 4326
rect 18206 3290 18262 3292
rect 18286 3290 18342 3292
rect 18366 3290 18422 3292
rect 18446 3290 18502 3292
rect 18206 3238 18232 3290
rect 18232 3238 18262 3290
rect 18286 3238 18296 3290
rect 18296 3238 18342 3290
rect 18366 3238 18412 3290
rect 18412 3238 18422 3290
rect 18446 3238 18476 3290
rect 18476 3238 18502 3290
rect 18206 3236 18262 3238
rect 18286 3236 18342 3238
rect 18366 3236 18422 3238
rect 18446 3236 18502 3238
rect 21362 20440 21418 20496
rect 21454 17740 21510 17776
rect 21454 17720 21456 17740
rect 21456 17720 21508 17740
rect 21508 17720 21510 17740
rect 21454 15680 21510 15736
rect 21454 12960 21510 13016
rect 21454 10240 21510 10296
rect 21454 8200 21510 8256
rect 21454 5480 21510 5536
rect 21454 2760 21510 2816
rect 18206 2202 18262 2204
rect 18286 2202 18342 2204
rect 18366 2202 18422 2204
rect 18446 2202 18502 2204
rect 18206 2150 18232 2202
rect 18232 2150 18262 2202
rect 18286 2150 18296 2202
rect 18296 2150 18342 2202
rect 18366 2150 18412 2202
rect 18412 2150 18422 2202
rect 18446 2150 18476 2202
rect 18476 2150 18502 2202
rect 18206 2148 18262 2150
rect 18286 2148 18342 2150
rect 18366 2148 18422 2150
rect 18446 2148 18502 2150
<< metal3 >>
rect 0 23218 800 23248
rect 1485 23218 1551 23221
rect 0 23216 1551 23218
rect 0 23160 1490 23216
rect 1546 23160 1551 23216
rect 0 23158 1551 23160
rect 0 23128 800 23158
rect 1485 23155 1551 23158
rect 21081 23218 21147 23221
rect 22179 23218 22979 23248
rect 21081 23216 22979 23218
rect 21081 23160 21086 23216
rect 21142 23160 22979 23216
rect 21081 23158 22979 23160
rect 21081 23155 21147 23158
rect 22179 23128 22979 23158
rect 4394 22880 4714 22881
rect 4394 22816 4402 22880
rect 4466 22816 4482 22880
rect 4546 22816 4562 22880
rect 4626 22816 4642 22880
rect 4706 22816 4714 22880
rect 4394 22815 4714 22816
rect 11294 22880 11614 22881
rect 11294 22816 11302 22880
rect 11366 22816 11382 22880
rect 11446 22816 11462 22880
rect 11526 22816 11542 22880
rect 11606 22816 11614 22880
rect 11294 22815 11614 22816
rect 18194 22880 18514 22881
rect 18194 22816 18202 22880
rect 18266 22816 18282 22880
rect 18346 22816 18362 22880
rect 18426 22816 18442 22880
rect 18506 22816 18514 22880
rect 18194 22815 18514 22816
rect 7844 22336 8164 22337
rect 7844 22272 7852 22336
rect 7916 22272 7932 22336
rect 7996 22272 8012 22336
rect 8076 22272 8092 22336
rect 8156 22272 8164 22336
rect 7844 22271 8164 22272
rect 14744 22336 15064 22337
rect 14744 22272 14752 22336
rect 14816 22272 14832 22336
rect 14896 22272 14912 22336
rect 14976 22272 14992 22336
rect 15056 22272 15064 22336
rect 14744 22271 15064 22272
rect 4394 21792 4714 21793
rect 4394 21728 4402 21792
rect 4466 21728 4482 21792
rect 4546 21728 4562 21792
rect 4626 21728 4642 21792
rect 4706 21728 4714 21792
rect 4394 21727 4714 21728
rect 11294 21792 11614 21793
rect 11294 21728 11302 21792
rect 11366 21728 11382 21792
rect 11446 21728 11462 21792
rect 11526 21728 11542 21792
rect 11606 21728 11614 21792
rect 11294 21727 11614 21728
rect 18194 21792 18514 21793
rect 18194 21728 18202 21792
rect 18266 21728 18282 21792
rect 18346 21728 18362 21792
rect 18426 21728 18442 21792
rect 18506 21728 18514 21792
rect 18194 21727 18514 21728
rect 7844 21248 8164 21249
rect 7844 21184 7852 21248
rect 7916 21184 7932 21248
rect 7996 21184 8012 21248
rect 8076 21184 8092 21248
rect 8156 21184 8164 21248
rect 7844 21183 8164 21184
rect 14744 21248 15064 21249
rect 14744 21184 14752 21248
rect 14816 21184 14832 21248
rect 14896 21184 14912 21248
rect 14976 21184 14992 21248
rect 15056 21184 15064 21248
rect 14744 21183 15064 21184
rect 4394 20704 4714 20705
rect 4394 20640 4402 20704
rect 4466 20640 4482 20704
rect 4546 20640 4562 20704
rect 4626 20640 4642 20704
rect 4706 20640 4714 20704
rect 4394 20639 4714 20640
rect 11294 20704 11614 20705
rect 11294 20640 11302 20704
rect 11366 20640 11382 20704
rect 11446 20640 11462 20704
rect 11526 20640 11542 20704
rect 11606 20640 11614 20704
rect 11294 20639 11614 20640
rect 18194 20704 18514 20705
rect 18194 20640 18202 20704
rect 18266 20640 18282 20704
rect 18346 20640 18362 20704
rect 18426 20640 18442 20704
rect 18506 20640 18514 20704
rect 18194 20639 18514 20640
rect 0 20498 800 20528
rect 1393 20498 1459 20501
rect 0 20496 1459 20498
rect 0 20440 1398 20496
rect 1454 20440 1459 20496
rect 0 20438 1459 20440
rect 0 20408 800 20438
rect 1393 20435 1459 20438
rect 21357 20498 21423 20501
rect 22179 20498 22979 20528
rect 21357 20496 22979 20498
rect 21357 20440 21362 20496
rect 21418 20440 22979 20496
rect 21357 20438 22979 20440
rect 21357 20435 21423 20438
rect 22179 20408 22979 20438
rect 7844 20160 8164 20161
rect 7844 20096 7852 20160
rect 7916 20096 7932 20160
rect 7996 20096 8012 20160
rect 8076 20096 8092 20160
rect 8156 20096 8164 20160
rect 7844 20095 8164 20096
rect 14744 20160 15064 20161
rect 14744 20096 14752 20160
rect 14816 20096 14832 20160
rect 14896 20096 14912 20160
rect 14976 20096 14992 20160
rect 15056 20096 15064 20160
rect 14744 20095 15064 20096
rect 4394 19616 4714 19617
rect 4394 19552 4402 19616
rect 4466 19552 4482 19616
rect 4546 19552 4562 19616
rect 4626 19552 4642 19616
rect 4706 19552 4714 19616
rect 4394 19551 4714 19552
rect 11294 19616 11614 19617
rect 11294 19552 11302 19616
rect 11366 19552 11382 19616
rect 11446 19552 11462 19616
rect 11526 19552 11542 19616
rect 11606 19552 11614 19616
rect 11294 19551 11614 19552
rect 18194 19616 18514 19617
rect 18194 19552 18202 19616
rect 18266 19552 18282 19616
rect 18346 19552 18362 19616
rect 18426 19552 18442 19616
rect 18506 19552 18514 19616
rect 18194 19551 18514 19552
rect 7557 19274 7623 19277
rect 8293 19274 8359 19277
rect 8569 19274 8635 19277
rect 7557 19272 8635 19274
rect 7557 19216 7562 19272
rect 7618 19216 8298 19272
rect 8354 19216 8574 19272
rect 8630 19216 8635 19272
rect 7557 19214 8635 19216
rect 7557 19211 7623 19214
rect 8293 19211 8359 19214
rect 8569 19211 8635 19214
rect 7844 19072 8164 19073
rect 7844 19008 7852 19072
rect 7916 19008 7932 19072
rect 7996 19008 8012 19072
rect 8076 19008 8092 19072
rect 8156 19008 8164 19072
rect 7844 19007 8164 19008
rect 14744 19072 15064 19073
rect 14744 19008 14752 19072
rect 14816 19008 14832 19072
rect 14896 19008 14912 19072
rect 14976 19008 14992 19072
rect 15056 19008 15064 19072
rect 14744 19007 15064 19008
rect 16481 18866 16547 18869
rect 18413 18866 18479 18869
rect 16481 18864 18479 18866
rect 16481 18808 16486 18864
rect 16542 18808 18418 18864
rect 18474 18808 18479 18864
rect 16481 18806 18479 18808
rect 16481 18803 16547 18806
rect 18413 18803 18479 18806
rect 4394 18528 4714 18529
rect 4394 18464 4402 18528
rect 4466 18464 4482 18528
rect 4546 18464 4562 18528
rect 4626 18464 4642 18528
rect 4706 18464 4714 18528
rect 4394 18463 4714 18464
rect 11294 18528 11614 18529
rect 11294 18464 11302 18528
rect 11366 18464 11382 18528
rect 11446 18464 11462 18528
rect 11526 18464 11542 18528
rect 11606 18464 11614 18528
rect 11294 18463 11614 18464
rect 18194 18528 18514 18529
rect 18194 18464 18202 18528
rect 18266 18464 18282 18528
rect 18346 18464 18362 18528
rect 18426 18464 18442 18528
rect 18506 18464 18514 18528
rect 18194 18463 18514 18464
rect 7844 17984 8164 17985
rect 7844 17920 7852 17984
rect 7916 17920 7932 17984
rect 7996 17920 8012 17984
rect 8076 17920 8092 17984
rect 8156 17920 8164 17984
rect 7844 17919 8164 17920
rect 14744 17984 15064 17985
rect 14744 17920 14752 17984
rect 14816 17920 14832 17984
rect 14896 17920 14912 17984
rect 14976 17920 14992 17984
rect 15056 17920 15064 17984
rect 14744 17919 15064 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 21449 17778 21515 17781
rect 22179 17778 22979 17808
rect 21449 17776 22979 17778
rect 21449 17720 21454 17776
rect 21510 17720 22979 17776
rect 21449 17718 22979 17720
rect 21449 17715 21515 17718
rect 22179 17688 22979 17718
rect 4394 17440 4714 17441
rect 4394 17376 4402 17440
rect 4466 17376 4482 17440
rect 4546 17376 4562 17440
rect 4626 17376 4642 17440
rect 4706 17376 4714 17440
rect 4394 17375 4714 17376
rect 11294 17440 11614 17441
rect 11294 17376 11302 17440
rect 11366 17376 11382 17440
rect 11446 17376 11462 17440
rect 11526 17376 11542 17440
rect 11606 17376 11614 17440
rect 11294 17375 11614 17376
rect 18194 17440 18514 17441
rect 18194 17376 18202 17440
rect 18266 17376 18282 17440
rect 18346 17376 18362 17440
rect 18426 17376 18442 17440
rect 18506 17376 18514 17440
rect 18194 17375 18514 17376
rect 7844 16896 8164 16897
rect 7844 16832 7852 16896
rect 7916 16832 7932 16896
rect 7996 16832 8012 16896
rect 8076 16832 8092 16896
rect 8156 16832 8164 16896
rect 7844 16831 8164 16832
rect 14744 16896 15064 16897
rect 14744 16832 14752 16896
rect 14816 16832 14832 16896
rect 14896 16832 14912 16896
rect 14976 16832 14992 16896
rect 15056 16832 15064 16896
rect 14744 16831 15064 16832
rect 4394 16352 4714 16353
rect 4394 16288 4402 16352
rect 4466 16288 4482 16352
rect 4546 16288 4562 16352
rect 4626 16288 4642 16352
rect 4706 16288 4714 16352
rect 4394 16287 4714 16288
rect 11294 16352 11614 16353
rect 11294 16288 11302 16352
rect 11366 16288 11382 16352
rect 11446 16288 11462 16352
rect 11526 16288 11542 16352
rect 11606 16288 11614 16352
rect 11294 16287 11614 16288
rect 18194 16352 18514 16353
rect 18194 16288 18202 16352
rect 18266 16288 18282 16352
rect 18346 16288 18362 16352
rect 18426 16288 18442 16352
rect 18506 16288 18514 16352
rect 18194 16287 18514 16288
rect 7844 15808 8164 15809
rect 0 15738 800 15768
rect 7844 15744 7852 15808
rect 7916 15744 7932 15808
rect 7996 15744 8012 15808
rect 8076 15744 8092 15808
rect 8156 15744 8164 15808
rect 7844 15743 8164 15744
rect 14744 15808 15064 15809
rect 14744 15744 14752 15808
rect 14816 15744 14832 15808
rect 14896 15744 14912 15808
rect 14976 15744 14992 15808
rect 15056 15744 15064 15808
rect 14744 15743 15064 15744
rect 1393 15738 1459 15741
rect 0 15736 1459 15738
rect 0 15680 1398 15736
rect 1454 15680 1459 15736
rect 0 15678 1459 15680
rect 0 15648 800 15678
rect 1393 15675 1459 15678
rect 21449 15738 21515 15741
rect 22179 15738 22979 15768
rect 21449 15736 22979 15738
rect 21449 15680 21454 15736
rect 21510 15680 22979 15736
rect 21449 15678 22979 15680
rect 21449 15675 21515 15678
rect 22179 15648 22979 15678
rect 4394 15264 4714 15265
rect 4394 15200 4402 15264
rect 4466 15200 4482 15264
rect 4546 15200 4562 15264
rect 4626 15200 4642 15264
rect 4706 15200 4714 15264
rect 4394 15199 4714 15200
rect 11294 15264 11614 15265
rect 11294 15200 11302 15264
rect 11366 15200 11382 15264
rect 11446 15200 11462 15264
rect 11526 15200 11542 15264
rect 11606 15200 11614 15264
rect 11294 15199 11614 15200
rect 18194 15264 18514 15265
rect 18194 15200 18202 15264
rect 18266 15200 18282 15264
rect 18346 15200 18362 15264
rect 18426 15200 18442 15264
rect 18506 15200 18514 15264
rect 18194 15199 18514 15200
rect 7844 14720 8164 14721
rect 7844 14656 7852 14720
rect 7916 14656 7932 14720
rect 7996 14656 8012 14720
rect 8076 14656 8092 14720
rect 8156 14656 8164 14720
rect 7844 14655 8164 14656
rect 14744 14720 15064 14721
rect 14744 14656 14752 14720
rect 14816 14656 14832 14720
rect 14896 14656 14912 14720
rect 14976 14656 14992 14720
rect 15056 14656 15064 14720
rect 14744 14655 15064 14656
rect 4394 14176 4714 14177
rect 4394 14112 4402 14176
rect 4466 14112 4482 14176
rect 4546 14112 4562 14176
rect 4626 14112 4642 14176
rect 4706 14112 4714 14176
rect 4394 14111 4714 14112
rect 11294 14176 11614 14177
rect 11294 14112 11302 14176
rect 11366 14112 11382 14176
rect 11446 14112 11462 14176
rect 11526 14112 11542 14176
rect 11606 14112 11614 14176
rect 11294 14111 11614 14112
rect 18194 14176 18514 14177
rect 18194 14112 18202 14176
rect 18266 14112 18282 14176
rect 18346 14112 18362 14176
rect 18426 14112 18442 14176
rect 18506 14112 18514 14176
rect 18194 14111 18514 14112
rect 7844 13632 8164 13633
rect 7844 13568 7852 13632
rect 7916 13568 7932 13632
rect 7996 13568 8012 13632
rect 8076 13568 8092 13632
rect 8156 13568 8164 13632
rect 7844 13567 8164 13568
rect 14744 13632 15064 13633
rect 14744 13568 14752 13632
rect 14816 13568 14832 13632
rect 14896 13568 14912 13632
rect 14976 13568 14992 13632
rect 15056 13568 15064 13632
rect 14744 13567 15064 13568
rect 4394 13088 4714 13089
rect 0 13018 800 13048
rect 4394 13024 4402 13088
rect 4466 13024 4482 13088
rect 4546 13024 4562 13088
rect 4626 13024 4642 13088
rect 4706 13024 4714 13088
rect 4394 13023 4714 13024
rect 11294 13088 11614 13089
rect 11294 13024 11302 13088
rect 11366 13024 11382 13088
rect 11446 13024 11462 13088
rect 11526 13024 11542 13088
rect 11606 13024 11614 13088
rect 11294 13023 11614 13024
rect 18194 13088 18514 13089
rect 18194 13024 18202 13088
rect 18266 13024 18282 13088
rect 18346 13024 18362 13088
rect 18426 13024 18442 13088
rect 18506 13024 18514 13088
rect 18194 13023 18514 13024
rect 1485 13018 1551 13021
rect 0 13016 1551 13018
rect 0 12960 1490 13016
rect 1546 12960 1551 13016
rect 0 12958 1551 12960
rect 0 12928 800 12958
rect 1485 12955 1551 12958
rect 21449 13018 21515 13021
rect 22179 13018 22979 13048
rect 21449 13016 22979 13018
rect 21449 12960 21454 13016
rect 21510 12960 22979 13016
rect 21449 12958 22979 12960
rect 21449 12955 21515 12958
rect 22179 12928 22979 12958
rect 7844 12544 8164 12545
rect 7844 12480 7852 12544
rect 7916 12480 7932 12544
rect 7996 12480 8012 12544
rect 8076 12480 8092 12544
rect 8156 12480 8164 12544
rect 7844 12479 8164 12480
rect 14744 12544 15064 12545
rect 14744 12480 14752 12544
rect 14816 12480 14832 12544
rect 14896 12480 14912 12544
rect 14976 12480 14992 12544
rect 15056 12480 15064 12544
rect 14744 12479 15064 12480
rect 4394 12000 4714 12001
rect 4394 11936 4402 12000
rect 4466 11936 4482 12000
rect 4546 11936 4562 12000
rect 4626 11936 4642 12000
rect 4706 11936 4714 12000
rect 4394 11935 4714 11936
rect 11294 12000 11614 12001
rect 11294 11936 11302 12000
rect 11366 11936 11382 12000
rect 11446 11936 11462 12000
rect 11526 11936 11542 12000
rect 11606 11936 11614 12000
rect 11294 11935 11614 11936
rect 18194 12000 18514 12001
rect 18194 11936 18202 12000
rect 18266 11936 18282 12000
rect 18346 11936 18362 12000
rect 18426 11936 18442 12000
rect 18506 11936 18514 12000
rect 18194 11935 18514 11936
rect 7844 11456 8164 11457
rect 7844 11392 7852 11456
rect 7916 11392 7932 11456
rect 7996 11392 8012 11456
rect 8076 11392 8092 11456
rect 8156 11392 8164 11456
rect 7844 11391 8164 11392
rect 14744 11456 15064 11457
rect 14744 11392 14752 11456
rect 14816 11392 14832 11456
rect 14896 11392 14912 11456
rect 14976 11392 14992 11456
rect 15056 11392 15064 11456
rect 14744 11391 15064 11392
rect 4394 10912 4714 10913
rect 4394 10848 4402 10912
rect 4466 10848 4482 10912
rect 4546 10848 4562 10912
rect 4626 10848 4642 10912
rect 4706 10848 4714 10912
rect 4394 10847 4714 10848
rect 11294 10912 11614 10913
rect 11294 10848 11302 10912
rect 11366 10848 11382 10912
rect 11446 10848 11462 10912
rect 11526 10848 11542 10912
rect 11606 10848 11614 10912
rect 11294 10847 11614 10848
rect 18194 10912 18514 10913
rect 18194 10848 18202 10912
rect 18266 10848 18282 10912
rect 18346 10848 18362 10912
rect 18426 10848 18442 10912
rect 18506 10848 18514 10912
rect 18194 10847 18514 10848
rect 7844 10368 8164 10369
rect 0 10298 800 10328
rect 7844 10304 7852 10368
rect 7916 10304 7932 10368
rect 7996 10304 8012 10368
rect 8076 10304 8092 10368
rect 8156 10304 8164 10368
rect 7844 10303 8164 10304
rect 14744 10368 15064 10369
rect 14744 10304 14752 10368
rect 14816 10304 14832 10368
rect 14896 10304 14912 10368
rect 14976 10304 14992 10368
rect 15056 10304 15064 10368
rect 14744 10303 15064 10304
rect 1485 10298 1551 10301
rect 0 10296 1551 10298
rect 0 10240 1490 10296
rect 1546 10240 1551 10296
rect 0 10238 1551 10240
rect 0 10208 800 10238
rect 1485 10235 1551 10238
rect 21449 10298 21515 10301
rect 22179 10298 22979 10328
rect 21449 10296 22979 10298
rect 21449 10240 21454 10296
rect 21510 10240 22979 10296
rect 21449 10238 22979 10240
rect 21449 10235 21515 10238
rect 22179 10208 22979 10238
rect 4394 9824 4714 9825
rect 4394 9760 4402 9824
rect 4466 9760 4482 9824
rect 4546 9760 4562 9824
rect 4626 9760 4642 9824
rect 4706 9760 4714 9824
rect 4394 9759 4714 9760
rect 11294 9824 11614 9825
rect 11294 9760 11302 9824
rect 11366 9760 11382 9824
rect 11446 9760 11462 9824
rect 11526 9760 11542 9824
rect 11606 9760 11614 9824
rect 11294 9759 11614 9760
rect 18194 9824 18514 9825
rect 18194 9760 18202 9824
rect 18266 9760 18282 9824
rect 18346 9760 18362 9824
rect 18426 9760 18442 9824
rect 18506 9760 18514 9824
rect 18194 9759 18514 9760
rect 7844 9280 8164 9281
rect 7844 9216 7852 9280
rect 7916 9216 7932 9280
rect 7996 9216 8012 9280
rect 8076 9216 8092 9280
rect 8156 9216 8164 9280
rect 7844 9215 8164 9216
rect 14744 9280 15064 9281
rect 14744 9216 14752 9280
rect 14816 9216 14832 9280
rect 14896 9216 14912 9280
rect 14976 9216 14992 9280
rect 15056 9216 15064 9280
rect 14744 9215 15064 9216
rect 4394 8736 4714 8737
rect 4394 8672 4402 8736
rect 4466 8672 4482 8736
rect 4546 8672 4562 8736
rect 4626 8672 4642 8736
rect 4706 8672 4714 8736
rect 4394 8671 4714 8672
rect 11294 8736 11614 8737
rect 11294 8672 11302 8736
rect 11366 8672 11382 8736
rect 11446 8672 11462 8736
rect 11526 8672 11542 8736
rect 11606 8672 11614 8736
rect 11294 8671 11614 8672
rect 18194 8736 18514 8737
rect 18194 8672 18202 8736
rect 18266 8672 18282 8736
rect 18346 8672 18362 8736
rect 18426 8672 18442 8736
rect 18506 8672 18514 8736
rect 18194 8671 18514 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 21449 8258 21515 8261
rect 22179 8258 22979 8288
rect 21449 8256 22979 8258
rect 21449 8200 21454 8256
rect 21510 8200 22979 8256
rect 21449 8198 22979 8200
rect 21449 8195 21515 8198
rect 7844 8192 8164 8193
rect 7844 8128 7852 8192
rect 7916 8128 7932 8192
rect 7996 8128 8012 8192
rect 8076 8128 8092 8192
rect 8156 8128 8164 8192
rect 7844 8127 8164 8128
rect 14744 8192 15064 8193
rect 14744 8128 14752 8192
rect 14816 8128 14832 8192
rect 14896 8128 14912 8192
rect 14976 8128 14992 8192
rect 15056 8128 15064 8192
rect 22179 8168 22979 8198
rect 14744 8127 15064 8128
rect 4394 7648 4714 7649
rect 4394 7584 4402 7648
rect 4466 7584 4482 7648
rect 4546 7584 4562 7648
rect 4626 7584 4642 7648
rect 4706 7584 4714 7648
rect 4394 7583 4714 7584
rect 11294 7648 11614 7649
rect 11294 7584 11302 7648
rect 11366 7584 11382 7648
rect 11446 7584 11462 7648
rect 11526 7584 11542 7648
rect 11606 7584 11614 7648
rect 11294 7583 11614 7584
rect 18194 7648 18514 7649
rect 18194 7584 18202 7648
rect 18266 7584 18282 7648
rect 18346 7584 18362 7648
rect 18426 7584 18442 7648
rect 18506 7584 18514 7648
rect 18194 7583 18514 7584
rect 7844 7104 8164 7105
rect 7844 7040 7852 7104
rect 7916 7040 7932 7104
rect 7996 7040 8012 7104
rect 8076 7040 8092 7104
rect 8156 7040 8164 7104
rect 7844 7039 8164 7040
rect 14744 7104 15064 7105
rect 14744 7040 14752 7104
rect 14816 7040 14832 7104
rect 14896 7040 14912 7104
rect 14976 7040 14992 7104
rect 15056 7040 15064 7104
rect 14744 7039 15064 7040
rect 4394 6560 4714 6561
rect 4394 6496 4402 6560
rect 4466 6496 4482 6560
rect 4546 6496 4562 6560
rect 4626 6496 4642 6560
rect 4706 6496 4714 6560
rect 4394 6495 4714 6496
rect 11294 6560 11614 6561
rect 11294 6496 11302 6560
rect 11366 6496 11382 6560
rect 11446 6496 11462 6560
rect 11526 6496 11542 6560
rect 11606 6496 11614 6560
rect 11294 6495 11614 6496
rect 18194 6560 18514 6561
rect 18194 6496 18202 6560
rect 18266 6496 18282 6560
rect 18346 6496 18362 6560
rect 18426 6496 18442 6560
rect 18506 6496 18514 6560
rect 18194 6495 18514 6496
rect 7844 6016 8164 6017
rect 7844 5952 7852 6016
rect 7916 5952 7932 6016
rect 7996 5952 8012 6016
rect 8076 5952 8092 6016
rect 8156 5952 8164 6016
rect 7844 5951 8164 5952
rect 14744 6016 15064 6017
rect 14744 5952 14752 6016
rect 14816 5952 14832 6016
rect 14896 5952 14912 6016
rect 14976 5952 14992 6016
rect 15056 5952 15064 6016
rect 14744 5951 15064 5952
rect 0 5538 800 5568
rect 1485 5538 1551 5541
rect 0 5536 1551 5538
rect 0 5480 1490 5536
rect 1546 5480 1551 5536
rect 0 5478 1551 5480
rect 0 5448 800 5478
rect 1485 5475 1551 5478
rect 21449 5538 21515 5541
rect 22179 5538 22979 5568
rect 21449 5536 22979 5538
rect 21449 5480 21454 5536
rect 21510 5480 22979 5536
rect 21449 5478 22979 5480
rect 21449 5475 21515 5478
rect 4394 5472 4714 5473
rect 4394 5408 4402 5472
rect 4466 5408 4482 5472
rect 4546 5408 4562 5472
rect 4626 5408 4642 5472
rect 4706 5408 4714 5472
rect 4394 5407 4714 5408
rect 11294 5472 11614 5473
rect 11294 5408 11302 5472
rect 11366 5408 11382 5472
rect 11446 5408 11462 5472
rect 11526 5408 11542 5472
rect 11606 5408 11614 5472
rect 11294 5407 11614 5408
rect 18194 5472 18514 5473
rect 18194 5408 18202 5472
rect 18266 5408 18282 5472
rect 18346 5408 18362 5472
rect 18426 5408 18442 5472
rect 18506 5408 18514 5472
rect 22179 5448 22979 5478
rect 18194 5407 18514 5408
rect 7844 4928 8164 4929
rect 7844 4864 7852 4928
rect 7916 4864 7932 4928
rect 7996 4864 8012 4928
rect 8076 4864 8092 4928
rect 8156 4864 8164 4928
rect 7844 4863 8164 4864
rect 14744 4928 15064 4929
rect 14744 4864 14752 4928
rect 14816 4864 14832 4928
rect 14896 4864 14912 4928
rect 14976 4864 14992 4928
rect 15056 4864 15064 4928
rect 14744 4863 15064 4864
rect 4394 4384 4714 4385
rect 4394 4320 4402 4384
rect 4466 4320 4482 4384
rect 4546 4320 4562 4384
rect 4626 4320 4642 4384
rect 4706 4320 4714 4384
rect 4394 4319 4714 4320
rect 11294 4384 11614 4385
rect 11294 4320 11302 4384
rect 11366 4320 11382 4384
rect 11446 4320 11462 4384
rect 11526 4320 11542 4384
rect 11606 4320 11614 4384
rect 11294 4319 11614 4320
rect 18194 4384 18514 4385
rect 18194 4320 18202 4384
rect 18266 4320 18282 4384
rect 18346 4320 18362 4384
rect 18426 4320 18442 4384
rect 18506 4320 18514 4384
rect 18194 4319 18514 4320
rect 7844 3840 8164 3841
rect 7844 3776 7852 3840
rect 7916 3776 7932 3840
rect 7996 3776 8012 3840
rect 8076 3776 8092 3840
rect 8156 3776 8164 3840
rect 7844 3775 8164 3776
rect 14744 3840 15064 3841
rect 14744 3776 14752 3840
rect 14816 3776 14832 3840
rect 14896 3776 14912 3840
rect 14976 3776 14992 3840
rect 15056 3776 15064 3840
rect 14744 3775 15064 3776
rect 4394 3296 4714 3297
rect 4394 3232 4402 3296
rect 4466 3232 4482 3296
rect 4546 3232 4562 3296
rect 4626 3232 4642 3296
rect 4706 3232 4714 3296
rect 4394 3231 4714 3232
rect 11294 3296 11614 3297
rect 11294 3232 11302 3296
rect 11366 3232 11382 3296
rect 11446 3232 11462 3296
rect 11526 3232 11542 3296
rect 11606 3232 11614 3296
rect 11294 3231 11614 3232
rect 18194 3296 18514 3297
rect 18194 3232 18202 3296
rect 18266 3232 18282 3296
rect 18346 3232 18362 3296
rect 18426 3232 18442 3296
rect 18506 3232 18514 3296
rect 18194 3231 18514 3232
rect 0 2818 800 2848
rect 1393 2818 1459 2821
rect 0 2816 1459 2818
rect 0 2760 1398 2816
rect 1454 2760 1459 2816
rect 0 2758 1459 2760
rect 0 2728 800 2758
rect 1393 2755 1459 2758
rect 21449 2818 21515 2821
rect 22179 2818 22979 2848
rect 21449 2816 22979 2818
rect 21449 2760 21454 2816
rect 21510 2760 22979 2816
rect 21449 2758 22979 2760
rect 21449 2755 21515 2758
rect 7844 2752 8164 2753
rect 7844 2688 7852 2752
rect 7916 2688 7932 2752
rect 7996 2688 8012 2752
rect 8076 2688 8092 2752
rect 8156 2688 8164 2752
rect 7844 2687 8164 2688
rect 14744 2752 15064 2753
rect 14744 2688 14752 2752
rect 14816 2688 14832 2752
rect 14896 2688 14912 2752
rect 14976 2688 14992 2752
rect 15056 2688 15064 2752
rect 22179 2728 22979 2758
rect 14744 2687 15064 2688
rect 4394 2208 4714 2209
rect 4394 2144 4402 2208
rect 4466 2144 4482 2208
rect 4546 2144 4562 2208
rect 4626 2144 4642 2208
rect 4706 2144 4714 2208
rect 4394 2143 4714 2144
rect 11294 2208 11614 2209
rect 11294 2144 11302 2208
rect 11366 2144 11382 2208
rect 11446 2144 11462 2208
rect 11526 2144 11542 2208
rect 11606 2144 11614 2208
rect 11294 2143 11614 2144
rect 18194 2208 18514 2209
rect 18194 2144 18202 2208
rect 18266 2144 18282 2208
rect 18346 2144 18362 2208
rect 18426 2144 18442 2208
rect 18506 2144 18514 2208
rect 18194 2143 18514 2144
<< via3 >>
rect 4402 22876 4466 22880
rect 4402 22820 4406 22876
rect 4406 22820 4462 22876
rect 4462 22820 4466 22876
rect 4402 22816 4466 22820
rect 4482 22876 4546 22880
rect 4482 22820 4486 22876
rect 4486 22820 4542 22876
rect 4542 22820 4546 22876
rect 4482 22816 4546 22820
rect 4562 22876 4626 22880
rect 4562 22820 4566 22876
rect 4566 22820 4622 22876
rect 4622 22820 4626 22876
rect 4562 22816 4626 22820
rect 4642 22876 4706 22880
rect 4642 22820 4646 22876
rect 4646 22820 4702 22876
rect 4702 22820 4706 22876
rect 4642 22816 4706 22820
rect 11302 22876 11366 22880
rect 11302 22820 11306 22876
rect 11306 22820 11362 22876
rect 11362 22820 11366 22876
rect 11302 22816 11366 22820
rect 11382 22876 11446 22880
rect 11382 22820 11386 22876
rect 11386 22820 11442 22876
rect 11442 22820 11446 22876
rect 11382 22816 11446 22820
rect 11462 22876 11526 22880
rect 11462 22820 11466 22876
rect 11466 22820 11522 22876
rect 11522 22820 11526 22876
rect 11462 22816 11526 22820
rect 11542 22876 11606 22880
rect 11542 22820 11546 22876
rect 11546 22820 11602 22876
rect 11602 22820 11606 22876
rect 11542 22816 11606 22820
rect 18202 22876 18266 22880
rect 18202 22820 18206 22876
rect 18206 22820 18262 22876
rect 18262 22820 18266 22876
rect 18202 22816 18266 22820
rect 18282 22876 18346 22880
rect 18282 22820 18286 22876
rect 18286 22820 18342 22876
rect 18342 22820 18346 22876
rect 18282 22816 18346 22820
rect 18362 22876 18426 22880
rect 18362 22820 18366 22876
rect 18366 22820 18422 22876
rect 18422 22820 18426 22876
rect 18362 22816 18426 22820
rect 18442 22876 18506 22880
rect 18442 22820 18446 22876
rect 18446 22820 18502 22876
rect 18502 22820 18506 22876
rect 18442 22816 18506 22820
rect 7852 22332 7916 22336
rect 7852 22276 7856 22332
rect 7856 22276 7912 22332
rect 7912 22276 7916 22332
rect 7852 22272 7916 22276
rect 7932 22332 7996 22336
rect 7932 22276 7936 22332
rect 7936 22276 7992 22332
rect 7992 22276 7996 22332
rect 7932 22272 7996 22276
rect 8012 22332 8076 22336
rect 8012 22276 8016 22332
rect 8016 22276 8072 22332
rect 8072 22276 8076 22332
rect 8012 22272 8076 22276
rect 8092 22332 8156 22336
rect 8092 22276 8096 22332
rect 8096 22276 8152 22332
rect 8152 22276 8156 22332
rect 8092 22272 8156 22276
rect 14752 22332 14816 22336
rect 14752 22276 14756 22332
rect 14756 22276 14812 22332
rect 14812 22276 14816 22332
rect 14752 22272 14816 22276
rect 14832 22332 14896 22336
rect 14832 22276 14836 22332
rect 14836 22276 14892 22332
rect 14892 22276 14896 22332
rect 14832 22272 14896 22276
rect 14912 22332 14976 22336
rect 14912 22276 14916 22332
rect 14916 22276 14972 22332
rect 14972 22276 14976 22332
rect 14912 22272 14976 22276
rect 14992 22332 15056 22336
rect 14992 22276 14996 22332
rect 14996 22276 15052 22332
rect 15052 22276 15056 22332
rect 14992 22272 15056 22276
rect 4402 21788 4466 21792
rect 4402 21732 4406 21788
rect 4406 21732 4462 21788
rect 4462 21732 4466 21788
rect 4402 21728 4466 21732
rect 4482 21788 4546 21792
rect 4482 21732 4486 21788
rect 4486 21732 4542 21788
rect 4542 21732 4546 21788
rect 4482 21728 4546 21732
rect 4562 21788 4626 21792
rect 4562 21732 4566 21788
rect 4566 21732 4622 21788
rect 4622 21732 4626 21788
rect 4562 21728 4626 21732
rect 4642 21788 4706 21792
rect 4642 21732 4646 21788
rect 4646 21732 4702 21788
rect 4702 21732 4706 21788
rect 4642 21728 4706 21732
rect 11302 21788 11366 21792
rect 11302 21732 11306 21788
rect 11306 21732 11362 21788
rect 11362 21732 11366 21788
rect 11302 21728 11366 21732
rect 11382 21788 11446 21792
rect 11382 21732 11386 21788
rect 11386 21732 11442 21788
rect 11442 21732 11446 21788
rect 11382 21728 11446 21732
rect 11462 21788 11526 21792
rect 11462 21732 11466 21788
rect 11466 21732 11522 21788
rect 11522 21732 11526 21788
rect 11462 21728 11526 21732
rect 11542 21788 11606 21792
rect 11542 21732 11546 21788
rect 11546 21732 11602 21788
rect 11602 21732 11606 21788
rect 11542 21728 11606 21732
rect 18202 21788 18266 21792
rect 18202 21732 18206 21788
rect 18206 21732 18262 21788
rect 18262 21732 18266 21788
rect 18202 21728 18266 21732
rect 18282 21788 18346 21792
rect 18282 21732 18286 21788
rect 18286 21732 18342 21788
rect 18342 21732 18346 21788
rect 18282 21728 18346 21732
rect 18362 21788 18426 21792
rect 18362 21732 18366 21788
rect 18366 21732 18422 21788
rect 18422 21732 18426 21788
rect 18362 21728 18426 21732
rect 18442 21788 18506 21792
rect 18442 21732 18446 21788
rect 18446 21732 18502 21788
rect 18502 21732 18506 21788
rect 18442 21728 18506 21732
rect 7852 21244 7916 21248
rect 7852 21188 7856 21244
rect 7856 21188 7912 21244
rect 7912 21188 7916 21244
rect 7852 21184 7916 21188
rect 7932 21244 7996 21248
rect 7932 21188 7936 21244
rect 7936 21188 7992 21244
rect 7992 21188 7996 21244
rect 7932 21184 7996 21188
rect 8012 21244 8076 21248
rect 8012 21188 8016 21244
rect 8016 21188 8072 21244
rect 8072 21188 8076 21244
rect 8012 21184 8076 21188
rect 8092 21244 8156 21248
rect 8092 21188 8096 21244
rect 8096 21188 8152 21244
rect 8152 21188 8156 21244
rect 8092 21184 8156 21188
rect 14752 21244 14816 21248
rect 14752 21188 14756 21244
rect 14756 21188 14812 21244
rect 14812 21188 14816 21244
rect 14752 21184 14816 21188
rect 14832 21244 14896 21248
rect 14832 21188 14836 21244
rect 14836 21188 14892 21244
rect 14892 21188 14896 21244
rect 14832 21184 14896 21188
rect 14912 21244 14976 21248
rect 14912 21188 14916 21244
rect 14916 21188 14972 21244
rect 14972 21188 14976 21244
rect 14912 21184 14976 21188
rect 14992 21244 15056 21248
rect 14992 21188 14996 21244
rect 14996 21188 15052 21244
rect 15052 21188 15056 21244
rect 14992 21184 15056 21188
rect 4402 20700 4466 20704
rect 4402 20644 4406 20700
rect 4406 20644 4462 20700
rect 4462 20644 4466 20700
rect 4402 20640 4466 20644
rect 4482 20700 4546 20704
rect 4482 20644 4486 20700
rect 4486 20644 4542 20700
rect 4542 20644 4546 20700
rect 4482 20640 4546 20644
rect 4562 20700 4626 20704
rect 4562 20644 4566 20700
rect 4566 20644 4622 20700
rect 4622 20644 4626 20700
rect 4562 20640 4626 20644
rect 4642 20700 4706 20704
rect 4642 20644 4646 20700
rect 4646 20644 4702 20700
rect 4702 20644 4706 20700
rect 4642 20640 4706 20644
rect 11302 20700 11366 20704
rect 11302 20644 11306 20700
rect 11306 20644 11362 20700
rect 11362 20644 11366 20700
rect 11302 20640 11366 20644
rect 11382 20700 11446 20704
rect 11382 20644 11386 20700
rect 11386 20644 11442 20700
rect 11442 20644 11446 20700
rect 11382 20640 11446 20644
rect 11462 20700 11526 20704
rect 11462 20644 11466 20700
rect 11466 20644 11522 20700
rect 11522 20644 11526 20700
rect 11462 20640 11526 20644
rect 11542 20700 11606 20704
rect 11542 20644 11546 20700
rect 11546 20644 11602 20700
rect 11602 20644 11606 20700
rect 11542 20640 11606 20644
rect 18202 20700 18266 20704
rect 18202 20644 18206 20700
rect 18206 20644 18262 20700
rect 18262 20644 18266 20700
rect 18202 20640 18266 20644
rect 18282 20700 18346 20704
rect 18282 20644 18286 20700
rect 18286 20644 18342 20700
rect 18342 20644 18346 20700
rect 18282 20640 18346 20644
rect 18362 20700 18426 20704
rect 18362 20644 18366 20700
rect 18366 20644 18422 20700
rect 18422 20644 18426 20700
rect 18362 20640 18426 20644
rect 18442 20700 18506 20704
rect 18442 20644 18446 20700
rect 18446 20644 18502 20700
rect 18502 20644 18506 20700
rect 18442 20640 18506 20644
rect 7852 20156 7916 20160
rect 7852 20100 7856 20156
rect 7856 20100 7912 20156
rect 7912 20100 7916 20156
rect 7852 20096 7916 20100
rect 7932 20156 7996 20160
rect 7932 20100 7936 20156
rect 7936 20100 7992 20156
rect 7992 20100 7996 20156
rect 7932 20096 7996 20100
rect 8012 20156 8076 20160
rect 8012 20100 8016 20156
rect 8016 20100 8072 20156
rect 8072 20100 8076 20156
rect 8012 20096 8076 20100
rect 8092 20156 8156 20160
rect 8092 20100 8096 20156
rect 8096 20100 8152 20156
rect 8152 20100 8156 20156
rect 8092 20096 8156 20100
rect 14752 20156 14816 20160
rect 14752 20100 14756 20156
rect 14756 20100 14812 20156
rect 14812 20100 14816 20156
rect 14752 20096 14816 20100
rect 14832 20156 14896 20160
rect 14832 20100 14836 20156
rect 14836 20100 14892 20156
rect 14892 20100 14896 20156
rect 14832 20096 14896 20100
rect 14912 20156 14976 20160
rect 14912 20100 14916 20156
rect 14916 20100 14972 20156
rect 14972 20100 14976 20156
rect 14912 20096 14976 20100
rect 14992 20156 15056 20160
rect 14992 20100 14996 20156
rect 14996 20100 15052 20156
rect 15052 20100 15056 20156
rect 14992 20096 15056 20100
rect 4402 19612 4466 19616
rect 4402 19556 4406 19612
rect 4406 19556 4462 19612
rect 4462 19556 4466 19612
rect 4402 19552 4466 19556
rect 4482 19612 4546 19616
rect 4482 19556 4486 19612
rect 4486 19556 4542 19612
rect 4542 19556 4546 19612
rect 4482 19552 4546 19556
rect 4562 19612 4626 19616
rect 4562 19556 4566 19612
rect 4566 19556 4622 19612
rect 4622 19556 4626 19612
rect 4562 19552 4626 19556
rect 4642 19612 4706 19616
rect 4642 19556 4646 19612
rect 4646 19556 4702 19612
rect 4702 19556 4706 19612
rect 4642 19552 4706 19556
rect 11302 19612 11366 19616
rect 11302 19556 11306 19612
rect 11306 19556 11362 19612
rect 11362 19556 11366 19612
rect 11302 19552 11366 19556
rect 11382 19612 11446 19616
rect 11382 19556 11386 19612
rect 11386 19556 11442 19612
rect 11442 19556 11446 19612
rect 11382 19552 11446 19556
rect 11462 19612 11526 19616
rect 11462 19556 11466 19612
rect 11466 19556 11522 19612
rect 11522 19556 11526 19612
rect 11462 19552 11526 19556
rect 11542 19612 11606 19616
rect 11542 19556 11546 19612
rect 11546 19556 11602 19612
rect 11602 19556 11606 19612
rect 11542 19552 11606 19556
rect 18202 19612 18266 19616
rect 18202 19556 18206 19612
rect 18206 19556 18262 19612
rect 18262 19556 18266 19612
rect 18202 19552 18266 19556
rect 18282 19612 18346 19616
rect 18282 19556 18286 19612
rect 18286 19556 18342 19612
rect 18342 19556 18346 19612
rect 18282 19552 18346 19556
rect 18362 19612 18426 19616
rect 18362 19556 18366 19612
rect 18366 19556 18422 19612
rect 18422 19556 18426 19612
rect 18362 19552 18426 19556
rect 18442 19612 18506 19616
rect 18442 19556 18446 19612
rect 18446 19556 18502 19612
rect 18502 19556 18506 19612
rect 18442 19552 18506 19556
rect 7852 19068 7916 19072
rect 7852 19012 7856 19068
rect 7856 19012 7912 19068
rect 7912 19012 7916 19068
rect 7852 19008 7916 19012
rect 7932 19068 7996 19072
rect 7932 19012 7936 19068
rect 7936 19012 7992 19068
rect 7992 19012 7996 19068
rect 7932 19008 7996 19012
rect 8012 19068 8076 19072
rect 8012 19012 8016 19068
rect 8016 19012 8072 19068
rect 8072 19012 8076 19068
rect 8012 19008 8076 19012
rect 8092 19068 8156 19072
rect 8092 19012 8096 19068
rect 8096 19012 8152 19068
rect 8152 19012 8156 19068
rect 8092 19008 8156 19012
rect 14752 19068 14816 19072
rect 14752 19012 14756 19068
rect 14756 19012 14812 19068
rect 14812 19012 14816 19068
rect 14752 19008 14816 19012
rect 14832 19068 14896 19072
rect 14832 19012 14836 19068
rect 14836 19012 14892 19068
rect 14892 19012 14896 19068
rect 14832 19008 14896 19012
rect 14912 19068 14976 19072
rect 14912 19012 14916 19068
rect 14916 19012 14972 19068
rect 14972 19012 14976 19068
rect 14912 19008 14976 19012
rect 14992 19068 15056 19072
rect 14992 19012 14996 19068
rect 14996 19012 15052 19068
rect 15052 19012 15056 19068
rect 14992 19008 15056 19012
rect 4402 18524 4466 18528
rect 4402 18468 4406 18524
rect 4406 18468 4462 18524
rect 4462 18468 4466 18524
rect 4402 18464 4466 18468
rect 4482 18524 4546 18528
rect 4482 18468 4486 18524
rect 4486 18468 4542 18524
rect 4542 18468 4546 18524
rect 4482 18464 4546 18468
rect 4562 18524 4626 18528
rect 4562 18468 4566 18524
rect 4566 18468 4622 18524
rect 4622 18468 4626 18524
rect 4562 18464 4626 18468
rect 4642 18524 4706 18528
rect 4642 18468 4646 18524
rect 4646 18468 4702 18524
rect 4702 18468 4706 18524
rect 4642 18464 4706 18468
rect 11302 18524 11366 18528
rect 11302 18468 11306 18524
rect 11306 18468 11362 18524
rect 11362 18468 11366 18524
rect 11302 18464 11366 18468
rect 11382 18524 11446 18528
rect 11382 18468 11386 18524
rect 11386 18468 11442 18524
rect 11442 18468 11446 18524
rect 11382 18464 11446 18468
rect 11462 18524 11526 18528
rect 11462 18468 11466 18524
rect 11466 18468 11522 18524
rect 11522 18468 11526 18524
rect 11462 18464 11526 18468
rect 11542 18524 11606 18528
rect 11542 18468 11546 18524
rect 11546 18468 11602 18524
rect 11602 18468 11606 18524
rect 11542 18464 11606 18468
rect 18202 18524 18266 18528
rect 18202 18468 18206 18524
rect 18206 18468 18262 18524
rect 18262 18468 18266 18524
rect 18202 18464 18266 18468
rect 18282 18524 18346 18528
rect 18282 18468 18286 18524
rect 18286 18468 18342 18524
rect 18342 18468 18346 18524
rect 18282 18464 18346 18468
rect 18362 18524 18426 18528
rect 18362 18468 18366 18524
rect 18366 18468 18422 18524
rect 18422 18468 18426 18524
rect 18362 18464 18426 18468
rect 18442 18524 18506 18528
rect 18442 18468 18446 18524
rect 18446 18468 18502 18524
rect 18502 18468 18506 18524
rect 18442 18464 18506 18468
rect 7852 17980 7916 17984
rect 7852 17924 7856 17980
rect 7856 17924 7912 17980
rect 7912 17924 7916 17980
rect 7852 17920 7916 17924
rect 7932 17980 7996 17984
rect 7932 17924 7936 17980
rect 7936 17924 7992 17980
rect 7992 17924 7996 17980
rect 7932 17920 7996 17924
rect 8012 17980 8076 17984
rect 8012 17924 8016 17980
rect 8016 17924 8072 17980
rect 8072 17924 8076 17980
rect 8012 17920 8076 17924
rect 8092 17980 8156 17984
rect 8092 17924 8096 17980
rect 8096 17924 8152 17980
rect 8152 17924 8156 17980
rect 8092 17920 8156 17924
rect 14752 17980 14816 17984
rect 14752 17924 14756 17980
rect 14756 17924 14812 17980
rect 14812 17924 14816 17980
rect 14752 17920 14816 17924
rect 14832 17980 14896 17984
rect 14832 17924 14836 17980
rect 14836 17924 14892 17980
rect 14892 17924 14896 17980
rect 14832 17920 14896 17924
rect 14912 17980 14976 17984
rect 14912 17924 14916 17980
rect 14916 17924 14972 17980
rect 14972 17924 14976 17980
rect 14912 17920 14976 17924
rect 14992 17980 15056 17984
rect 14992 17924 14996 17980
rect 14996 17924 15052 17980
rect 15052 17924 15056 17980
rect 14992 17920 15056 17924
rect 4402 17436 4466 17440
rect 4402 17380 4406 17436
rect 4406 17380 4462 17436
rect 4462 17380 4466 17436
rect 4402 17376 4466 17380
rect 4482 17436 4546 17440
rect 4482 17380 4486 17436
rect 4486 17380 4542 17436
rect 4542 17380 4546 17436
rect 4482 17376 4546 17380
rect 4562 17436 4626 17440
rect 4562 17380 4566 17436
rect 4566 17380 4622 17436
rect 4622 17380 4626 17436
rect 4562 17376 4626 17380
rect 4642 17436 4706 17440
rect 4642 17380 4646 17436
rect 4646 17380 4702 17436
rect 4702 17380 4706 17436
rect 4642 17376 4706 17380
rect 11302 17436 11366 17440
rect 11302 17380 11306 17436
rect 11306 17380 11362 17436
rect 11362 17380 11366 17436
rect 11302 17376 11366 17380
rect 11382 17436 11446 17440
rect 11382 17380 11386 17436
rect 11386 17380 11442 17436
rect 11442 17380 11446 17436
rect 11382 17376 11446 17380
rect 11462 17436 11526 17440
rect 11462 17380 11466 17436
rect 11466 17380 11522 17436
rect 11522 17380 11526 17436
rect 11462 17376 11526 17380
rect 11542 17436 11606 17440
rect 11542 17380 11546 17436
rect 11546 17380 11602 17436
rect 11602 17380 11606 17436
rect 11542 17376 11606 17380
rect 18202 17436 18266 17440
rect 18202 17380 18206 17436
rect 18206 17380 18262 17436
rect 18262 17380 18266 17436
rect 18202 17376 18266 17380
rect 18282 17436 18346 17440
rect 18282 17380 18286 17436
rect 18286 17380 18342 17436
rect 18342 17380 18346 17436
rect 18282 17376 18346 17380
rect 18362 17436 18426 17440
rect 18362 17380 18366 17436
rect 18366 17380 18422 17436
rect 18422 17380 18426 17436
rect 18362 17376 18426 17380
rect 18442 17436 18506 17440
rect 18442 17380 18446 17436
rect 18446 17380 18502 17436
rect 18502 17380 18506 17436
rect 18442 17376 18506 17380
rect 7852 16892 7916 16896
rect 7852 16836 7856 16892
rect 7856 16836 7912 16892
rect 7912 16836 7916 16892
rect 7852 16832 7916 16836
rect 7932 16892 7996 16896
rect 7932 16836 7936 16892
rect 7936 16836 7992 16892
rect 7992 16836 7996 16892
rect 7932 16832 7996 16836
rect 8012 16892 8076 16896
rect 8012 16836 8016 16892
rect 8016 16836 8072 16892
rect 8072 16836 8076 16892
rect 8012 16832 8076 16836
rect 8092 16892 8156 16896
rect 8092 16836 8096 16892
rect 8096 16836 8152 16892
rect 8152 16836 8156 16892
rect 8092 16832 8156 16836
rect 14752 16892 14816 16896
rect 14752 16836 14756 16892
rect 14756 16836 14812 16892
rect 14812 16836 14816 16892
rect 14752 16832 14816 16836
rect 14832 16892 14896 16896
rect 14832 16836 14836 16892
rect 14836 16836 14892 16892
rect 14892 16836 14896 16892
rect 14832 16832 14896 16836
rect 14912 16892 14976 16896
rect 14912 16836 14916 16892
rect 14916 16836 14972 16892
rect 14972 16836 14976 16892
rect 14912 16832 14976 16836
rect 14992 16892 15056 16896
rect 14992 16836 14996 16892
rect 14996 16836 15052 16892
rect 15052 16836 15056 16892
rect 14992 16832 15056 16836
rect 4402 16348 4466 16352
rect 4402 16292 4406 16348
rect 4406 16292 4462 16348
rect 4462 16292 4466 16348
rect 4402 16288 4466 16292
rect 4482 16348 4546 16352
rect 4482 16292 4486 16348
rect 4486 16292 4542 16348
rect 4542 16292 4546 16348
rect 4482 16288 4546 16292
rect 4562 16348 4626 16352
rect 4562 16292 4566 16348
rect 4566 16292 4622 16348
rect 4622 16292 4626 16348
rect 4562 16288 4626 16292
rect 4642 16348 4706 16352
rect 4642 16292 4646 16348
rect 4646 16292 4702 16348
rect 4702 16292 4706 16348
rect 4642 16288 4706 16292
rect 11302 16348 11366 16352
rect 11302 16292 11306 16348
rect 11306 16292 11362 16348
rect 11362 16292 11366 16348
rect 11302 16288 11366 16292
rect 11382 16348 11446 16352
rect 11382 16292 11386 16348
rect 11386 16292 11442 16348
rect 11442 16292 11446 16348
rect 11382 16288 11446 16292
rect 11462 16348 11526 16352
rect 11462 16292 11466 16348
rect 11466 16292 11522 16348
rect 11522 16292 11526 16348
rect 11462 16288 11526 16292
rect 11542 16348 11606 16352
rect 11542 16292 11546 16348
rect 11546 16292 11602 16348
rect 11602 16292 11606 16348
rect 11542 16288 11606 16292
rect 18202 16348 18266 16352
rect 18202 16292 18206 16348
rect 18206 16292 18262 16348
rect 18262 16292 18266 16348
rect 18202 16288 18266 16292
rect 18282 16348 18346 16352
rect 18282 16292 18286 16348
rect 18286 16292 18342 16348
rect 18342 16292 18346 16348
rect 18282 16288 18346 16292
rect 18362 16348 18426 16352
rect 18362 16292 18366 16348
rect 18366 16292 18422 16348
rect 18422 16292 18426 16348
rect 18362 16288 18426 16292
rect 18442 16348 18506 16352
rect 18442 16292 18446 16348
rect 18446 16292 18502 16348
rect 18502 16292 18506 16348
rect 18442 16288 18506 16292
rect 7852 15804 7916 15808
rect 7852 15748 7856 15804
rect 7856 15748 7912 15804
rect 7912 15748 7916 15804
rect 7852 15744 7916 15748
rect 7932 15804 7996 15808
rect 7932 15748 7936 15804
rect 7936 15748 7992 15804
rect 7992 15748 7996 15804
rect 7932 15744 7996 15748
rect 8012 15804 8076 15808
rect 8012 15748 8016 15804
rect 8016 15748 8072 15804
rect 8072 15748 8076 15804
rect 8012 15744 8076 15748
rect 8092 15804 8156 15808
rect 8092 15748 8096 15804
rect 8096 15748 8152 15804
rect 8152 15748 8156 15804
rect 8092 15744 8156 15748
rect 14752 15804 14816 15808
rect 14752 15748 14756 15804
rect 14756 15748 14812 15804
rect 14812 15748 14816 15804
rect 14752 15744 14816 15748
rect 14832 15804 14896 15808
rect 14832 15748 14836 15804
rect 14836 15748 14892 15804
rect 14892 15748 14896 15804
rect 14832 15744 14896 15748
rect 14912 15804 14976 15808
rect 14912 15748 14916 15804
rect 14916 15748 14972 15804
rect 14972 15748 14976 15804
rect 14912 15744 14976 15748
rect 14992 15804 15056 15808
rect 14992 15748 14996 15804
rect 14996 15748 15052 15804
rect 15052 15748 15056 15804
rect 14992 15744 15056 15748
rect 4402 15260 4466 15264
rect 4402 15204 4406 15260
rect 4406 15204 4462 15260
rect 4462 15204 4466 15260
rect 4402 15200 4466 15204
rect 4482 15260 4546 15264
rect 4482 15204 4486 15260
rect 4486 15204 4542 15260
rect 4542 15204 4546 15260
rect 4482 15200 4546 15204
rect 4562 15260 4626 15264
rect 4562 15204 4566 15260
rect 4566 15204 4622 15260
rect 4622 15204 4626 15260
rect 4562 15200 4626 15204
rect 4642 15260 4706 15264
rect 4642 15204 4646 15260
rect 4646 15204 4702 15260
rect 4702 15204 4706 15260
rect 4642 15200 4706 15204
rect 11302 15260 11366 15264
rect 11302 15204 11306 15260
rect 11306 15204 11362 15260
rect 11362 15204 11366 15260
rect 11302 15200 11366 15204
rect 11382 15260 11446 15264
rect 11382 15204 11386 15260
rect 11386 15204 11442 15260
rect 11442 15204 11446 15260
rect 11382 15200 11446 15204
rect 11462 15260 11526 15264
rect 11462 15204 11466 15260
rect 11466 15204 11522 15260
rect 11522 15204 11526 15260
rect 11462 15200 11526 15204
rect 11542 15260 11606 15264
rect 11542 15204 11546 15260
rect 11546 15204 11602 15260
rect 11602 15204 11606 15260
rect 11542 15200 11606 15204
rect 18202 15260 18266 15264
rect 18202 15204 18206 15260
rect 18206 15204 18262 15260
rect 18262 15204 18266 15260
rect 18202 15200 18266 15204
rect 18282 15260 18346 15264
rect 18282 15204 18286 15260
rect 18286 15204 18342 15260
rect 18342 15204 18346 15260
rect 18282 15200 18346 15204
rect 18362 15260 18426 15264
rect 18362 15204 18366 15260
rect 18366 15204 18422 15260
rect 18422 15204 18426 15260
rect 18362 15200 18426 15204
rect 18442 15260 18506 15264
rect 18442 15204 18446 15260
rect 18446 15204 18502 15260
rect 18502 15204 18506 15260
rect 18442 15200 18506 15204
rect 7852 14716 7916 14720
rect 7852 14660 7856 14716
rect 7856 14660 7912 14716
rect 7912 14660 7916 14716
rect 7852 14656 7916 14660
rect 7932 14716 7996 14720
rect 7932 14660 7936 14716
rect 7936 14660 7992 14716
rect 7992 14660 7996 14716
rect 7932 14656 7996 14660
rect 8012 14716 8076 14720
rect 8012 14660 8016 14716
rect 8016 14660 8072 14716
rect 8072 14660 8076 14716
rect 8012 14656 8076 14660
rect 8092 14716 8156 14720
rect 8092 14660 8096 14716
rect 8096 14660 8152 14716
rect 8152 14660 8156 14716
rect 8092 14656 8156 14660
rect 14752 14716 14816 14720
rect 14752 14660 14756 14716
rect 14756 14660 14812 14716
rect 14812 14660 14816 14716
rect 14752 14656 14816 14660
rect 14832 14716 14896 14720
rect 14832 14660 14836 14716
rect 14836 14660 14892 14716
rect 14892 14660 14896 14716
rect 14832 14656 14896 14660
rect 14912 14716 14976 14720
rect 14912 14660 14916 14716
rect 14916 14660 14972 14716
rect 14972 14660 14976 14716
rect 14912 14656 14976 14660
rect 14992 14716 15056 14720
rect 14992 14660 14996 14716
rect 14996 14660 15052 14716
rect 15052 14660 15056 14716
rect 14992 14656 15056 14660
rect 4402 14172 4466 14176
rect 4402 14116 4406 14172
rect 4406 14116 4462 14172
rect 4462 14116 4466 14172
rect 4402 14112 4466 14116
rect 4482 14172 4546 14176
rect 4482 14116 4486 14172
rect 4486 14116 4542 14172
rect 4542 14116 4546 14172
rect 4482 14112 4546 14116
rect 4562 14172 4626 14176
rect 4562 14116 4566 14172
rect 4566 14116 4622 14172
rect 4622 14116 4626 14172
rect 4562 14112 4626 14116
rect 4642 14172 4706 14176
rect 4642 14116 4646 14172
rect 4646 14116 4702 14172
rect 4702 14116 4706 14172
rect 4642 14112 4706 14116
rect 11302 14172 11366 14176
rect 11302 14116 11306 14172
rect 11306 14116 11362 14172
rect 11362 14116 11366 14172
rect 11302 14112 11366 14116
rect 11382 14172 11446 14176
rect 11382 14116 11386 14172
rect 11386 14116 11442 14172
rect 11442 14116 11446 14172
rect 11382 14112 11446 14116
rect 11462 14172 11526 14176
rect 11462 14116 11466 14172
rect 11466 14116 11522 14172
rect 11522 14116 11526 14172
rect 11462 14112 11526 14116
rect 11542 14172 11606 14176
rect 11542 14116 11546 14172
rect 11546 14116 11602 14172
rect 11602 14116 11606 14172
rect 11542 14112 11606 14116
rect 18202 14172 18266 14176
rect 18202 14116 18206 14172
rect 18206 14116 18262 14172
rect 18262 14116 18266 14172
rect 18202 14112 18266 14116
rect 18282 14172 18346 14176
rect 18282 14116 18286 14172
rect 18286 14116 18342 14172
rect 18342 14116 18346 14172
rect 18282 14112 18346 14116
rect 18362 14172 18426 14176
rect 18362 14116 18366 14172
rect 18366 14116 18422 14172
rect 18422 14116 18426 14172
rect 18362 14112 18426 14116
rect 18442 14172 18506 14176
rect 18442 14116 18446 14172
rect 18446 14116 18502 14172
rect 18502 14116 18506 14172
rect 18442 14112 18506 14116
rect 7852 13628 7916 13632
rect 7852 13572 7856 13628
rect 7856 13572 7912 13628
rect 7912 13572 7916 13628
rect 7852 13568 7916 13572
rect 7932 13628 7996 13632
rect 7932 13572 7936 13628
rect 7936 13572 7992 13628
rect 7992 13572 7996 13628
rect 7932 13568 7996 13572
rect 8012 13628 8076 13632
rect 8012 13572 8016 13628
rect 8016 13572 8072 13628
rect 8072 13572 8076 13628
rect 8012 13568 8076 13572
rect 8092 13628 8156 13632
rect 8092 13572 8096 13628
rect 8096 13572 8152 13628
rect 8152 13572 8156 13628
rect 8092 13568 8156 13572
rect 14752 13628 14816 13632
rect 14752 13572 14756 13628
rect 14756 13572 14812 13628
rect 14812 13572 14816 13628
rect 14752 13568 14816 13572
rect 14832 13628 14896 13632
rect 14832 13572 14836 13628
rect 14836 13572 14892 13628
rect 14892 13572 14896 13628
rect 14832 13568 14896 13572
rect 14912 13628 14976 13632
rect 14912 13572 14916 13628
rect 14916 13572 14972 13628
rect 14972 13572 14976 13628
rect 14912 13568 14976 13572
rect 14992 13628 15056 13632
rect 14992 13572 14996 13628
rect 14996 13572 15052 13628
rect 15052 13572 15056 13628
rect 14992 13568 15056 13572
rect 4402 13084 4466 13088
rect 4402 13028 4406 13084
rect 4406 13028 4462 13084
rect 4462 13028 4466 13084
rect 4402 13024 4466 13028
rect 4482 13084 4546 13088
rect 4482 13028 4486 13084
rect 4486 13028 4542 13084
rect 4542 13028 4546 13084
rect 4482 13024 4546 13028
rect 4562 13084 4626 13088
rect 4562 13028 4566 13084
rect 4566 13028 4622 13084
rect 4622 13028 4626 13084
rect 4562 13024 4626 13028
rect 4642 13084 4706 13088
rect 4642 13028 4646 13084
rect 4646 13028 4702 13084
rect 4702 13028 4706 13084
rect 4642 13024 4706 13028
rect 11302 13084 11366 13088
rect 11302 13028 11306 13084
rect 11306 13028 11362 13084
rect 11362 13028 11366 13084
rect 11302 13024 11366 13028
rect 11382 13084 11446 13088
rect 11382 13028 11386 13084
rect 11386 13028 11442 13084
rect 11442 13028 11446 13084
rect 11382 13024 11446 13028
rect 11462 13084 11526 13088
rect 11462 13028 11466 13084
rect 11466 13028 11522 13084
rect 11522 13028 11526 13084
rect 11462 13024 11526 13028
rect 11542 13084 11606 13088
rect 11542 13028 11546 13084
rect 11546 13028 11602 13084
rect 11602 13028 11606 13084
rect 11542 13024 11606 13028
rect 18202 13084 18266 13088
rect 18202 13028 18206 13084
rect 18206 13028 18262 13084
rect 18262 13028 18266 13084
rect 18202 13024 18266 13028
rect 18282 13084 18346 13088
rect 18282 13028 18286 13084
rect 18286 13028 18342 13084
rect 18342 13028 18346 13084
rect 18282 13024 18346 13028
rect 18362 13084 18426 13088
rect 18362 13028 18366 13084
rect 18366 13028 18422 13084
rect 18422 13028 18426 13084
rect 18362 13024 18426 13028
rect 18442 13084 18506 13088
rect 18442 13028 18446 13084
rect 18446 13028 18502 13084
rect 18502 13028 18506 13084
rect 18442 13024 18506 13028
rect 7852 12540 7916 12544
rect 7852 12484 7856 12540
rect 7856 12484 7912 12540
rect 7912 12484 7916 12540
rect 7852 12480 7916 12484
rect 7932 12540 7996 12544
rect 7932 12484 7936 12540
rect 7936 12484 7992 12540
rect 7992 12484 7996 12540
rect 7932 12480 7996 12484
rect 8012 12540 8076 12544
rect 8012 12484 8016 12540
rect 8016 12484 8072 12540
rect 8072 12484 8076 12540
rect 8012 12480 8076 12484
rect 8092 12540 8156 12544
rect 8092 12484 8096 12540
rect 8096 12484 8152 12540
rect 8152 12484 8156 12540
rect 8092 12480 8156 12484
rect 14752 12540 14816 12544
rect 14752 12484 14756 12540
rect 14756 12484 14812 12540
rect 14812 12484 14816 12540
rect 14752 12480 14816 12484
rect 14832 12540 14896 12544
rect 14832 12484 14836 12540
rect 14836 12484 14892 12540
rect 14892 12484 14896 12540
rect 14832 12480 14896 12484
rect 14912 12540 14976 12544
rect 14912 12484 14916 12540
rect 14916 12484 14972 12540
rect 14972 12484 14976 12540
rect 14912 12480 14976 12484
rect 14992 12540 15056 12544
rect 14992 12484 14996 12540
rect 14996 12484 15052 12540
rect 15052 12484 15056 12540
rect 14992 12480 15056 12484
rect 4402 11996 4466 12000
rect 4402 11940 4406 11996
rect 4406 11940 4462 11996
rect 4462 11940 4466 11996
rect 4402 11936 4466 11940
rect 4482 11996 4546 12000
rect 4482 11940 4486 11996
rect 4486 11940 4542 11996
rect 4542 11940 4546 11996
rect 4482 11936 4546 11940
rect 4562 11996 4626 12000
rect 4562 11940 4566 11996
rect 4566 11940 4622 11996
rect 4622 11940 4626 11996
rect 4562 11936 4626 11940
rect 4642 11996 4706 12000
rect 4642 11940 4646 11996
rect 4646 11940 4702 11996
rect 4702 11940 4706 11996
rect 4642 11936 4706 11940
rect 11302 11996 11366 12000
rect 11302 11940 11306 11996
rect 11306 11940 11362 11996
rect 11362 11940 11366 11996
rect 11302 11936 11366 11940
rect 11382 11996 11446 12000
rect 11382 11940 11386 11996
rect 11386 11940 11442 11996
rect 11442 11940 11446 11996
rect 11382 11936 11446 11940
rect 11462 11996 11526 12000
rect 11462 11940 11466 11996
rect 11466 11940 11522 11996
rect 11522 11940 11526 11996
rect 11462 11936 11526 11940
rect 11542 11996 11606 12000
rect 11542 11940 11546 11996
rect 11546 11940 11602 11996
rect 11602 11940 11606 11996
rect 11542 11936 11606 11940
rect 18202 11996 18266 12000
rect 18202 11940 18206 11996
rect 18206 11940 18262 11996
rect 18262 11940 18266 11996
rect 18202 11936 18266 11940
rect 18282 11996 18346 12000
rect 18282 11940 18286 11996
rect 18286 11940 18342 11996
rect 18342 11940 18346 11996
rect 18282 11936 18346 11940
rect 18362 11996 18426 12000
rect 18362 11940 18366 11996
rect 18366 11940 18422 11996
rect 18422 11940 18426 11996
rect 18362 11936 18426 11940
rect 18442 11996 18506 12000
rect 18442 11940 18446 11996
rect 18446 11940 18502 11996
rect 18502 11940 18506 11996
rect 18442 11936 18506 11940
rect 7852 11452 7916 11456
rect 7852 11396 7856 11452
rect 7856 11396 7912 11452
rect 7912 11396 7916 11452
rect 7852 11392 7916 11396
rect 7932 11452 7996 11456
rect 7932 11396 7936 11452
rect 7936 11396 7992 11452
rect 7992 11396 7996 11452
rect 7932 11392 7996 11396
rect 8012 11452 8076 11456
rect 8012 11396 8016 11452
rect 8016 11396 8072 11452
rect 8072 11396 8076 11452
rect 8012 11392 8076 11396
rect 8092 11452 8156 11456
rect 8092 11396 8096 11452
rect 8096 11396 8152 11452
rect 8152 11396 8156 11452
rect 8092 11392 8156 11396
rect 14752 11452 14816 11456
rect 14752 11396 14756 11452
rect 14756 11396 14812 11452
rect 14812 11396 14816 11452
rect 14752 11392 14816 11396
rect 14832 11452 14896 11456
rect 14832 11396 14836 11452
rect 14836 11396 14892 11452
rect 14892 11396 14896 11452
rect 14832 11392 14896 11396
rect 14912 11452 14976 11456
rect 14912 11396 14916 11452
rect 14916 11396 14972 11452
rect 14972 11396 14976 11452
rect 14912 11392 14976 11396
rect 14992 11452 15056 11456
rect 14992 11396 14996 11452
rect 14996 11396 15052 11452
rect 15052 11396 15056 11452
rect 14992 11392 15056 11396
rect 4402 10908 4466 10912
rect 4402 10852 4406 10908
rect 4406 10852 4462 10908
rect 4462 10852 4466 10908
rect 4402 10848 4466 10852
rect 4482 10908 4546 10912
rect 4482 10852 4486 10908
rect 4486 10852 4542 10908
rect 4542 10852 4546 10908
rect 4482 10848 4546 10852
rect 4562 10908 4626 10912
rect 4562 10852 4566 10908
rect 4566 10852 4622 10908
rect 4622 10852 4626 10908
rect 4562 10848 4626 10852
rect 4642 10908 4706 10912
rect 4642 10852 4646 10908
rect 4646 10852 4702 10908
rect 4702 10852 4706 10908
rect 4642 10848 4706 10852
rect 11302 10908 11366 10912
rect 11302 10852 11306 10908
rect 11306 10852 11362 10908
rect 11362 10852 11366 10908
rect 11302 10848 11366 10852
rect 11382 10908 11446 10912
rect 11382 10852 11386 10908
rect 11386 10852 11442 10908
rect 11442 10852 11446 10908
rect 11382 10848 11446 10852
rect 11462 10908 11526 10912
rect 11462 10852 11466 10908
rect 11466 10852 11522 10908
rect 11522 10852 11526 10908
rect 11462 10848 11526 10852
rect 11542 10908 11606 10912
rect 11542 10852 11546 10908
rect 11546 10852 11602 10908
rect 11602 10852 11606 10908
rect 11542 10848 11606 10852
rect 18202 10908 18266 10912
rect 18202 10852 18206 10908
rect 18206 10852 18262 10908
rect 18262 10852 18266 10908
rect 18202 10848 18266 10852
rect 18282 10908 18346 10912
rect 18282 10852 18286 10908
rect 18286 10852 18342 10908
rect 18342 10852 18346 10908
rect 18282 10848 18346 10852
rect 18362 10908 18426 10912
rect 18362 10852 18366 10908
rect 18366 10852 18422 10908
rect 18422 10852 18426 10908
rect 18362 10848 18426 10852
rect 18442 10908 18506 10912
rect 18442 10852 18446 10908
rect 18446 10852 18502 10908
rect 18502 10852 18506 10908
rect 18442 10848 18506 10852
rect 7852 10364 7916 10368
rect 7852 10308 7856 10364
rect 7856 10308 7912 10364
rect 7912 10308 7916 10364
rect 7852 10304 7916 10308
rect 7932 10364 7996 10368
rect 7932 10308 7936 10364
rect 7936 10308 7992 10364
rect 7992 10308 7996 10364
rect 7932 10304 7996 10308
rect 8012 10364 8076 10368
rect 8012 10308 8016 10364
rect 8016 10308 8072 10364
rect 8072 10308 8076 10364
rect 8012 10304 8076 10308
rect 8092 10364 8156 10368
rect 8092 10308 8096 10364
rect 8096 10308 8152 10364
rect 8152 10308 8156 10364
rect 8092 10304 8156 10308
rect 14752 10364 14816 10368
rect 14752 10308 14756 10364
rect 14756 10308 14812 10364
rect 14812 10308 14816 10364
rect 14752 10304 14816 10308
rect 14832 10364 14896 10368
rect 14832 10308 14836 10364
rect 14836 10308 14892 10364
rect 14892 10308 14896 10364
rect 14832 10304 14896 10308
rect 14912 10364 14976 10368
rect 14912 10308 14916 10364
rect 14916 10308 14972 10364
rect 14972 10308 14976 10364
rect 14912 10304 14976 10308
rect 14992 10364 15056 10368
rect 14992 10308 14996 10364
rect 14996 10308 15052 10364
rect 15052 10308 15056 10364
rect 14992 10304 15056 10308
rect 4402 9820 4466 9824
rect 4402 9764 4406 9820
rect 4406 9764 4462 9820
rect 4462 9764 4466 9820
rect 4402 9760 4466 9764
rect 4482 9820 4546 9824
rect 4482 9764 4486 9820
rect 4486 9764 4542 9820
rect 4542 9764 4546 9820
rect 4482 9760 4546 9764
rect 4562 9820 4626 9824
rect 4562 9764 4566 9820
rect 4566 9764 4622 9820
rect 4622 9764 4626 9820
rect 4562 9760 4626 9764
rect 4642 9820 4706 9824
rect 4642 9764 4646 9820
rect 4646 9764 4702 9820
rect 4702 9764 4706 9820
rect 4642 9760 4706 9764
rect 11302 9820 11366 9824
rect 11302 9764 11306 9820
rect 11306 9764 11362 9820
rect 11362 9764 11366 9820
rect 11302 9760 11366 9764
rect 11382 9820 11446 9824
rect 11382 9764 11386 9820
rect 11386 9764 11442 9820
rect 11442 9764 11446 9820
rect 11382 9760 11446 9764
rect 11462 9820 11526 9824
rect 11462 9764 11466 9820
rect 11466 9764 11522 9820
rect 11522 9764 11526 9820
rect 11462 9760 11526 9764
rect 11542 9820 11606 9824
rect 11542 9764 11546 9820
rect 11546 9764 11602 9820
rect 11602 9764 11606 9820
rect 11542 9760 11606 9764
rect 18202 9820 18266 9824
rect 18202 9764 18206 9820
rect 18206 9764 18262 9820
rect 18262 9764 18266 9820
rect 18202 9760 18266 9764
rect 18282 9820 18346 9824
rect 18282 9764 18286 9820
rect 18286 9764 18342 9820
rect 18342 9764 18346 9820
rect 18282 9760 18346 9764
rect 18362 9820 18426 9824
rect 18362 9764 18366 9820
rect 18366 9764 18422 9820
rect 18422 9764 18426 9820
rect 18362 9760 18426 9764
rect 18442 9820 18506 9824
rect 18442 9764 18446 9820
rect 18446 9764 18502 9820
rect 18502 9764 18506 9820
rect 18442 9760 18506 9764
rect 7852 9276 7916 9280
rect 7852 9220 7856 9276
rect 7856 9220 7912 9276
rect 7912 9220 7916 9276
rect 7852 9216 7916 9220
rect 7932 9276 7996 9280
rect 7932 9220 7936 9276
rect 7936 9220 7992 9276
rect 7992 9220 7996 9276
rect 7932 9216 7996 9220
rect 8012 9276 8076 9280
rect 8012 9220 8016 9276
rect 8016 9220 8072 9276
rect 8072 9220 8076 9276
rect 8012 9216 8076 9220
rect 8092 9276 8156 9280
rect 8092 9220 8096 9276
rect 8096 9220 8152 9276
rect 8152 9220 8156 9276
rect 8092 9216 8156 9220
rect 14752 9276 14816 9280
rect 14752 9220 14756 9276
rect 14756 9220 14812 9276
rect 14812 9220 14816 9276
rect 14752 9216 14816 9220
rect 14832 9276 14896 9280
rect 14832 9220 14836 9276
rect 14836 9220 14892 9276
rect 14892 9220 14896 9276
rect 14832 9216 14896 9220
rect 14912 9276 14976 9280
rect 14912 9220 14916 9276
rect 14916 9220 14972 9276
rect 14972 9220 14976 9276
rect 14912 9216 14976 9220
rect 14992 9276 15056 9280
rect 14992 9220 14996 9276
rect 14996 9220 15052 9276
rect 15052 9220 15056 9276
rect 14992 9216 15056 9220
rect 4402 8732 4466 8736
rect 4402 8676 4406 8732
rect 4406 8676 4462 8732
rect 4462 8676 4466 8732
rect 4402 8672 4466 8676
rect 4482 8732 4546 8736
rect 4482 8676 4486 8732
rect 4486 8676 4542 8732
rect 4542 8676 4546 8732
rect 4482 8672 4546 8676
rect 4562 8732 4626 8736
rect 4562 8676 4566 8732
rect 4566 8676 4622 8732
rect 4622 8676 4626 8732
rect 4562 8672 4626 8676
rect 4642 8732 4706 8736
rect 4642 8676 4646 8732
rect 4646 8676 4702 8732
rect 4702 8676 4706 8732
rect 4642 8672 4706 8676
rect 11302 8732 11366 8736
rect 11302 8676 11306 8732
rect 11306 8676 11362 8732
rect 11362 8676 11366 8732
rect 11302 8672 11366 8676
rect 11382 8732 11446 8736
rect 11382 8676 11386 8732
rect 11386 8676 11442 8732
rect 11442 8676 11446 8732
rect 11382 8672 11446 8676
rect 11462 8732 11526 8736
rect 11462 8676 11466 8732
rect 11466 8676 11522 8732
rect 11522 8676 11526 8732
rect 11462 8672 11526 8676
rect 11542 8732 11606 8736
rect 11542 8676 11546 8732
rect 11546 8676 11602 8732
rect 11602 8676 11606 8732
rect 11542 8672 11606 8676
rect 18202 8732 18266 8736
rect 18202 8676 18206 8732
rect 18206 8676 18262 8732
rect 18262 8676 18266 8732
rect 18202 8672 18266 8676
rect 18282 8732 18346 8736
rect 18282 8676 18286 8732
rect 18286 8676 18342 8732
rect 18342 8676 18346 8732
rect 18282 8672 18346 8676
rect 18362 8732 18426 8736
rect 18362 8676 18366 8732
rect 18366 8676 18422 8732
rect 18422 8676 18426 8732
rect 18362 8672 18426 8676
rect 18442 8732 18506 8736
rect 18442 8676 18446 8732
rect 18446 8676 18502 8732
rect 18502 8676 18506 8732
rect 18442 8672 18506 8676
rect 7852 8188 7916 8192
rect 7852 8132 7856 8188
rect 7856 8132 7912 8188
rect 7912 8132 7916 8188
rect 7852 8128 7916 8132
rect 7932 8188 7996 8192
rect 7932 8132 7936 8188
rect 7936 8132 7992 8188
rect 7992 8132 7996 8188
rect 7932 8128 7996 8132
rect 8012 8188 8076 8192
rect 8012 8132 8016 8188
rect 8016 8132 8072 8188
rect 8072 8132 8076 8188
rect 8012 8128 8076 8132
rect 8092 8188 8156 8192
rect 8092 8132 8096 8188
rect 8096 8132 8152 8188
rect 8152 8132 8156 8188
rect 8092 8128 8156 8132
rect 14752 8188 14816 8192
rect 14752 8132 14756 8188
rect 14756 8132 14812 8188
rect 14812 8132 14816 8188
rect 14752 8128 14816 8132
rect 14832 8188 14896 8192
rect 14832 8132 14836 8188
rect 14836 8132 14892 8188
rect 14892 8132 14896 8188
rect 14832 8128 14896 8132
rect 14912 8188 14976 8192
rect 14912 8132 14916 8188
rect 14916 8132 14972 8188
rect 14972 8132 14976 8188
rect 14912 8128 14976 8132
rect 14992 8188 15056 8192
rect 14992 8132 14996 8188
rect 14996 8132 15052 8188
rect 15052 8132 15056 8188
rect 14992 8128 15056 8132
rect 4402 7644 4466 7648
rect 4402 7588 4406 7644
rect 4406 7588 4462 7644
rect 4462 7588 4466 7644
rect 4402 7584 4466 7588
rect 4482 7644 4546 7648
rect 4482 7588 4486 7644
rect 4486 7588 4542 7644
rect 4542 7588 4546 7644
rect 4482 7584 4546 7588
rect 4562 7644 4626 7648
rect 4562 7588 4566 7644
rect 4566 7588 4622 7644
rect 4622 7588 4626 7644
rect 4562 7584 4626 7588
rect 4642 7644 4706 7648
rect 4642 7588 4646 7644
rect 4646 7588 4702 7644
rect 4702 7588 4706 7644
rect 4642 7584 4706 7588
rect 11302 7644 11366 7648
rect 11302 7588 11306 7644
rect 11306 7588 11362 7644
rect 11362 7588 11366 7644
rect 11302 7584 11366 7588
rect 11382 7644 11446 7648
rect 11382 7588 11386 7644
rect 11386 7588 11442 7644
rect 11442 7588 11446 7644
rect 11382 7584 11446 7588
rect 11462 7644 11526 7648
rect 11462 7588 11466 7644
rect 11466 7588 11522 7644
rect 11522 7588 11526 7644
rect 11462 7584 11526 7588
rect 11542 7644 11606 7648
rect 11542 7588 11546 7644
rect 11546 7588 11602 7644
rect 11602 7588 11606 7644
rect 11542 7584 11606 7588
rect 18202 7644 18266 7648
rect 18202 7588 18206 7644
rect 18206 7588 18262 7644
rect 18262 7588 18266 7644
rect 18202 7584 18266 7588
rect 18282 7644 18346 7648
rect 18282 7588 18286 7644
rect 18286 7588 18342 7644
rect 18342 7588 18346 7644
rect 18282 7584 18346 7588
rect 18362 7644 18426 7648
rect 18362 7588 18366 7644
rect 18366 7588 18422 7644
rect 18422 7588 18426 7644
rect 18362 7584 18426 7588
rect 18442 7644 18506 7648
rect 18442 7588 18446 7644
rect 18446 7588 18502 7644
rect 18502 7588 18506 7644
rect 18442 7584 18506 7588
rect 7852 7100 7916 7104
rect 7852 7044 7856 7100
rect 7856 7044 7912 7100
rect 7912 7044 7916 7100
rect 7852 7040 7916 7044
rect 7932 7100 7996 7104
rect 7932 7044 7936 7100
rect 7936 7044 7992 7100
rect 7992 7044 7996 7100
rect 7932 7040 7996 7044
rect 8012 7100 8076 7104
rect 8012 7044 8016 7100
rect 8016 7044 8072 7100
rect 8072 7044 8076 7100
rect 8012 7040 8076 7044
rect 8092 7100 8156 7104
rect 8092 7044 8096 7100
rect 8096 7044 8152 7100
rect 8152 7044 8156 7100
rect 8092 7040 8156 7044
rect 14752 7100 14816 7104
rect 14752 7044 14756 7100
rect 14756 7044 14812 7100
rect 14812 7044 14816 7100
rect 14752 7040 14816 7044
rect 14832 7100 14896 7104
rect 14832 7044 14836 7100
rect 14836 7044 14892 7100
rect 14892 7044 14896 7100
rect 14832 7040 14896 7044
rect 14912 7100 14976 7104
rect 14912 7044 14916 7100
rect 14916 7044 14972 7100
rect 14972 7044 14976 7100
rect 14912 7040 14976 7044
rect 14992 7100 15056 7104
rect 14992 7044 14996 7100
rect 14996 7044 15052 7100
rect 15052 7044 15056 7100
rect 14992 7040 15056 7044
rect 4402 6556 4466 6560
rect 4402 6500 4406 6556
rect 4406 6500 4462 6556
rect 4462 6500 4466 6556
rect 4402 6496 4466 6500
rect 4482 6556 4546 6560
rect 4482 6500 4486 6556
rect 4486 6500 4542 6556
rect 4542 6500 4546 6556
rect 4482 6496 4546 6500
rect 4562 6556 4626 6560
rect 4562 6500 4566 6556
rect 4566 6500 4622 6556
rect 4622 6500 4626 6556
rect 4562 6496 4626 6500
rect 4642 6556 4706 6560
rect 4642 6500 4646 6556
rect 4646 6500 4702 6556
rect 4702 6500 4706 6556
rect 4642 6496 4706 6500
rect 11302 6556 11366 6560
rect 11302 6500 11306 6556
rect 11306 6500 11362 6556
rect 11362 6500 11366 6556
rect 11302 6496 11366 6500
rect 11382 6556 11446 6560
rect 11382 6500 11386 6556
rect 11386 6500 11442 6556
rect 11442 6500 11446 6556
rect 11382 6496 11446 6500
rect 11462 6556 11526 6560
rect 11462 6500 11466 6556
rect 11466 6500 11522 6556
rect 11522 6500 11526 6556
rect 11462 6496 11526 6500
rect 11542 6556 11606 6560
rect 11542 6500 11546 6556
rect 11546 6500 11602 6556
rect 11602 6500 11606 6556
rect 11542 6496 11606 6500
rect 18202 6556 18266 6560
rect 18202 6500 18206 6556
rect 18206 6500 18262 6556
rect 18262 6500 18266 6556
rect 18202 6496 18266 6500
rect 18282 6556 18346 6560
rect 18282 6500 18286 6556
rect 18286 6500 18342 6556
rect 18342 6500 18346 6556
rect 18282 6496 18346 6500
rect 18362 6556 18426 6560
rect 18362 6500 18366 6556
rect 18366 6500 18422 6556
rect 18422 6500 18426 6556
rect 18362 6496 18426 6500
rect 18442 6556 18506 6560
rect 18442 6500 18446 6556
rect 18446 6500 18502 6556
rect 18502 6500 18506 6556
rect 18442 6496 18506 6500
rect 7852 6012 7916 6016
rect 7852 5956 7856 6012
rect 7856 5956 7912 6012
rect 7912 5956 7916 6012
rect 7852 5952 7916 5956
rect 7932 6012 7996 6016
rect 7932 5956 7936 6012
rect 7936 5956 7992 6012
rect 7992 5956 7996 6012
rect 7932 5952 7996 5956
rect 8012 6012 8076 6016
rect 8012 5956 8016 6012
rect 8016 5956 8072 6012
rect 8072 5956 8076 6012
rect 8012 5952 8076 5956
rect 8092 6012 8156 6016
rect 8092 5956 8096 6012
rect 8096 5956 8152 6012
rect 8152 5956 8156 6012
rect 8092 5952 8156 5956
rect 14752 6012 14816 6016
rect 14752 5956 14756 6012
rect 14756 5956 14812 6012
rect 14812 5956 14816 6012
rect 14752 5952 14816 5956
rect 14832 6012 14896 6016
rect 14832 5956 14836 6012
rect 14836 5956 14892 6012
rect 14892 5956 14896 6012
rect 14832 5952 14896 5956
rect 14912 6012 14976 6016
rect 14912 5956 14916 6012
rect 14916 5956 14972 6012
rect 14972 5956 14976 6012
rect 14912 5952 14976 5956
rect 14992 6012 15056 6016
rect 14992 5956 14996 6012
rect 14996 5956 15052 6012
rect 15052 5956 15056 6012
rect 14992 5952 15056 5956
rect 4402 5468 4466 5472
rect 4402 5412 4406 5468
rect 4406 5412 4462 5468
rect 4462 5412 4466 5468
rect 4402 5408 4466 5412
rect 4482 5468 4546 5472
rect 4482 5412 4486 5468
rect 4486 5412 4542 5468
rect 4542 5412 4546 5468
rect 4482 5408 4546 5412
rect 4562 5468 4626 5472
rect 4562 5412 4566 5468
rect 4566 5412 4622 5468
rect 4622 5412 4626 5468
rect 4562 5408 4626 5412
rect 4642 5468 4706 5472
rect 4642 5412 4646 5468
rect 4646 5412 4702 5468
rect 4702 5412 4706 5468
rect 4642 5408 4706 5412
rect 11302 5468 11366 5472
rect 11302 5412 11306 5468
rect 11306 5412 11362 5468
rect 11362 5412 11366 5468
rect 11302 5408 11366 5412
rect 11382 5468 11446 5472
rect 11382 5412 11386 5468
rect 11386 5412 11442 5468
rect 11442 5412 11446 5468
rect 11382 5408 11446 5412
rect 11462 5468 11526 5472
rect 11462 5412 11466 5468
rect 11466 5412 11522 5468
rect 11522 5412 11526 5468
rect 11462 5408 11526 5412
rect 11542 5468 11606 5472
rect 11542 5412 11546 5468
rect 11546 5412 11602 5468
rect 11602 5412 11606 5468
rect 11542 5408 11606 5412
rect 18202 5468 18266 5472
rect 18202 5412 18206 5468
rect 18206 5412 18262 5468
rect 18262 5412 18266 5468
rect 18202 5408 18266 5412
rect 18282 5468 18346 5472
rect 18282 5412 18286 5468
rect 18286 5412 18342 5468
rect 18342 5412 18346 5468
rect 18282 5408 18346 5412
rect 18362 5468 18426 5472
rect 18362 5412 18366 5468
rect 18366 5412 18422 5468
rect 18422 5412 18426 5468
rect 18362 5408 18426 5412
rect 18442 5468 18506 5472
rect 18442 5412 18446 5468
rect 18446 5412 18502 5468
rect 18502 5412 18506 5468
rect 18442 5408 18506 5412
rect 7852 4924 7916 4928
rect 7852 4868 7856 4924
rect 7856 4868 7912 4924
rect 7912 4868 7916 4924
rect 7852 4864 7916 4868
rect 7932 4924 7996 4928
rect 7932 4868 7936 4924
rect 7936 4868 7992 4924
rect 7992 4868 7996 4924
rect 7932 4864 7996 4868
rect 8012 4924 8076 4928
rect 8012 4868 8016 4924
rect 8016 4868 8072 4924
rect 8072 4868 8076 4924
rect 8012 4864 8076 4868
rect 8092 4924 8156 4928
rect 8092 4868 8096 4924
rect 8096 4868 8152 4924
rect 8152 4868 8156 4924
rect 8092 4864 8156 4868
rect 14752 4924 14816 4928
rect 14752 4868 14756 4924
rect 14756 4868 14812 4924
rect 14812 4868 14816 4924
rect 14752 4864 14816 4868
rect 14832 4924 14896 4928
rect 14832 4868 14836 4924
rect 14836 4868 14892 4924
rect 14892 4868 14896 4924
rect 14832 4864 14896 4868
rect 14912 4924 14976 4928
rect 14912 4868 14916 4924
rect 14916 4868 14972 4924
rect 14972 4868 14976 4924
rect 14912 4864 14976 4868
rect 14992 4924 15056 4928
rect 14992 4868 14996 4924
rect 14996 4868 15052 4924
rect 15052 4868 15056 4924
rect 14992 4864 15056 4868
rect 4402 4380 4466 4384
rect 4402 4324 4406 4380
rect 4406 4324 4462 4380
rect 4462 4324 4466 4380
rect 4402 4320 4466 4324
rect 4482 4380 4546 4384
rect 4482 4324 4486 4380
rect 4486 4324 4542 4380
rect 4542 4324 4546 4380
rect 4482 4320 4546 4324
rect 4562 4380 4626 4384
rect 4562 4324 4566 4380
rect 4566 4324 4622 4380
rect 4622 4324 4626 4380
rect 4562 4320 4626 4324
rect 4642 4380 4706 4384
rect 4642 4324 4646 4380
rect 4646 4324 4702 4380
rect 4702 4324 4706 4380
rect 4642 4320 4706 4324
rect 11302 4380 11366 4384
rect 11302 4324 11306 4380
rect 11306 4324 11362 4380
rect 11362 4324 11366 4380
rect 11302 4320 11366 4324
rect 11382 4380 11446 4384
rect 11382 4324 11386 4380
rect 11386 4324 11442 4380
rect 11442 4324 11446 4380
rect 11382 4320 11446 4324
rect 11462 4380 11526 4384
rect 11462 4324 11466 4380
rect 11466 4324 11522 4380
rect 11522 4324 11526 4380
rect 11462 4320 11526 4324
rect 11542 4380 11606 4384
rect 11542 4324 11546 4380
rect 11546 4324 11602 4380
rect 11602 4324 11606 4380
rect 11542 4320 11606 4324
rect 18202 4380 18266 4384
rect 18202 4324 18206 4380
rect 18206 4324 18262 4380
rect 18262 4324 18266 4380
rect 18202 4320 18266 4324
rect 18282 4380 18346 4384
rect 18282 4324 18286 4380
rect 18286 4324 18342 4380
rect 18342 4324 18346 4380
rect 18282 4320 18346 4324
rect 18362 4380 18426 4384
rect 18362 4324 18366 4380
rect 18366 4324 18422 4380
rect 18422 4324 18426 4380
rect 18362 4320 18426 4324
rect 18442 4380 18506 4384
rect 18442 4324 18446 4380
rect 18446 4324 18502 4380
rect 18502 4324 18506 4380
rect 18442 4320 18506 4324
rect 7852 3836 7916 3840
rect 7852 3780 7856 3836
rect 7856 3780 7912 3836
rect 7912 3780 7916 3836
rect 7852 3776 7916 3780
rect 7932 3836 7996 3840
rect 7932 3780 7936 3836
rect 7936 3780 7992 3836
rect 7992 3780 7996 3836
rect 7932 3776 7996 3780
rect 8012 3836 8076 3840
rect 8012 3780 8016 3836
rect 8016 3780 8072 3836
rect 8072 3780 8076 3836
rect 8012 3776 8076 3780
rect 8092 3836 8156 3840
rect 8092 3780 8096 3836
rect 8096 3780 8152 3836
rect 8152 3780 8156 3836
rect 8092 3776 8156 3780
rect 14752 3836 14816 3840
rect 14752 3780 14756 3836
rect 14756 3780 14812 3836
rect 14812 3780 14816 3836
rect 14752 3776 14816 3780
rect 14832 3836 14896 3840
rect 14832 3780 14836 3836
rect 14836 3780 14892 3836
rect 14892 3780 14896 3836
rect 14832 3776 14896 3780
rect 14912 3836 14976 3840
rect 14912 3780 14916 3836
rect 14916 3780 14972 3836
rect 14972 3780 14976 3836
rect 14912 3776 14976 3780
rect 14992 3836 15056 3840
rect 14992 3780 14996 3836
rect 14996 3780 15052 3836
rect 15052 3780 15056 3836
rect 14992 3776 15056 3780
rect 4402 3292 4466 3296
rect 4402 3236 4406 3292
rect 4406 3236 4462 3292
rect 4462 3236 4466 3292
rect 4402 3232 4466 3236
rect 4482 3292 4546 3296
rect 4482 3236 4486 3292
rect 4486 3236 4542 3292
rect 4542 3236 4546 3292
rect 4482 3232 4546 3236
rect 4562 3292 4626 3296
rect 4562 3236 4566 3292
rect 4566 3236 4622 3292
rect 4622 3236 4626 3292
rect 4562 3232 4626 3236
rect 4642 3292 4706 3296
rect 4642 3236 4646 3292
rect 4646 3236 4702 3292
rect 4702 3236 4706 3292
rect 4642 3232 4706 3236
rect 11302 3292 11366 3296
rect 11302 3236 11306 3292
rect 11306 3236 11362 3292
rect 11362 3236 11366 3292
rect 11302 3232 11366 3236
rect 11382 3292 11446 3296
rect 11382 3236 11386 3292
rect 11386 3236 11442 3292
rect 11442 3236 11446 3292
rect 11382 3232 11446 3236
rect 11462 3292 11526 3296
rect 11462 3236 11466 3292
rect 11466 3236 11522 3292
rect 11522 3236 11526 3292
rect 11462 3232 11526 3236
rect 11542 3292 11606 3296
rect 11542 3236 11546 3292
rect 11546 3236 11602 3292
rect 11602 3236 11606 3292
rect 11542 3232 11606 3236
rect 18202 3292 18266 3296
rect 18202 3236 18206 3292
rect 18206 3236 18262 3292
rect 18262 3236 18266 3292
rect 18202 3232 18266 3236
rect 18282 3292 18346 3296
rect 18282 3236 18286 3292
rect 18286 3236 18342 3292
rect 18342 3236 18346 3292
rect 18282 3232 18346 3236
rect 18362 3292 18426 3296
rect 18362 3236 18366 3292
rect 18366 3236 18422 3292
rect 18422 3236 18426 3292
rect 18362 3232 18426 3236
rect 18442 3292 18506 3296
rect 18442 3236 18446 3292
rect 18446 3236 18502 3292
rect 18502 3236 18506 3292
rect 18442 3232 18506 3236
rect 7852 2748 7916 2752
rect 7852 2692 7856 2748
rect 7856 2692 7912 2748
rect 7912 2692 7916 2748
rect 7852 2688 7916 2692
rect 7932 2748 7996 2752
rect 7932 2692 7936 2748
rect 7936 2692 7992 2748
rect 7992 2692 7996 2748
rect 7932 2688 7996 2692
rect 8012 2748 8076 2752
rect 8012 2692 8016 2748
rect 8016 2692 8072 2748
rect 8072 2692 8076 2748
rect 8012 2688 8076 2692
rect 8092 2748 8156 2752
rect 8092 2692 8096 2748
rect 8096 2692 8152 2748
rect 8152 2692 8156 2748
rect 8092 2688 8156 2692
rect 14752 2748 14816 2752
rect 14752 2692 14756 2748
rect 14756 2692 14812 2748
rect 14812 2692 14816 2748
rect 14752 2688 14816 2692
rect 14832 2748 14896 2752
rect 14832 2692 14836 2748
rect 14836 2692 14892 2748
rect 14892 2692 14896 2748
rect 14832 2688 14896 2692
rect 14912 2748 14976 2752
rect 14912 2692 14916 2748
rect 14916 2692 14972 2748
rect 14972 2692 14976 2748
rect 14912 2688 14976 2692
rect 14992 2748 15056 2752
rect 14992 2692 14996 2748
rect 14996 2692 15052 2748
rect 15052 2692 15056 2748
rect 14992 2688 15056 2692
rect 4402 2204 4466 2208
rect 4402 2148 4406 2204
rect 4406 2148 4462 2204
rect 4462 2148 4466 2204
rect 4402 2144 4466 2148
rect 4482 2204 4546 2208
rect 4482 2148 4486 2204
rect 4486 2148 4542 2204
rect 4542 2148 4546 2204
rect 4482 2144 4546 2148
rect 4562 2204 4626 2208
rect 4562 2148 4566 2204
rect 4566 2148 4622 2204
rect 4622 2148 4626 2204
rect 4562 2144 4626 2148
rect 4642 2204 4706 2208
rect 4642 2148 4646 2204
rect 4646 2148 4702 2204
rect 4702 2148 4706 2204
rect 4642 2144 4706 2148
rect 11302 2204 11366 2208
rect 11302 2148 11306 2204
rect 11306 2148 11362 2204
rect 11362 2148 11366 2204
rect 11302 2144 11366 2148
rect 11382 2204 11446 2208
rect 11382 2148 11386 2204
rect 11386 2148 11442 2204
rect 11442 2148 11446 2204
rect 11382 2144 11446 2148
rect 11462 2204 11526 2208
rect 11462 2148 11466 2204
rect 11466 2148 11522 2204
rect 11522 2148 11526 2204
rect 11462 2144 11526 2148
rect 11542 2204 11606 2208
rect 11542 2148 11546 2204
rect 11546 2148 11602 2204
rect 11602 2148 11606 2204
rect 11542 2144 11606 2148
rect 18202 2204 18266 2208
rect 18202 2148 18206 2204
rect 18206 2148 18262 2204
rect 18262 2148 18266 2204
rect 18202 2144 18266 2148
rect 18282 2204 18346 2208
rect 18282 2148 18286 2204
rect 18286 2148 18342 2204
rect 18342 2148 18346 2204
rect 18282 2144 18346 2148
rect 18362 2204 18426 2208
rect 18362 2148 18366 2204
rect 18366 2148 18422 2204
rect 18422 2148 18426 2204
rect 18362 2144 18426 2148
rect 18442 2204 18506 2208
rect 18442 2148 18446 2204
rect 18446 2148 18502 2204
rect 18502 2148 18506 2204
rect 18442 2144 18506 2148
<< metal4 >>
rect 4394 22880 4714 22896
rect 4394 22816 4402 22880
rect 4466 22816 4482 22880
rect 4546 22816 4562 22880
rect 4626 22816 4642 22880
rect 4706 22816 4714 22880
rect 4394 21792 4714 22816
rect 4394 21728 4402 21792
rect 4466 21728 4482 21792
rect 4546 21728 4562 21792
rect 4626 21728 4642 21792
rect 4706 21728 4714 21792
rect 4394 20704 4714 21728
rect 4394 20640 4402 20704
rect 4466 20640 4482 20704
rect 4546 20640 4562 20704
rect 4626 20640 4642 20704
rect 4706 20640 4714 20704
rect 4394 19616 4714 20640
rect 4394 19552 4402 19616
rect 4466 19552 4482 19616
rect 4546 19552 4562 19616
rect 4626 19552 4642 19616
rect 4706 19552 4714 19616
rect 4394 19472 4714 19552
rect 4394 19236 4436 19472
rect 4672 19236 4714 19472
rect 4394 18528 4714 19236
rect 4394 18464 4402 18528
rect 4466 18464 4482 18528
rect 4546 18464 4562 18528
rect 4626 18464 4642 18528
rect 4706 18464 4714 18528
rect 4394 17440 4714 18464
rect 4394 17376 4402 17440
rect 4466 17376 4482 17440
rect 4546 17376 4562 17440
rect 4626 17376 4642 17440
rect 4706 17376 4714 17440
rect 4394 16352 4714 17376
rect 4394 16288 4402 16352
rect 4466 16288 4482 16352
rect 4546 16288 4562 16352
rect 4626 16288 4642 16352
rect 4706 16288 4714 16352
rect 4394 15264 4714 16288
rect 4394 15200 4402 15264
rect 4466 15200 4482 15264
rect 4546 15200 4562 15264
rect 4626 15200 4642 15264
rect 4706 15200 4714 15264
rect 4394 14176 4714 15200
rect 4394 14112 4402 14176
rect 4466 14112 4482 14176
rect 4546 14112 4562 14176
rect 4626 14112 4642 14176
rect 4706 14112 4714 14176
rect 4394 13088 4714 14112
rect 4394 13024 4402 13088
rect 4466 13024 4482 13088
rect 4546 13024 4562 13088
rect 4626 13024 4642 13088
rect 4706 13024 4714 13088
rect 4394 12582 4714 13024
rect 4394 12346 4436 12582
rect 4672 12346 4714 12582
rect 4394 12000 4714 12346
rect 4394 11936 4402 12000
rect 4466 11936 4482 12000
rect 4546 11936 4562 12000
rect 4626 11936 4642 12000
rect 4706 11936 4714 12000
rect 4394 10912 4714 11936
rect 4394 10848 4402 10912
rect 4466 10848 4482 10912
rect 4546 10848 4562 10912
rect 4626 10848 4642 10912
rect 4706 10848 4714 10912
rect 4394 9824 4714 10848
rect 4394 9760 4402 9824
rect 4466 9760 4482 9824
rect 4546 9760 4562 9824
rect 4626 9760 4642 9824
rect 4706 9760 4714 9824
rect 4394 8736 4714 9760
rect 4394 8672 4402 8736
rect 4466 8672 4482 8736
rect 4546 8672 4562 8736
rect 4626 8672 4642 8736
rect 4706 8672 4714 8736
rect 4394 7648 4714 8672
rect 4394 7584 4402 7648
rect 4466 7584 4482 7648
rect 4546 7584 4562 7648
rect 4626 7584 4642 7648
rect 4706 7584 4714 7648
rect 4394 6560 4714 7584
rect 4394 6496 4402 6560
rect 4466 6496 4482 6560
rect 4546 6496 4562 6560
rect 4626 6496 4642 6560
rect 4706 6496 4714 6560
rect 4394 5691 4714 6496
rect 4394 5472 4436 5691
rect 4672 5472 4714 5691
rect 4394 5408 4402 5472
rect 4466 5408 4482 5455
rect 4546 5408 4562 5455
rect 4626 5408 4642 5455
rect 4706 5408 4714 5472
rect 4394 4384 4714 5408
rect 4394 4320 4402 4384
rect 4466 4320 4482 4384
rect 4546 4320 4562 4384
rect 4626 4320 4642 4384
rect 4706 4320 4714 4384
rect 4394 3296 4714 4320
rect 4394 3232 4402 3296
rect 4466 3232 4482 3296
rect 4546 3232 4562 3296
rect 4626 3232 4642 3296
rect 4706 3232 4714 3296
rect 4394 2208 4714 3232
rect 4394 2144 4402 2208
rect 4466 2144 4482 2208
rect 4546 2144 4562 2208
rect 4626 2144 4642 2208
rect 4706 2144 4714 2208
rect 4394 2128 4714 2144
rect 7844 22336 8164 22896
rect 7844 22272 7852 22336
rect 7916 22272 7932 22336
rect 7996 22272 8012 22336
rect 8076 22272 8092 22336
rect 8156 22272 8164 22336
rect 7844 21248 8164 22272
rect 7844 21184 7852 21248
rect 7916 21184 7932 21248
rect 7996 21184 8012 21248
rect 8076 21184 8092 21248
rect 8156 21184 8164 21248
rect 7844 20160 8164 21184
rect 7844 20096 7852 20160
rect 7916 20096 7932 20160
rect 7996 20096 8012 20160
rect 8076 20096 8092 20160
rect 8156 20096 8164 20160
rect 7844 19072 8164 20096
rect 7844 19008 7852 19072
rect 7916 19008 7932 19072
rect 7996 19008 8012 19072
rect 8076 19008 8092 19072
rect 8156 19008 8164 19072
rect 7844 17984 8164 19008
rect 7844 17920 7852 17984
rect 7916 17920 7932 17984
rect 7996 17920 8012 17984
rect 8076 17920 8092 17984
rect 8156 17920 8164 17984
rect 7844 16896 8164 17920
rect 7844 16832 7852 16896
rect 7916 16832 7932 16896
rect 7996 16832 8012 16896
rect 8076 16832 8092 16896
rect 8156 16832 8164 16896
rect 7844 16027 8164 16832
rect 7844 15808 7886 16027
rect 8122 15808 8164 16027
rect 7844 15744 7852 15808
rect 7916 15744 7932 15791
rect 7996 15744 8012 15791
rect 8076 15744 8092 15791
rect 8156 15744 8164 15808
rect 7844 14720 8164 15744
rect 7844 14656 7852 14720
rect 7916 14656 7932 14720
rect 7996 14656 8012 14720
rect 8076 14656 8092 14720
rect 8156 14656 8164 14720
rect 7844 13632 8164 14656
rect 7844 13568 7852 13632
rect 7916 13568 7932 13632
rect 7996 13568 8012 13632
rect 8076 13568 8092 13632
rect 8156 13568 8164 13632
rect 7844 12544 8164 13568
rect 7844 12480 7852 12544
rect 7916 12480 7932 12544
rect 7996 12480 8012 12544
rect 8076 12480 8092 12544
rect 8156 12480 8164 12544
rect 7844 11456 8164 12480
rect 7844 11392 7852 11456
rect 7916 11392 7932 11456
rect 7996 11392 8012 11456
rect 8076 11392 8092 11456
rect 8156 11392 8164 11456
rect 7844 10368 8164 11392
rect 7844 10304 7852 10368
rect 7916 10304 7932 10368
rect 7996 10304 8012 10368
rect 8076 10304 8092 10368
rect 8156 10304 8164 10368
rect 7844 9280 8164 10304
rect 7844 9216 7852 9280
rect 7916 9216 7932 9280
rect 7996 9216 8012 9280
rect 8076 9216 8092 9280
rect 8156 9216 8164 9280
rect 7844 9136 8164 9216
rect 7844 8900 7886 9136
rect 8122 8900 8164 9136
rect 7844 8192 8164 8900
rect 7844 8128 7852 8192
rect 7916 8128 7932 8192
rect 7996 8128 8012 8192
rect 8076 8128 8092 8192
rect 8156 8128 8164 8192
rect 7844 7104 8164 8128
rect 7844 7040 7852 7104
rect 7916 7040 7932 7104
rect 7996 7040 8012 7104
rect 8076 7040 8092 7104
rect 8156 7040 8164 7104
rect 7844 6016 8164 7040
rect 7844 5952 7852 6016
rect 7916 5952 7932 6016
rect 7996 5952 8012 6016
rect 8076 5952 8092 6016
rect 8156 5952 8164 6016
rect 7844 4928 8164 5952
rect 7844 4864 7852 4928
rect 7916 4864 7932 4928
rect 7996 4864 8012 4928
rect 8076 4864 8092 4928
rect 8156 4864 8164 4928
rect 7844 3840 8164 4864
rect 7844 3776 7852 3840
rect 7916 3776 7932 3840
rect 7996 3776 8012 3840
rect 8076 3776 8092 3840
rect 8156 3776 8164 3840
rect 7844 2752 8164 3776
rect 7844 2688 7852 2752
rect 7916 2688 7932 2752
rect 7996 2688 8012 2752
rect 8076 2688 8092 2752
rect 8156 2688 8164 2752
rect 7844 2128 8164 2688
rect 11294 22880 11614 22896
rect 11294 22816 11302 22880
rect 11366 22816 11382 22880
rect 11446 22816 11462 22880
rect 11526 22816 11542 22880
rect 11606 22816 11614 22880
rect 11294 21792 11614 22816
rect 11294 21728 11302 21792
rect 11366 21728 11382 21792
rect 11446 21728 11462 21792
rect 11526 21728 11542 21792
rect 11606 21728 11614 21792
rect 11294 20704 11614 21728
rect 11294 20640 11302 20704
rect 11366 20640 11382 20704
rect 11446 20640 11462 20704
rect 11526 20640 11542 20704
rect 11606 20640 11614 20704
rect 11294 19616 11614 20640
rect 11294 19552 11302 19616
rect 11366 19552 11382 19616
rect 11446 19552 11462 19616
rect 11526 19552 11542 19616
rect 11606 19552 11614 19616
rect 11294 19472 11614 19552
rect 11294 19236 11336 19472
rect 11572 19236 11614 19472
rect 11294 18528 11614 19236
rect 11294 18464 11302 18528
rect 11366 18464 11382 18528
rect 11446 18464 11462 18528
rect 11526 18464 11542 18528
rect 11606 18464 11614 18528
rect 11294 17440 11614 18464
rect 11294 17376 11302 17440
rect 11366 17376 11382 17440
rect 11446 17376 11462 17440
rect 11526 17376 11542 17440
rect 11606 17376 11614 17440
rect 11294 16352 11614 17376
rect 11294 16288 11302 16352
rect 11366 16288 11382 16352
rect 11446 16288 11462 16352
rect 11526 16288 11542 16352
rect 11606 16288 11614 16352
rect 11294 15264 11614 16288
rect 11294 15200 11302 15264
rect 11366 15200 11382 15264
rect 11446 15200 11462 15264
rect 11526 15200 11542 15264
rect 11606 15200 11614 15264
rect 11294 14176 11614 15200
rect 11294 14112 11302 14176
rect 11366 14112 11382 14176
rect 11446 14112 11462 14176
rect 11526 14112 11542 14176
rect 11606 14112 11614 14176
rect 11294 13088 11614 14112
rect 11294 13024 11302 13088
rect 11366 13024 11382 13088
rect 11446 13024 11462 13088
rect 11526 13024 11542 13088
rect 11606 13024 11614 13088
rect 11294 12582 11614 13024
rect 11294 12346 11336 12582
rect 11572 12346 11614 12582
rect 11294 12000 11614 12346
rect 11294 11936 11302 12000
rect 11366 11936 11382 12000
rect 11446 11936 11462 12000
rect 11526 11936 11542 12000
rect 11606 11936 11614 12000
rect 11294 10912 11614 11936
rect 11294 10848 11302 10912
rect 11366 10848 11382 10912
rect 11446 10848 11462 10912
rect 11526 10848 11542 10912
rect 11606 10848 11614 10912
rect 11294 9824 11614 10848
rect 11294 9760 11302 9824
rect 11366 9760 11382 9824
rect 11446 9760 11462 9824
rect 11526 9760 11542 9824
rect 11606 9760 11614 9824
rect 11294 8736 11614 9760
rect 11294 8672 11302 8736
rect 11366 8672 11382 8736
rect 11446 8672 11462 8736
rect 11526 8672 11542 8736
rect 11606 8672 11614 8736
rect 11294 7648 11614 8672
rect 11294 7584 11302 7648
rect 11366 7584 11382 7648
rect 11446 7584 11462 7648
rect 11526 7584 11542 7648
rect 11606 7584 11614 7648
rect 11294 6560 11614 7584
rect 11294 6496 11302 6560
rect 11366 6496 11382 6560
rect 11446 6496 11462 6560
rect 11526 6496 11542 6560
rect 11606 6496 11614 6560
rect 11294 5691 11614 6496
rect 11294 5472 11336 5691
rect 11572 5472 11614 5691
rect 11294 5408 11302 5472
rect 11366 5408 11382 5455
rect 11446 5408 11462 5455
rect 11526 5408 11542 5455
rect 11606 5408 11614 5472
rect 11294 4384 11614 5408
rect 11294 4320 11302 4384
rect 11366 4320 11382 4384
rect 11446 4320 11462 4384
rect 11526 4320 11542 4384
rect 11606 4320 11614 4384
rect 11294 3296 11614 4320
rect 11294 3232 11302 3296
rect 11366 3232 11382 3296
rect 11446 3232 11462 3296
rect 11526 3232 11542 3296
rect 11606 3232 11614 3296
rect 11294 2208 11614 3232
rect 11294 2144 11302 2208
rect 11366 2144 11382 2208
rect 11446 2144 11462 2208
rect 11526 2144 11542 2208
rect 11606 2144 11614 2208
rect 11294 2128 11614 2144
rect 14744 22336 15064 22896
rect 14744 22272 14752 22336
rect 14816 22272 14832 22336
rect 14896 22272 14912 22336
rect 14976 22272 14992 22336
rect 15056 22272 15064 22336
rect 14744 21248 15064 22272
rect 14744 21184 14752 21248
rect 14816 21184 14832 21248
rect 14896 21184 14912 21248
rect 14976 21184 14992 21248
rect 15056 21184 15064 21248
rect 14744 20160 15064 21184
rect 14744 20096 14752 20160
rect 14816 20096 14832 20160
rect 14896 20096 14912 20160
rect 14976 20096 14992 20160
rect 15056 20096 15064 20160
rect 14744 19072 15064 20096
rect 14744 19008 14752 19072
rect 14816 19008 14832 19072
rect 14896 19008 14912 19072
rect 14976 19008 14992 19072
rect 15056 19008 15064 19072
rect 14744 17984 15064 19008
rect 14744 17920 14752 17984
rect 14816 17920 14832 17984
rect 14896 17920 14912 17984
rect 14976 17920 14992 17984
rect 15056 17920 15064 17984
rect 14744 16896 15064 17920
rect 14744 16832 14752 16896
rect 14816 16832 14832 16896
rect 14896 16832 14912 16896
rect 14976 16832 14992 16896
rect 15056 16832 15064 16896
rect 14744 16027 15064 16832
rect 14744 15808 14786 16027
rect 15022 15808 15064 16027
rect 14744 15744 14752 15808
rect 14816 15744 14832 15791
rect 14896 15744 14912 15791
rect 14976 15744 14992 15791
rect 15056 15744 15064 15808
rect 14744 14720 15064 15744
rect 14744 14656 14752 14720
rect 14816 14656 14832 14720
rect 14896 14656 14912 14720
rect 14976 14656 14992 14720
rect 15056 14656 15064 14720
rect 14744 13632 15064 14656
rect 14744 13568 14752 13632
rect 14816 13568 14832 13632
rect 14896 13568 14912 13632
rect 14976 13568 14992 13632
rect 15056 13568 15064 13632
rect 14744 12544 15064 13568
rect 14744 12480 14752 12544
rect 14816 12480 14832 12544
rect 14896 12480 14912 12544
rect 14976 12480 14992 12544
rect 15056 12480 15064 12544
rect 14744 11456 15064 12480
rect 14744 11392 14752 11456
rect 14816 11392 14832 11456
rect 14896 11392 14912 11456
rect 14976 11392 14992 11456
rect 15056 11392 15064 11456
rect 14744 10368 15064 11392
rect 14744 10304 14752 10368
rect 14816 10304 14832 10368
rect 14896 10304 14912 10368
rect 14976 10304 14992 10368
rect 15056 10304 15064 10368
rect 14744 9280 15064 10304
rect 14744 9216 14752 9280
rect 14816 9216 14832 9280
rect 14896 9216 14912 9280
rect 14976 9216 14992 9280
rect 15056 9216 15064 9280
rect 14744 9136 15064 9216
rect 14744 8900 14786 9136
rect 15022 8900 15064 9136
rect 14744 8192 15064 8900
rect 14744 8128 14752 8192
rect 14816 8128 14832 8192
rect 14896 8128 14912 8192
rect 14976 8128 14992 8192
rect 15056 8128 15064 8192
rect 14744 7104 15064 8128
rect 14744 7040 14752 7104
rect 14816 7040 14832 7104
rect 14896 7040 14912 7104
rect 14976 7040 14992 7104
rect 15056 7040 15064 7104
rect 14744 6016 15064 7040
rect 14744 5952 14752 6016
rect 14816 5952 14832 6016
rect 14896 5952 14912 6016
rect 14976 5952 14992 6016
rect 15056 5952 15064 6016
rect 14744 4928 15064 5952
rect 14744 4864 14752 4928
rect 14816 4864 14832 4928
rect 14896 4864 14912 4928
rect 14976 4864 14992 4928
rect 15056 4864 15064 4928
rect 14744 3840 15064 4864
rect 14744 3776 14752 3840
rect 14816 3776 14832 3840
rect 14896 3776 14912 3840
rect 14976 3776 14992 3840
rect 15056 3776 15064 3840
rect 14744 2752 15064 3776
rect 14744 2688 14752 2752
rect 14816 2688 14832 2752
rect 14896 2688 14912 2752
rect 14976 2688 14992 2752
rect 15056 2688 15064 2752
rect 14744 2128 15064 2688
rect 18194 22880 18514 22896
rect 18194 22816 18202 22880
rect 18266 22816 18282 22880
rect 18346 22816 18362 22880
rect 18426 22816 18442 22880
rect 18506 22816 18514 22880
rect 18194 21792 18514 22816
rect 18194 21728 18202 21792
rect 18266 21728 18282 21792
rect 18346 21728 18362 21792
rect 18426 21728 18442 21792
rect 18506 21728 18514 21792
rect 18194 20704 18514 21728
rect 18194 20640 18202 20704
rect 18266 20640 18282 20704
rect 18346 20640 18362 20704
rect 18426 20640 18442 20704
rect 18506 20640 18514 20704
rect 18194 19616 18514 20640
rect 18194 19552 18202 19616
rect 18266 19552 18282 19616
rect 18346 19552 18362 19616
rect 18426 19552 18442 19616
rect 18506 19552 18514 19616
rect 18194 19472 18514 19552
rect 18194 19236 18236 19472
rect 18472 19236 18514 19472
rect 18194 18528 18514 19236
rect 18194 18464 18202 18528
rect 18266 18464 18282 18528
rect 18346 18464 18362 18528
rect 18426 18464 18442 18528
rect 18506 18464 18514 18528
rect 18194 17440 18514 18464
rect 18194 17376 18202 17440
rect 18266 17376 18282 17440
rect 18346 17376 18362 17440
rect 18426 17376 18442 17440
rect 18506 17376 18514 17440
rect 18194 16352 18514 17376
rect 18194 16288 18202 16352
rect 18266 16288 18282 16352
rect 18346 16288 18362 16352
rect 18426 16288 18442 16352
rect 18506 16288 18514 16352
rect 18194 15264 18514 16288
rect 18194 15200 18202 15264
rect 18266 15200 18282 15264
rect 18346 15200 18362 15264
rect 18426 15200 18442 15264
rect 18506 15200 18514 15264
rect 18194 14176 18514 15200
rect 18194 14112 18202 14176
rect 18266 14112 18282 14176
rect 18346 14112 18362 14176
rect 18426 14112 18442 14176
rect 18506 14112 18514 14176
rect 18194 13088 18514 14112
rect 18194 13024 18202 13088
rect 18266 13024 18282 13088
rect 18346 13024 18362 13088
rect 18426 13024 18442 13088
rect 18506 13024 18514 13088
rect 18194 12582 18514 13024
rect 18194 12346 18236 12582
rect 18472 12346 18514 12582
rect 18194 12000 18514 12346
rect 18194 11936 18202 12000
rect 18266 11936 18282 12000
rect 18346 11936 18362 12000
rect 18426 11936 18442 12000
rect 18506 11936 18514 12000
rect 18194 10912 18514 11936
rect 18194 10848 18202 10912
rect 18266 10848 18282 10912
rect 18346 10848 18362 10912
rect 18426 10848 18442 10912
rect 18506 10848 18514 10912
rect 18194 9824 18514 10848
rect 18194 9760 18202 9824
rect 18266 9760 18282 9824
rect 18346 9760 18362 9824
rect 18426 9760 18442 9824
rect 18506 9760 18514 9824
rect 18194 8736 18514 9760
rect 18194 8672 18202 8736
rect 18266 8672 18282 8736
rect 18346 8672 18362 8736
rect 18426 8672 18442 8736
rect 18506 8672 18514 8736
rect 18194 7648 18514 8672
rect 18194 7584 18202 7648
rect 18266 7584 18282 7648
rect 18346 7584 18362 7648
rect 18426 7584 18442 7648
rect 18506 7584 18514 7648
rect 18194 6560 18514 7584
rect 18194 6496 18202 6560
rect 18266 6496 18282 6560
rect 18346 6496 18362 6560
rect 18426 6496 18442 6560
rect 18506 6496 18514 6560
rect 18194 5691 18514 6496
rect 18194 5472 18236 5691
rect 18472 5472 18514 5691
rect 18194 5408 18202 5472
rect 18266 5408 18282 5455
rect 18346 5408 18362 5455
rect 18426 5408 18442 5455
rect 18506 5408 18514 5472
rect 18194 4384 18514 5408
rect 18194 4320 18202 4384
rect 18266 4320 18282 4384
rect 18346 4320 18362 4384
rect 18426 4320 18442 4384
rect 18506 4320 18514 4384
rect 18194 3296 18514 4320
rect 18194 3232 18202 3296
rect 18266 3232 18282 3296
rect 18346 3232 18362 3296
rect 18426 3232 18442 3296
rect 18506 3232 18514 3296
rect 18194 2208 18514 3232
rect 18194 2144 18202 2208
rect 18266 2144 18282 2208
rect 18346 2144 18362 2208
rect 18426 2144 18442 2208
rect 18506 2144 18514 2208
rect 18194 2128 18514 2144
<< via4 >>
rect 4436 19236 4672 19472
rect 4436 12346 4672 12582
rect 4436 5472 4672 5691
rect 4436 5455 4466 5472
rect 4466 5455 4482 5472
rect 4482 5455 4546 5472
rect 4546 5455 4562 5472
rect 4562 5455 4626 5472
rect 4626 5455 4642 5472
rect 4642 5455 4672 5472
rect 7886 15808 8122 16027
rect 7886 15791 7916 15808
rect 7916 15791 7932 15808
rect 7932 15791 7996 15808
rect 7996 15791 8012 15808
rect 8012 15791 8076 15808
rect 8076 15791 8092 15808
rect 8092 15791 8122 15808
rect 7886 8900 8122 9136
rect 11336 19236 11572 19472
rect 11336 12346 11572 12582
rect 11336 5472 11572 5691
rect 11336 5455 11366 5472
rect 11366 5455 11382 5472
rect 11382 5455 11446 5472
rect 11446 5455 11462 5472
rect 11462 5455 11526 5472
rect 11526 5455 11542 5472
rect 11542 5455 11572 5472
rect 14786 15808 15022 16027
rect 14786 15791 14816 15808
rect 14816 15791 14832 15808
rect 14832 15791 14896 15808
rect 14896 15791 14912 15808
rect 14912 15791 14976 15808
rect 14976 15791 14992 15808
rect 14992 15791 15022 15808
rect 14786 8900 15022 9136
rect 18236 19236 18472 19472
rect 18236 12346 18472 12582
rect 18236 5472 18472 5691
rect 18236 5455 18266 5472
rect 18266 5455 18282 5472
rect 18282 5455 18346 5472
rect 18346 5455 18362 5472
rect 18362 5455 18426 5472
rect 18426 5455 18442 5472
rect 18442 5455 18472 5472
<< metal5 >>
rect 1104 19472 21804 19515
rect 1104 19236 4436 19472
rect 4672 19236 11336 19472
rect 11572 19236 18236 19472
rect 18472 19236 21804 19472
rect 1104 19194 21804 19236
rect 1104 16027 21804 16069
rect 1104 15791 7886 16027
rect 8122 15791 14786 16027
rect 15022 15791 21804 16027
rect 1104 15749 21804 15791
rect 1104 12582 21804 12624
rect 1104 12346 4436 12582
rect 4672 12346 11336 12582
rect 11572 12346 18236 12582
rect 18472 12346 21804 12582
rect 1104 12304 21804 12346
rect 1104 9136 21804 9179
rect 1104 8900 7886 9136
rect 8122 8900 14786 9136
rect 15022 8900 21804 9136
rect 1104 8858 21804 8900
rect 1104 5691 21804 5733
rect 1104 5455 4436 5691
rect 4672 5455 11336 5691
rect 11572 5455 18236 5691
rect 18472 5455 21804 5691
rect 1104 5413 21804 5455
use sky130_fd_sc_hd__fill_2  FILLER_0_6
timestamp 1619617919
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output45
timestamp 1619617919
transform -1 0 2208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1619617919
transform -1 0 1656 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1619617919
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1619617919
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1619617919
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1619617919
transform 1 0 3312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_18
timestamp 1619617919
transform 1 0 2760 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_6
timestamp 1619617919
transform 1 0 1656 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_12
timestamp 1619617919
transform 1 0 2208 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1619617919
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1619617919
transform -1 0 4140 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1619617919
transform -1 0 5796 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28
timestamp 1619617919
transform 1 0 3680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_33
timestamp 1619617919
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45
timestamp 1619617919
transform 1 0 5244 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_30
timestamp 1619617919
transform 1 0 3864 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_42
timestamp 1619617919
transform 1 0 4968 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_54
timestamp 1619617919
transform 1 0 6072 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1619617919
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1619617919
transform 1 0 6348 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51
timestamp 1619617919
transform 1 0 5796 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1619617919
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1619617919
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_70
timestamp 1619617919
transform 1 0 7544 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1619617919
transform -1 0 7268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_58
timestamp 1619617919
transform 1 0 6440 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_67
timestamp 1619617919
transform 1 0 7268 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _369_
timestamp 1619617919
transform -1 0 9108 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1619617919
transform 1 0 9752 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb1
timestamp 1619617919
transform 1 0 9108 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1619617919
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1619617919
transform -1 0 9016 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79
timestamp 1619617919
transform 1 0 8372 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86
timestamp 1619617919
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_88
timestamp 1619617919
transform 1 0 9200 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_97
timestamp 1619617919
transform 1 0 10028 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_105
timestamp 1619617919
transform 1 0 10764 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_107
timestamp 1619617919
transform 1 0 10948 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100
timestamp 1619617919
transform 1 0 10304 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1619617919
transform 1 0 10580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[11\].id.delayenb1
timestamp 1619617919
transform 1 0 10856 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_1_113
timestamp 1619617919
transform 1 0 11500 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1619617919
transform 1 0 11868 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115
timestamp 1619617919
transform 1 0 11684 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1619617919
transform -1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1619617919
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1619617919
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1619617919
transform 1 0 11684 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1619617919
transform 1 0 12512 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_121
timestamp 1619617919
transform 1 0 12236 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_127
timestamp 1619617919
transform 1 0 12788 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_133
timestamp 1619617919
transform 1 0 13340 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp 1619617919
transform -1 0 13892 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_149
timestamp 1619617919
transform 1 0 14812 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1619617919
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_137
timestamp 1619617919
transform 1 0 13708 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1619617919
transform 1 0 13800 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1619617919
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb1
timestamp 1619617919
transform 1 0 13892 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1619617919
transform 1 0 14536 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_146
timestamp 1619617919
transform 1 0 14536 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1619617919
transform 1 0 15548 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfrbp_2  idiv8
timestamp 1619617919
transform 1 0 16928 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb0
timestamp 1619617919
transform -1 0 15548 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1619617919
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  input1
timestamp 1619617919
transform 1 0 15640 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_170
timestamp 1619617919
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_166
timestamp 1619617919
transform 1 0 16376 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_170
timestamp 1619617919
transform 1 0 16744 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfrbp_1  idiv16
timestamp 1619617919
transform -1 0 21252 0 1 2720
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1619617919
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1619617919
transform 1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1619617919
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_179
timestamp 1619617919
transform 1 0 17572 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_191
timestamp 1619617919
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_196
timestamp 1619617919
transform 1 0 19136 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_204
timestamp 1619617919
transform 1 0 19872 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_202
timestamp 1619617919
transform 1 0 19688 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1619617919
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_212
timestamp 1619617919
transform 1 0 20608 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output43
timestamp 1619617919
transform -1 0 21068 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_217
timestamp 1619617919
transform 1 0 21068 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1619617919
transform 1 0 21252 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1619617919
transform -1 0 21528 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1619617919
transform -1 0 21804 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1619617919
transform -1 0 21804 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1619617919
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1619617919
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1619617919
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1619617919
transform 1 0 3864 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1619617919
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1619617919
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_34
timestamp 1619617919
transform 1 0 4232 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_46
timestamp 1619617919
transform 1 0 5336 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_4  irb
timestamp 1619617919
transform 1 0 6624 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_2_58
timestamp 1619617919
transform 1 0 6440 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1619617919
transform 1 0 7084 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen1
timestamp 1619617919
transform 1 0 8464 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1619617919
transform -1 0 9384 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1619617919
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_77
timestamp 1619617919
transform 1 0 8188 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1619617919
transform 1 0 8924 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_90
timestamp 1619617919
transform 1 0 9384 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1619617919
transform 1 0 11684 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[11\].id.delayen1
timestamp 1619617919
transform 1 0 10948 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1619617919
transform 1 0 11408 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_102
timestamp 1619617919
transform 1 0 10488 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_106
timestamp 1619617919
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_118
timestamp 1619617919
transform 1 0 11960 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen1
timestamp 1619617919
transform 1 0 13524 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1619617919
transform 1 0 14812 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1619617919
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_130
timestamp 1619617919
transform 1 0 13064 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_134
timestamp 1619617919
transform 1 0 13432 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_140
timestamp 1619617919
transform 1 0 13984 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_144
timestamp 1619617919
transform 1 0 14352 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_148
timestamp 1619617919
transform 1 0 14720 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen0
timestamp 1619617919
transform -1 0 15548 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_2_157
timestamp 1619617919
transform 1 0 15548 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_169
timestamp 1619617919
transform 1 0 16652 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_181
timestamp 1619617919
transform 1 0 17756 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_193
timestamp 1619617919
transform 1 0 18860 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1619617919
transform -1 0 21804 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1619617919
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_199
timestamp 1619617919
transform 1 0 19412 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_201
timestamp 1619617919
transform 1 0 19596 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_213
timestamp 1619617919
transform 1 0 20700 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_221
timestamp 1619617919
transform 1 0 21436 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1619617919
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1619617919
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1619617919
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1619617919
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1619617919
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1619617919
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1619617919
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1619617919
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1619617919
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_82
timestamp 1619617919
transform 1 0 8648 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_94
timestamp 1619617919
transform 1 0 9752 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1619617919
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_106
timestamp 1619617919
transform 1 0 10856 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_115
timestamp 1619617919
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_127
timestamp 1619617919
transform 1 0 12788 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_139
timestamp 1619617919
transform 1 0 13892 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1619617919
transform -1 0 15732 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1619617919
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_151
timestamp 1619617919
transform 1 0 14996 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1619617919
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_172
timestamp 1619617919
transform 1 0 16928 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1619617919
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1619617919
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1619617919
transform -1 0 21804 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1619617919
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_220
timestamp 1619617919
transform 1 0 21344 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1619617919
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1619617919
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1619617919
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrbp_2  idiv4
timestamp 1619617919
transform -1 0 7084 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1619617919
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1619617919
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_30
timestamp 1619617919
transform 1 0 3864 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_38
timestamp 1619617919
transform 1 0 4600 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _368_
timestamp 1619617919
transform 1 0 7820 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_65
timestamp 1619617919
transform 1 0 7084 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _356_
timestamp 1619617919
transform -1 0 10304 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1619617919
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_82
timestamp 1619617919
transform 1 0 8648 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1619617919
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_4  ringosc.dstage\[11\].id.delayen0
timestamp 1619617919
transform 1 0 10488 0 -1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_4_100
timestamp 1619617919
transform 1 0 10304 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_113
timestamp 1619617919
transform 1 0 11500 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1619617919
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_125
timestamp 1619617919
transform 1 0 12604 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_137
timestamp 1619617919
transform 1 0 13708 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144
timestamp 1619617919
transform 1 0 14352 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_156
timestamp 1619617919
transform 1 0 15456 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_168
timestamp 1619617919
transform 1 0 16560 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1619617919
transform 1 0 17940 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_180
timestamp 1619617919
transform 1 0 17664 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_192
timestamp 1619617919
transform 1 0 18768 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1619617919
transform -1 0 21804 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1619617919
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_201
timestamp 1619617919
transform 1 0 19596 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_213
timestamp 1619617919
transform 1 0 20700 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_221
timestamp 1619617919
transform 1 0 21436 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfrbp_2  idiv2
timestamp 1619617919
transform 1 0 2944 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1619617919
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1619617919
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1619617919
transform 1 0 2484 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_19
timestamp 1619617919
transform 1 0 2852 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1619617919
transform 1 0 5152 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb0
timestamp 1619617919
transform 1 0 7544 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1619617919
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_56
timestamp 1619617919
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1619617919
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen0
timestamp 1619617919
transform 1 0 8188 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_5_82
timestamp 1619617919
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_94
timestamp 1619617919
transform 1 0 9752 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb0
timestamp 1619617919
transform 1 0 12420 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1619617919
transform -1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb0
timestamp 1619617919
transform 1 0 10304 0 1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1619617919
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_111
timestamp 1619617919
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_115
timestamp 1619617919
transform 1 0 11684 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen0
timestamp 1619617919
transform 1 0 13064 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1619617919
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_135
timestamp 1619617919
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_143
timestamp 1619617919
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_149
timestamp 1619617919
transform 1 0 14812 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1619617919
transform 1 0 16928 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1619617919
transform 1 0 15088 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1619617919
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_155
timestamp 1619617919
transform 1 0 15364 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_167
timestamp 1619617919
transform 1 0 16468 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1619617919
transform -1 0 18216 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1619617919
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_186
timestamp 1619617919
transform 1 0 18216 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_198
timestamp 1619617919
transform 1 0 19320 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1619617919
transform -1 0 21804 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_210
timestamp 1619617919
transform 1 0 20424 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_7
timestamp 1619617919
transform 1 0 1748 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output41
timestamp 1619617919
transform -1 0 1748 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1619617919
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1619617919
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_23
timestamp 1619617919
transform 1 0 3220 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_15
timestamp 1619617919
transform 1 0 2484 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_19
timestamp 1619617919
transform 1 0 2852 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_15
timestamp 1619617919
transform 1 0 2484 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  ringosc.ibufp11
timestamp 1619617919
transform -1 0 2852 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  ringosc.ibufp10
timestamp 1619617919
transform -1 0 3588 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1619617919
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[5\].id.delayenb1
timestamp 1619617919
transform -1 0 6164 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1619617919
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1619617919
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1619617919
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1619617919
transform 1 0 4968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1619617919
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_39
timestamp 1619617919
transform 1 0 4692 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_47
timestamp 1619617919
transform 1 0 5428 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1619617919
transform -1 0 7176 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1619617919
transform 1 0 6900 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[5\].id.delayen1
timestamp 1619617919
transform 1 0 6440 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1619617919
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_54
timestamp 1619617919
transform 1 0 6072 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_66
timestamp 1619617919
transform 1 0 7176 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_55
timestamp 1619617919
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_66
timestamp 1619617919
transform 1 0 7176 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1619617919
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_78
timestamp 1619617919
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_87
timestamp 1619617919
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_99
timestamp 1619617919
transform 1 0 10212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_78
timestamp 1619617919
transform 1 0 8280 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_90
timestamp 1619617919
transform 1 0 9384 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1619617919
transform -1 0 12880 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1619617919
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_111
timestamp 1619617919
transform 1 0 11316 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_123
timestamp 1619617919
transform 1 0 12420 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_102
timestamp 1619617919
transform 1 0 10488 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_115
timestamp 1619617919
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb1
timestamp 1619617919
transform -1 0 15180 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1619617919
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_128
timestamp 1619617919
transform 1 0 12880 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_140
timestamp 1619617919
transform 1 0 13984 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_144
timestamp 1619617919
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1619617919
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_139
timestamp 1619617919
transform 1 0 13892 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1619617919
transform 1 0 16100 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen1
timestamp 1619617919
transform -1 0 15640 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1619617919
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_158
timestamp 1619617919
transform 1 0 15640 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_162
timestamp 1619617919
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_172
timestamp 1619617919
transform 1 0 16928 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_151
timestamp 1619617919
transform 1 0 14996 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_163
timestamp 1619617919
transform 1 0 16100 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_172
timestamp 1619617919
transform 1 0 16928 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1619617919
transform -1 0 19136 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _322_
timestamp 1619617919
transform -1 0 17940 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _323_
timestamp 1619617919
transform 1 0 17388 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _324_
timestamp 1619617919
transform -1 0 18860 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _325_
timestamp 1619617919
transform -1 0 18676 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_176
timestamp 1619617919
transform 1 0 17296 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_196
timestamp 1619617919
transform 1 0 19136 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_191
timestamp 1619617919
transform 1 0 18676 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1619617919
transform -1 0 21804 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1619617919
transform -1 0 21804 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1619617919
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1619617919
transform -1 0 21528 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_201
timestamp 1619617919
transform 1 0 19596 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_213
timestamp 1619617919
transform 1 0 20700 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_203
timestamp 1619617919
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_215
timestamp 1619617919
transform 1 0 20884 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_221
timestamp 1619617919
transform 1 0 21436 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1619617919
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1619617919
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1619617919
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1619617919
transform 1 0 5244 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb0
timestamp 1619617919
transform 1 0 4232 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1619617919
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1619617919
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_30
timestamp 1619617919
transform 1 0 3864 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1619617919
transform -1 0 8740 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1619617919
transform -1 0 6164 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_55
timestamp 1619617919
transform 1 0 6164 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_67
timestamp 1619617919
transform 1 0 7268 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_73
timestamp 1619617919
transform 1 0 7820 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.iss.delayenb1
timestamp 1619617919
transform 1 0 9844 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1619617919
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_83
timestamp 1619617919
transform 1 0 8740 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_87
timestamp 1619617919
transform 1 0 9108 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1619617919
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.delayen1
timestamp 1619617919
transform 1 0 10488 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_8_110
timestamp 1619617919
transform 1 0 11224 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_122
timestamp 1619617919
transform 1 0 12328 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1619617919
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_134
timestamp 1619617919
transform 1 0 13432 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_142
timestamp 1619617919
transform 1 0 14168 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1619617919
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1619617919
transform 1 0 15548 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_156
timestamp 1619617919
transform 1 0 15456 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1619617919
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1619617919
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_190
timestamp 1619617919
transform 1 0 18584 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_198
timestamp 1619617919
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1619617919
transform -1 0 21804 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1619617919
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_201
timestamp 1619617919
transform 1 0 19596 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_213
timestamp 1619617919
transform 1 0 20700 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_221
timestamp 1619617919
transform 1 0 21436 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1619617919
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1619617919
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1619617919
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1619617919
transform -1 0 4048 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1619617919
transform 1 0 3588 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_32
timestamp 1619617919
transform 1 0 4048 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_44
timestamp 1619617919
transform 1 0 5152 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00
timestamp 1619617919
transform -1 0 7912 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1619617919
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_56
timestamp 1619617919
transform 1 0 6256 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1619617919
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_74
timestamp 1619617919
transform 1 0 7912 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.delayen0
timestamp 1619617919
transform 1 0 8556 0 1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb0
timestamp 1619617919
transform 1 0 9660 0 1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_9_80
timestamp 1619617919
transform 1 0 8464 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_92
timestamp 1619617919
transform 1 0 9568 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb0
timestamp 1619617919
transform 1 0 12236 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1619617919
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_104
timestamp 1619617919
transform 1 0 10672 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_112
timestamp 1619617919
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_115
timestamp 1619617919
transform 1 0 11684 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen0
timestamp 1619617919
transform 1 0 12880 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1619617919
transform -1 0 14352 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_133
timestamp 1619617919
transform 1 0 13340 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_144
timestamp 1619617919
transform 1 0 14352 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1619617919
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_156
timestamp 1619617919
transform 1 0 15456 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_168
timestamp 1619617919
transform 1 0 16560 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_172
timestamp 1619617919
transform 1 0 16928 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1619617919
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1619617919
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1619617919
transform -1 0 21804 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1619617919
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_220
timestamp 1619617919
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb0
timestamp 1619617919
transform 1 0 2116 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1619617919
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1619617919
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_18
timestamp 1619617919
transform 1 0 2760 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1619617919
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_26
timestamp 1619617919
transform 1 0 3496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1619617919
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1619617919
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01
timestamp 1619617919
transform -1 0 8096 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_10_54
timestamp 1619617919
transform 1 0 6072 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_62
timestamp 1619617919
transform 1 0 6808 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0
timestamp 1619617919
transform -1 0 8648 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1619617919
transform -1 0 9936 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1619617919
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_76
timestamp 1619617919
transform 1 0 8096 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_82
timestamp 1619617919
transform 1 0 8648 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_87
timestamp 1619617919
transform 1 0 9108 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_96
timestamp 1619617919
transform 1 0 9936 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1619617919
transform 1 0 12420 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_108
timestamp 1619617919
transform 1 0 11040 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_120
timestamp 1619617919
transform 1 0 12144 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb1
timestamp 1619617919
transform -1 0 14996 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1619617919
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_132
timestamp 1619617919
transform 1 0 13248 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_140
timestamp 1619617919
transform 1 0 13984 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1619617919
transform -1 0 16560 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1619617919
transform 1 0 15456 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen1
timestamp 1619617919
transform 1 0 14996 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_10_159
timestamp 1619617919
transform 1 0 15732 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_163
timestamp 1619617919
transform 1 0 16100 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_168
timestamp 1619617919
transform 1 0 16560 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_180
timestamp 1619617919
transform 1 0 17664 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_192
timestamp 1619617919
transform 1 0 18768 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1619617919
transform -1 0 21804 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1619617919
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1619617919
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_213
timestamp 1619617919
transform 1 0 20700 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_221
timestamp 1619617919
transform 1 0 21436 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _360_
timestamp 1619617919
transform 1 0 2116 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1619617919
transform 1 0 2944 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1619617919
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1619617919
transform -1 0 1656 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_6
timestamp 1619617919
transform 1 0 1656 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_10
timestamp 1619617919
transform 1 0 2024 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1619617919
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1619617919
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _372_
timestamp 1619617919
transform -1 0 7268 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.reseten0
timestamp 1619617919
transform 1 0 7544 0 1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1619617919
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_51
timestamp 1619617919
transform 1 0 5796 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_67
timestamp 1619617919
transform 1 0 7268 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1
timestamp 1619617919
transform 1 0 8556 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_84
timestamp 1619617919
transform 1 0 8832 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_96
timestamp 1619617919
transform 1 0 9936 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _291_
timestamp 1619617919
transform 1 0 11868 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1619617919
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_108
timestamp 1619617919
transform 1 0 11040 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1619617919
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_122
timestamp 1619617919
transform 1 0 12328 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_134
timestamp 1619617919
transform 1 0 13432 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_146
timestamp 1619617919
transform 1 0 14536 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen0
timestamp 1619617919
transform 1 0 16928 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb0
timestamp 1619617919
transform 1 0 16192 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1619617919
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_158
timestamp 1619617919
transform 1 0 15640 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1619617919
transform 1 0 19228 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen1
timestamp 1619617919
transform 1 0 18768 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb1
timestamp 1619617919
transform -1 0 18768 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_11_177
timestamp 1619617919
transform 1 0 17388 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1619617919
transform -1 0 21804 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1619617919
transform 1 0 21252 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_200
timestamp 1619617919
transform 1 0 19504 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_212
timestamp 1619617919
transform 1 0 20608 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_218
timestamp 1619617919
transform 1 0 21160 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1619617919
transform 1 0 2668 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1619617919
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1619617919
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_15
timestamp 1619617919
transform 1 0 2484 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1619617919
transform 1 0 2944 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _303_
timestamp 1619617919
transform 1 0 4508 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1619617919
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_28
timestamp 1619617919
transform 1 0 3680 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_30
timestamp 1619617919
transform 1 0 3864 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_36
timestamp 1619617919
transform 1 0 4416 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_43
timestamp 1619617919
transform 1 0 5060 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _196_
timestamp 1619617919
transform 1 0 6624 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_12_55
timestamp 1619617919
transform 1 0 6164 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_59
timestamp 1619617919
transform 1 0 6532 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_67
timestamp 1619617919
transform 1 0 7268 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_1  _306_
timestamp 1619617919
transform 1 0 9476 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1619617919
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_79
timestamp 1619617919
transform 1 0 8372 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1619617919
transform 1 0 8924 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1619617919
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_96
timestamp 1619617919
transform 1 0 9936 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0
timestamp 1619617919
transform 1 0 11408 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_108
timestamp 1619617919
transform 1 0 11040 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_116
timestamp 1619617919
transform 1 0 11776 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _347_
timestamp 1619617919
transform -1 0 14628 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1619617919
transform 1 0 14812 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1619617919
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_128
timestamp 1619617919
transform 1 0 12880 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_140
timestamp 1619617919
transform 1 0 13984 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_147
timestamp 1619617919
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1619617919
transform 1 0 16652 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_158
timestamp 1619617919
transform 1 0 15640 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_166
timestamp 1619617919
transform 1 0 16376 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_173
timestamp 1619617919
transform 1 0 17020 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1619617919
transform -1 0 18492 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_185
timestamp 1619617919
transform 1 0 18124 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_189
timestamp 1619617919
transform 1 0 18492 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_197
timestamp 1619617919
transform 1 0 19228 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1619617919
transform -1 0 21804 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1619617919
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1619617919
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_213
timestamp 1619617919
transform 1 0 20700 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_221
timestamp 1619617919
transform 1 0 21436 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1619617919
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output39
timestamp 1619617919
transform -1 0 1748 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1619617919
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1619617919
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb1
timestamp 1619617919
transform 1 0 1748 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp 1619617919
transform 1 0 2852 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen1
timestamp 1619617919
transform 1 0 2392 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1619617919
transform 1 0 2852 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_7
timestamp 1619617919
transform 1 0 1748 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_22
timestamp 1619617919
transform 1 0 3128 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _354_
timestamp 1619617919
transform -1 0 5888 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _377_
timestamp 1619617919
transform -1 0 5428 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1619617919
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_34
timestamp 1619617919
transform 1 0 4232 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1619617919
transform 1 0 5428 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1619617919
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1619617919
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_42
timestamp 1619617919
transform 1 0 4968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_8  _197_
timestamp 1619617919
transform -1 0 8832 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1619617919
transform 1 0 5888 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1619617919
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_55
timestamp 1619617919
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_58
timestamp 1619617919
transform 1 0 6440 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_66
timestamp 1619617919
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_61
timestamp 1619617919
transform 1 0 6716 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_73
timestamp 1619617919
transform 1 0 7820 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _312_
timestamp 1619617919
transform -1 0 10488 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _321_
timestamp 1619617919
transform 1 0 10212 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1619617919
transform -1 0 10212 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1619617919
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  repeater46
timestamp 1619617919
transform -1 0 9936 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_13_84
timestamp 1619617919
transform 1 0 8832 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1619617919
transform 1 0 8924 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen1
timestamp 1619617919
transform 1 0 12328 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb1
timestamp 1619617919
transform 1 0 11684 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1619617919
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_105
timestamp 1619617919
transform 1 0 10764 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1619617919
transform 1 0 11500 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_102
timestamp 1619617919
transform 1 0 10488 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_114
timestamp 1619617919
transform 1 0 11592 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_126
timestamp 1619617919
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 1619617919
transform 1 0 13524 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb0
timestamp 1619617919
transform 1 0 12880 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1619617919
transform 1 0 12788 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_142
timestamp 1619617919
transform 1 0 14168 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_138
timestamp 1619617919
transform 1 0 13800 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1619617919
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_144
timestamp 1619617919
transform 1 0 14352 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_142
timestamp 1619617919
transform 1 0 14168 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_130
timestamp 1619617919
transform 1 0 13064 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1619617919
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_154
timestamp 1619617919
transform 1 0 15272 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_166
timestamp 1619617919
transform 1 0 16376 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_170
timestamp 1619617919
transform 1 0 16744 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1619617919
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_156
timestamp 1619617919
transform 1 0 15456 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_168
timestamp 1619617919
transform 1 0 16560 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1619617919
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1619617919
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_180
timestamp 1619617919
transform 1 0 17664 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_192
timestamp 1619617919
transform 1 0 18768 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1619617919
transform -1 0 21804 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1619617919
transform -1 0 21804 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1619617919
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1619617919
transform 1 0 21252 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1619617919
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_220
timestamp 1619617919
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1619617919
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_213
timestamp 1619617919
transform 1 0 20700 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1619617919
transform 1 0 2576 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1619617919
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1619617919
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_15
timestamp 1619617919
transform 1 0 2484 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_20
timestamp 1619617919
transform 1 0 2944 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _314_
timestamp 1619617919
transform 1 0 4600 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_32
timestamp 1619617919
transform 1 0 4048 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1619617919
transform 1 0 5152 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1619617919
transform -1 0 8096 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _307_
timestamp 1619617919
transform 1 0 6440 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1619617919
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_56
timestamp 1619617919
transform 1 0 6256 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_65
timestamp 1619617919
transform 1 0 7084 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1619617919
transform 1 0 9476 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _319_
timestamp 1619617919
transform 1 0 8924 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_76
timestamp 1619617919
transform 1 0 8096 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_84
timestamp 1619617919
transform 1 0 8832 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_94
timestamp 1619617919
transform 1 0 9752 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1619617919
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_106
timestamp 1619617919
transform 1 0 10856 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_115
timestamp 1619617919
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen0
timestamp 1619617919
transform 1 0 13064 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb0
timestamp 1619617919
transform 1 0 14812 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_15_127
timestamp 1619617919
transform 1 0 12788 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1619617919
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_147
timestamp 1619617919
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen0
timestamp 1619617919
transform 1 0 15732 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1619617919
transform -1 0 17204 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1619617919
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_156
timestamp 1619617919
transform 1 0 15456 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_164
timestamp 1619617919
transform 1 0 16192 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_170
timestamp 1619617919
transform 1 0 16744 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp 1619617919
transform 1 0 17664 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _385_
timestamp 1619617919
transform 1 0 19136 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1619617919
transform 1 0 18492 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen1
timestamp 1619617919
transform -1 0 17664 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_15_192
timestamp 1619617919
transform 1 0 18768 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1619617919
transform -1 0 21804 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_217
timestamp 1619617919
transform 1 0 21068 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_221
timestamp 1619617919
transform 1 0 21436 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1619617919
transform -1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb1
timestamp 1619617919
transform -1 0 3588 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1619617919
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1619617919
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_14
timestamp 1619617919
transform 1 0 2392 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1619617919
transform 1 0 4324 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen1
timestamp 1619617919
transform 1 0 3864 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1619617919
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1619617919
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_38
timestamp 1619617919
transform 1 0 4600 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1619617919
transform 1 0 6900 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 7544 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _302_
timestamp 1619617919
transform 1 0 7176 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_50
timestamp 1619617919
transform 1 0 5704 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_62
timestamp 1619617919
transform 1 0 6808 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _300_
timestamp 1619617919
transform -1 0 8556 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _315_
timestamp 1619617919
transform 1 0 10028 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1619617919
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_81
timestamp 1619617919
transform 1 0 8556 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1619617919
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_87
timestamp 1619617919
transform 1 0 9108 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_95
timestamp 1619617919
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_2  _365_
timestamp 1619617919
transform 1 0 11224 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_102
timestamp 1619617919
transform 1 0 10488 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_119
timestamp 1619617919
transform 1 0 12052 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1619617919
transform -1 0 13432 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1619617919
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_134
timestamp 1619617919
transform 1 0 13432 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_142
timestamp 1619617919
transform 1 0 14168 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_144
timestamp 1619617919
transform 1 0 14352 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1619617919
transform 1 0 14904 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1619617919
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_166
timestamp 1619617919
transform 1 0 16376 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _373_
timestamp 1619617919
transform -1 0 18860 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb1
timestamp 1619617919
transform -1 0 17848 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_16_174
timestamp 1619617919
transform 1 0 17112 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_182
timestamp 1619617919
transform 1 0 17848 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_193
timestamp 1619617919
transform 1 0 18860 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1619617919
transform -1 0 20332 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1619617919
transform -1 0 21804 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1619617919
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_199
timestamp 1619617919
transform 1 0 19412 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_201
timestamp 1619617919
transform 1 0 19596 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_205
timestamp 1619617919
transform 1 0 19964 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1619617919
transform 1 0 20332 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_221
timestamp 1619617919
transform 1 0 21436 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1619617919
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1619617919
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1619617919
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _308_
timestamp 1619617919
transform 1 0 5428 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1619617919
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_39
timestamp 1619617919
transform 1 0 4692 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _296_
timestamp 1619617919
transform -1 0 6900 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _298_
timestamp 1619617919
transform -1 0 8464 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1619617919
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_54
timestamp 1619617919
transform 1 0 6072 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_63
timestamp 1619617919
transform 1 0 6900 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_71
timestamp 1619617919
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _311_
timestamp 1619617919
transform 1 0 9292 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _317_
timestamp 1619617919
transform -1 0 10672 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_80
timestamp 1619617919
transform 1 0 8464 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_88
timestamp 1619617919
transform 1 0 9200 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1619617919
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_104
timestamp 1619617919
transform 1 0 10672 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_112
timestamp 1619617919
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_115
timestamp 1619617919
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_127
timestamp 1619617919
transform 1 0 12788 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_139
timestamp 1619617919
transform 1 0 13892 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1619617919
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_151
timestamp 1619617919
transform 1 0 14996 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_163
timestamp 1619617919
transform 1 0 16100 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_172
timestamp 1619617919
transform 1 0 16928 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1619617919
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1619617919
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1619617919
transform -1 0 21804 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1619617919
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_220
timestamp 1619617919
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1619617919
transform -1 0 3588 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1619617919
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1619617919
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_15
timestamp 1619617919
transform 1 0 2484 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_23
timestamp 1619617919
transform 1 0 3220 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _366_
timestamp 1619617919
transform 1 0 4968 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1619617919
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1619617919
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1619617919
transform 1 0 3864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _304_
timestamp 1619617919
transform 1 0 5796 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_18_58
timestamp 1619617919
transform 1 0 6440 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_70
timestamp 1619617919
transform 1 0 7544 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1619617919
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_82
timestamp 1619617919
transform 1 0 8648 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1619617919
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_99
timestamp 1619617919
transform 1 0 10212 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _318_
timestamp 1619617919
transform 1 0 11592 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_18_111
timestamp 1619617919
transform 1 0 11316 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_119
timestamp 1619617919
transform 1 0 12052 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _401_
timestamp 1619617919
transform -1 0 16192 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1619617919
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_131
timestamp 1619617919
transform 1 0 13156 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_164
timestamp 1619617919
transform 1 0 16192 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_176
timestamp 1619617919
transform 1 0 17296 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_188
timestamp 1619617919
transform 1 0 18400 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1619617919
transform -1 0 21804 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1619617919
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_201
timestamp 1619617919
transform 1 0 19596 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_213
timestamp 1619617919
transform 1 0 20700 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_221
timestamp 1619617919
transform 1 0 21436 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1619617919
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_7
timestamp 1619617919
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output40
timestamp 1619617919
transform -1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1619617919
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1619617919
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb0
timestamp 1619617919
transform 1 0 2116 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _364_
timestamp 1619617919
transform -1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_14
timestamp 1619617919
transform 1 0 2392 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1619617919
transform 1 0 3128 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen0
timestamp 1619617919
transform 1 0 2760 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_19_23
timestamp 1619617919
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_1  _293_
timestamp 1619617919
transform -1 0 5336 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1619617919
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_35
timestamp 1619617919
transform 1 0 4324 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_46
timestamp 1619617919
transform 1 0 5336 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_26
timestamp 1619617919
transform 1 0 3496 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1619617919
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_42
timestamp 1619617919
transform 1 0 4968 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_54
timestamp 1619617919
transform 1 0 6072 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1619617919
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _248_
timestamp 1619617919
transform 1 0 6440 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_20_70
timestamp 1619617919
transform 1 0 7544 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_66
timestamp 1619617919
transform 1 0 7176 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_69
timestamp 1619617919
transform 1 0 7452 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_63
timestamp 1619617919
transform 1 0 6900 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _254_
timestamp 1619617919
transform 1 0 7544 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1619617919
transform 1 0 7268 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_54
timestamp 1619617919
transform 1 0 6072 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_80
timestamp 1619617919
transform 1 0 8464 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_76
timestamp 1619617919
transform 1 0 8096 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_82
timestamp 1619617919
transform 1 0 8648 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1619617919
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _310_
timestamp 1619617919
transform -1 0 8648 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1619617919
transform 1 0 8188 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _316_
timestamp 1619617919
transform -1 0 10488 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _309_
timestamp 1619617919
transform 1 0 9200 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_20_99
timestamp 1619617919
transform 1 0 10212 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_87
timestamp 1619617919
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_102
timestamp 1619617919
transform 1 0 10488 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _313_
timestamp 1619617919
transform -1 0 11040 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _290_
timestamp 1619617919
transform 1 0 11040 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_20_117
timestamp 1619617919
transform 1 0 11868 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_111
timestamp 1619617919
transform 1 0 11316 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1619617919
transform 1 0 11500 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1619617919
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1619617919
transform 1 0 11684 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _371_
timestamp 1619617919
transform -1 0 12788 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_124
timestamp 1619617919
transform 1 0 12512 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _199_
timestamp 1619617919
transform -1 0 14996 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _292_
timestamp 1619617919
transform 1 0 12788 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1619617919
transform -1 0 14996 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1619617919
transform 1 0 12880 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1619617919
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_137
timestamp 1619617919
transform 1 0 13708 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_145
timestamp 1619617919
transform 1 0 14444 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_132
timestamp 1619617919
transform 1 0 13248 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_140
timestamp 1619617919
transform 1 0 13984 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _341_
timestamp 1619617919
transform 1 0 16560 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _386_
timestamp 1619617919
transform -1 0 17756 0 -1 13600
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1619617919
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_151
timestamp 1619617919
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_163
timestamp 1619617919
transform 1 0 16100 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1619617919
transform 1 0 16468 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_172
timestamp 1619617919
transform 1 0 16928 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_151
timestamp 1619617919
transform 1 0 14996 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_157
timestamp 1619617919
transform 1 0 15548 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1619617919
transform 1 0 17296 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _286_
timestamp 1619617919
transform 1 0 17756 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _287_
timestamp 1619617919
transform -1 0 19320 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _288_
timestamp 1619617919
transform 1 0 18860 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_19_179
timestamp 1619617919
transform 1 0 17572 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_191
timestamp 1619617919
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_198
timestamp 1619617919
transform 1 0 19320 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_188
timestamp 1619617919
transform 1 0 18400 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_198
timestamp 1619617919
transform 1 0 19320 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _200_
timestamp 1619617919
transform 1 0 19596 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1619617919
transform -1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _400_
timestamp 1619617919
transform 1 0 19688 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1619617919
transform -1 0 21804 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1619617919
transform -1 0 21804 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1619617919
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1619617919
transform -1 0 21528 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_208
timestamp 1619617919
transform 1 0 20240 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1619617919
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1619617919
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1619617919
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1619617919
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1619617919
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1619617919
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1619617919
transform 1 0 7728 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1619617919
transform 1 0 6072 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _294_
timestamp 1619617919
transform 1 0 7268 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _305_
timestamp 1619617919
transform 1 0 6440 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1619617919
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_51
timestamp 1619617919
transform 1 0 5796 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_65
timestamp 1619617919
transform 1 0 7084 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1619617919
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _320_
timestamp 1619617919
transform -1 0 10304 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_78
timestamp 1619617919
transform 1 0 8280 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_90
timestamp 1619617919
transform 1 0 9384 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1619617919
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_100
timestamp 1619617919
transform 1 0 10304 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_112
timestamp 1619617919
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_115
timestamp 1619617919
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1619617919
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1619617919
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1619617919
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_151
timestamp 1619617919
transform 1 0 14996 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_163
timestamp 1619617919
transform 1 0 16100 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_172
timestamp 1619617919
transform 1 0 16928 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1619617919
transform 1 0 18768 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _279_
timestamp 1619617919
transform -1 0 17940 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _285_
timestamp 1619617919
transform -1 0 18308 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_187
timestamp 1619617919
transform 1 0 18308 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_191
timestamp 1619617919
transform 1 0 18676 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_195
timestamp 1619617919
transform 1 0 19044 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1619617919
transform -1 0 21804 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_207
timestamp 1619617919
transform 1 0 20148 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_219
timestamp 1619617919
transform 1 0 21252 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1619617919
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1619617919
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1619617919
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _392_
timestamp 1619617919
transform -1 0 5980 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1619617919
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1619617919
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_30
timestamp 1619617919
transform 1 0 3864 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1619617919
transform 1 0 5980 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1619617919
transform 1 0 7084 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1619617919
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_77
timestamp 1619617919
transform 1 0 8188 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1619617919
transform 1 0 8924 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_87
timestamp 1619617919
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1619617919
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_4  _194_
timestamp 1619617919
transform 1 0 12328 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_22_111
timestamp 1619617919
transform 1 0 11316 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_119
timestamp 1619617919
transform 1 0 12052 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _212_
timestamp 1619617919
transform 1 0 14536 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1619617919
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1619617919
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1619617919
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_144
timestamp 1619617919
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _207_
timestamp 1619617919
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1619617919
transform -1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_160
timestamp 1619617919
transform 1 0 15824 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_172
timestamp 1619617919
transform 1 0 16928 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1619617919
transform 1 0 18860 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1619617919
transform -1 0 17480 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1619617919
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_190
timestamp 1619617919
transform 1 0 18584 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_196
timestamp 1619617919
transform 1 0 19136 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _209_
timestamp 1619617919
transform 1 0 20148 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1619617919
transform -1 0 21804 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1619617919
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_201
timestamp 1619617919
transform 1 0 19596 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_215
timestamp 1619617919
transform 1 0 20884 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_221
timestamp 1619617919
transform 1 0 21436 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1619617919
transform 1 0 1564 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb1
timestamp 1619617919
transform -1 0 3496 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1619617919
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1619617919
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_14
timestamp 1619617919
transform 1 0 2392 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_18
timestamp 1619617919
transform 1 0 2760 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1619617919
transform 1 0 4876 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1619617919
transform 1 0 3956 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen1
timestamp 1619617919
transform 1 0 3496 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_23_34
timestamp 1619617919
transform 1 0 4232 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_40
timestamp 1619617919
transform 1 0 4784 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_44
timestamp 1619617919
transform 1 0 5152 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _246_
timestamp 1619617919
transform 1 0 6808 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _273_
timestamp 1619617919
transform -1 0 6808 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1619617919
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_56
timestamp 1619617919
transform 1 0 6256 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1619617919
transform 1 0 7452 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1619617919
transform 1 0 10212 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _363_
timestamp 1619617919
transform 1 0 9384 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1619617919
transform 1 0 8556 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_89
timestamp 1619617919
transform 1 0 9292 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1619617919
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_102
timestamp 1619617919
transform 1 0 10488 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_115
timestamp 1619617919
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _223_
timestamp 1619617919
transform 1 0 14260 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _224_
timestamp 1619617919
transform 1 0 13064 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_127
timestamp 1619617919
transform 1 0 12788 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1619617919
transform 1 0 13800 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_142
timestamp 1619617919
transform 1 0 14168 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1619617919
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1619617919
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1619617919
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_172
timestamp 1619617919
transform 1 0 16928 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1619617919
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_196
timestamp 1619617919
transform 1 0 19136 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _210_
timestamp 1619617919
transform -1 0 20240 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1619617919
transform -1 0 21804 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_200
timestamp 1619617919
transform 1 0 19504 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1619617919
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_220
timestamp 1619617919
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1619617919
transform 1 0 2024 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1619617919
transform -1 0 3312 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1619617919
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1619617919
transform -1 0 1656 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_6
timestamp 1619617919
transform 1 0 1656 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_17
timestamp 1619617919
transform 1 0 2668 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1619617919
transform 1 0 3312 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1619617919
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_28
timestamp 1619617919
transform 1 0 3680 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1619617919
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_42
timestamp 1619617919
transform 1 0 4968 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_54
timestamp 1619617919
transform 1 0 6072 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_66
timestamp 1619617919
transform 1 0 7176 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _258_
timestamp 1619617919
transform -1 0 8924 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _261_
timestamp 1619617919
transform -1 0 9476 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _395_
timestamp 1619617919
transform 1 0 9936 0 -1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1619617919
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1619617919
transform 1 0 8924 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_91
timestamp 1619617919
transform 1 0 9476 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_95
timestamp 1619617919
transform 1 0 9844 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _222_
timestamp 1619617919
transform -1 0 12880 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_117
timestamp 1619617919
transform 1 0 11868 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _220_
timestamp 1619617919
transform 1 0 14352 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _221_
timestamp 1619617919
transform -1 0 13340 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1619617919
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_133
timestamp 1619617919
transform 1 0 13340 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1619617919
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__and4_1  _284_
timestamp 1619617919
transform 1 0 16928 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_24_152
timestamp 1619617919
transform 1 0 15088 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_164
timestamp 1619617919
transform 1 0 16192 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_179
timestamp 1619617919
transform 1 0 17572 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_191
timestamp 1619617919
transform 1 0 18676 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2ai_1  _228_
timestamp 1619617919
transform -1 0 20240 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1619617919
transform -1 0 21804 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1619617919
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1619617919
transform -1 0 21528 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_199
timestamp 1619617919
transform 1 0 19412 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_208
timestamp 1619617919
transform 1 0 20240 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_216
timestamp 1619617919
transform 1 0 20976 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb0
timestamp 1619617919
transform 1 0 1564 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1619617919
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1619617919
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_12
timestamp 1619617919
transform 1 0 2208 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_24
timestamp 1619617919
transform 1 0 3312 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_36
timestamp 1619617919
transform 1 0 4416 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_48
timestamp 1619617919
transform 1 0 5520 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1619617919
transform 1 0 7176 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _272_
timestamp 1619617919
transform 1 0 6440 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1619617919
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_56
timestamp 1619617919
transform 1 0 6256 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_69
timestamp 1619617919
transform 1 0 7452 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1619617919
transform -1 0 8372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _260_
timestamp 1619617919
transform 1 0 8464 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_75
timestamp 1619617919
transform 1 0 8004 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_79
timestamp 1619617919
transform 1 0 8372 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_88
timestamp 1619617919
transform 1 0 9200 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1619617919
transform -1 0 11224 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1619617919
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_100
timestamp 1619617919
transform 1 0 10304 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_106
timestamp 1619617919
transform 1 0 10856 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_110
timestamp 1619617919
transform 1 0 11224 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1619617919
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__o2bb2a_1  _213_
timestamp 1619617919
transform 1 0 14444 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_127
timestamp 1619617919
transform 1 0 12788 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_139
timestamp 1619617919
transform 1 0 13892 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _206_
timestamp 1619617919
transform 1 0 15732 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _219_
timestamp 1619617919
transform 1 0 15180 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _384_
timestamp 1619617919
transform 1 0 16928 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1619617919
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_162
timestamp 1619617919
transform 1 0 16008 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_170
timestamp 1619617919
transform 1 0 16744 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_1  _227_
timestamp 1619617919
transform 1 0 19044 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_25_192
timestamp 1619617919
transform 1 0 18768 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _208_
timestamp 1619617919
transform 1 0 19596 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1619617919
transform -1 0 21804 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_206
timestamp 1619617919
transform 1 0 20056 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_218
timestamp 1619617919
transform 1 0 21160 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1619617919
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1619617919
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1619617919
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1619617919
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1619617919
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1619617919
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _244_
timestamp 1619617919
transform 1 0 5336 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1619617919
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1619617919
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1619617919
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_42
timestamp 1619617919
transform 1 0 4968 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1619617919
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_39
timestamp 1619617919
transform 1 0 4692 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_45
timestamp 1619617919
transform 1 0 5244 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_56
timestamp 1619617919
transform 1 0 6256 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_55
timestamp 1619617919
transform 1 0 6164 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_50
timestamp 1619617919
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1619617919
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1619617919
transform 1 0 6256 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _270_
timestamp 1619617919
transform 1 0 5796 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _250_
timestamp 1619617919
transform -1 0 7176 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1619617919
transform 1 0 5980 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_71
timestamp 1619617919
transform 1 0 7636 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_66
timestamp 1619617919
transform 1 0 7176 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_59
timestamp 1619617919
transform 1 0 6532 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1619617919
transform 1 0 8924 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_79
timestamp 1619617919
transform 1 0 8372 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_75
timestamp 1619617919
transform 1 0 8004 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1619617919
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1619617919
transform 1 0 8096 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_90
timestamp 1619617919
transform 1 0 9384 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1619617919
transform 1 0 10120 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_78
timestamp 1619617919
transform 1 0 8280 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_99
timestamp 1619617919
transform 1 0 10212 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1619617919
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__a221oi_2  _226_
timestamp 1619617919
transform 1 0 11868 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1619617919
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_111
timestamp 1619617919
transform 1 0 11316 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_123
timestamp 1619617919
transform 1 0 12420 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_101
timestamp 1619617919
transform 1 0 10396 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1619617919
transform 1 0 11500 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_115
timestamp 1619617919
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__or3_1  _237_
timestamp 1619617919
transform 1 0 12972 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _402_
timestamp 1619617919
transform 1 0 14444 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1619617919
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_135
timestamp 1619617919
transform 1 0 13524 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1619617919
transform 1 0 14352 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_134
timestamp 1619617919
transform 1 0 13432 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_142
timestamp 1619617919
transform 1 0 14168 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _289_
timestamp 1619617919
transform 1 0 16836 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1619617919
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_156
timestamp 1619617919
transform 1 0 15456 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_168
timestamp 1619617919
transform 1 0 16560 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_165
timestamp 1619617919
transform 1 0 16284 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1619617919
transform 1 0 16928 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _343_
timestamp 1619617919
transform -1 0 17848 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_182
timestamp 1619617919
transform 1 0 17848 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_194
timestamp 1619617919
transform 1 0 18952 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1619617919
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_196
timestamp 1619617919
transform 1 0 19136 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1619617919
transform -1 0 20516 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _201_
timestamp 1619617919
transform 1 0 19596 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _399_
timestamp 1619617919
transform 1 0 19688 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1619617919
transform -1 0 21804 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1619617919
transform -1 0 21804 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1619617919
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_211
timestamp 1619617919
transform 1 0 20516 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_219
timestamp 1619617919
transform 1 0 21252 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1619617919
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1619617919
transform -1 0 1656 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_6
timestamp 1619617919
transform 1 0 1656 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_18
timestamp 1619617919
transform 1 0 2760 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _274_
timestamp 1619617919
transform -1 0 5796 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _275_
timestamp 1619617919
transform 1 0 4600 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1619617919
transform 1 0 3864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1619617919
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_26
timestamp 1619617919
transform 1 0 3496 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_33
timestamp 1619617919
transform 1 0 4140 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_37
timestamp 1619617919
transform 1 0 4508 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1619617919
transform 1 0 6440 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _256_
timestamp 1619617919
transform 1 0 7820 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _269_
timestamp 1619617919
transform -1 0 6440 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_28_51
timestamp 1619617919
transform 1 0 5796 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_61
timestamp 1619617919
transform 1 0 6716 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _394_
timestamp 1619617919
transform 1 0 9292 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1619617919
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_81
timestamp 1619617919
transform 1 0 8556 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 1619617919
transform 1 0 8924 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_87
timestamp 1619617919
transform 1 0 9108 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1619617919
transform 1 0 12144 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1619617919
transform 1 0 12512 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_110
timestamp 1619617919
transform 1 0 11224 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_118
timestamp 1619617919
transform 1 0 11960 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_123
timestamp 1619617919
transform 1 0 12420 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _198_
timestamp 1619617919
transform -1 0 15180 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1619617919
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_127
timestamp 1619617919
transform 1 0 12788 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_139
timestamp 1619617919
transform 1 0 13892 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_144
timestamp 1619617919
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1619617919
transform 1 0 15180 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1619617919
transform 1 0 16284 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1619617919
transform 1 0 17388 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_189
timestamp 1619617919
transform 1 0 18492 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_197
timestamp 1619617919
transform 1 0 19228 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1619617919
transform -1 0 20976 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1619617919
transform -1 0 21804 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1619617919
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1619617919
transform 1 0 21252 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_201
timestamp 1619617919
transform 1 0 19596 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_216
timestamp 1619617919
transform 1 0 20976 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _391_
timestamp 1619617919
transform 1 0 2668 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1619617919
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1619617919
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_15
timestamp 1619617919
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_38
timestamp 1619617919
transform 1 0 4600 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1619617919
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1619617919
transform 1 0 5704 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_56
timestamp 1619617919
transform 1 0 6256 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_58
timestamp 1619617919
transform 1 0 6440 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_70
timestamp 1619617919
transform 1 0 7544 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _252_
timestamp 1619617919
transform 1 0 8464 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _266_
timestamp 1619617919
transform 1 0 9108 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 1619617919
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_91
timestamp 1619617919
transform 1 0 9476 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_99
timestamp 1619617919
transform 1 0 10212 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _238_
timestamp 1619617919
transform 1 0 12144 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp 1619617919
transform -1 0 10580 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1619617919
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_103
timestamp 1619617919
transform 1 0 10580 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_111
timestamp 1619617919
transform 1 0 11316 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_115
timestamp 1619617919
transform 1 0 11684 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_119
timestamp 1619617919
transform 1 0 12052 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1619617919
transform 1 0 13708 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1619617919
transform 1 0 14812 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1619617919
transform -1 0 16836 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1619617919
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1619617919
transform 1 0 15916 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1619617919
transform 1 0 16468 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_172
timestamp 1619617919
transform 1 0 16928 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1619617919
transform -1 0 18860 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _231_
timestamp 1619617919
transform -1 0 19872 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_29_184
timestamp 1619617919
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_193
timestamp 1619617919
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1619617919
transform -1 0 21804 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_204
timestamp 1619617919
transform 1 0 19872 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_216
timestamp 1619617919
transform 1 0 20976 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1619617919
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1619617919
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1619617919
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1619617919
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1619617919
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_30
timestamp 1619617919
transform 1 0 3864 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_42
timestamp 1619617919
transform 1 0 4968 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1619617919
transform 1 0 6532 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_54
timestamp 1619617919
transform 1 0 6072 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_58
timestamp 1619617919
transform 1 0 6440 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_62
timestamp 1619617919
transform 1 0 6808 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_74
timestamp 1619617919
transform 1 0 7912 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1619617919
transform 1 0 8648 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _265_
timestamp 1619617919
transform 1 0 9108 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1619617919
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1619617919
transform 1 0 8924 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_95
timestamp 1619617919
transform 1 0 9844 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__a41o_2  _234_
timestamp 1619617919
transform 1 0 12236 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_30_107
timestamp 1619617919
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_119
timestamp 1619617919
transform 1 0 12052 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _236_
timestamp 1619617919
transform -1 0 13432 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1619617919
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_134
timestamp 1619617919
transform 1 0 13432 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_142
timestamp 1619617919
transform 1 0 14168 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_144
timestamp 1619617919
transform 1 0 14352 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _283_
timestamp 1619617919
transform 1 0 15824 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _387_
timestamp 1619617919
transform 1 0 16652 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_30_156
timestamp 1619617919
transform 1 0 15456 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _232_
timestamp 1619617919
transform 1 0 18768 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_190
timestamp 1619617919
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_198
timestamp 1619617919
transform 1 0 19320 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _229_
timestamp 1619617919
transform -1 0 19872 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1619617919
transform -1 0 21804 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1619617919
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_204
timestamp 1619617919
transform 1 0 19872 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_216
timestamp 1619617919
transform 1 0 20976 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1619617919
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1619617919
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1619617919
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _240_
timestamp 1619617919
transform 1 0 5152 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1619617919
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_39
timestamp 1619617919
transform 1 0 4692 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_43
timestamp 1619617919
transform 1 0 5060 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _242_
timestamp 1619617919
transform -1 0 6164 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _251_
timestamp 1619617919
transform 1 0 7360 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1619617919
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_55
timestamp 1619617919
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_58
timestamp 1619617919
transform 1 0 6440 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_66
timestamp 1619617919
transform 1 0 7176 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _263_
timestamp 1619617919
transform -1 0 8372 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1619617919
transform 1 0 8556 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_79
timestamp 1619617919
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_84
timestamp 1619617919
transform 1 0 8832 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_96
timestamp 1619617919
transform 1 0 9936 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1619617919
transform -1 0 12788 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1619617919
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_108
timestamp 1619617919
transform 1 0 11040 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_115
timestamp 1619617919
transform 1 0 11684 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_123
timestamp 1619617919
transform 1 0 12420 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _216_
timestamp 1619617919
transform -1 0 14996 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _218_
timestamp 1619617919
transform -1 0 14076 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_127
timestamp 1619617919
transform 1 0 12788 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_135
timestamp 1619617919
transform 1 0 13524 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_141
timestamp 1619617919
transform 1 0 14076 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _214_
timestamp 1619617919
transform 1 0 14996 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1619617919
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_156
timestamp 1619617919
transform 1 0 15456 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_168
timestamp 1619617919
transform 1 0 16560 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_172
timestamp 1619617919
transform 1 0 16928 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp 1619617919
transform -1 0 17848 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_178
timestamp 1619617919
transform 1 0 17480 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_182
timestamp 1619617919
transform 1 0 17848 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_194
timestamp 1619617919
transform 1 0 18952 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp 1619617919
transform -1 0 20700 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1619617919
transform -1 0 21804 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_206
timestamp 1619617919
transform 1 0 20056 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_213
timestamp 1619617919
transform 1 0 20700 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_221
timestamp 1619617919
transform 1 0 21436 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1619617919
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1619617919
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_15
timestamp 1619617919
transform 1 0 2484 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_23
timestamp 1619617919
transform 1 0 3220 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _276_
timestamp 1619617919
transform 1 0 5428 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _277_
timestamp 1619617919
transform 1 0 4692 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1619617919
transform 1 0 3496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1619617919
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_30
timestamp 1619617919
transform 1 0 3864 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_38
timestamp 1619617919
transform 1 0 4600 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1619617919
transform 1 0 5888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _262_
timestamp 1619617919
transform -1 0 8188 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_32_55
timestamp 1619617919
transform 1 0 6164 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_67
timestamp 1619617919
transform 1 0 7268 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_71
timestamp 1619617919
transform 1 0 7636 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _267_
timestamp 1619617919
transform -1 0 8464 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1619617919
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_80
timestamp 1619617919
transform 1 0 8464 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_87
timestamp 1619617919
transform 1 0 9108 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_99
timestamp 1619617919
transform 1 0 10212 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1619617919
transform -1 0 10580 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_103
timestamp 1619617919
transform 1 0 10580 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_115
timestamp 1619617919
transform 1 0 11684 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_1  _215_
timestamp 1619617919
transform -1 0 15088 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1619617919
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_127
timestamp 1619617919
transform 1 0 12788 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_139
timestamp 1619617919
transform 1 0 13892 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1619617919
transform 1 0 15732 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _205_
timestamp 1619617919
transform 1 0 15088 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _282_
timestamp 1619617919
transform -1 0 16468 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_162
timestamp 1619617919
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_167
timestamp 1619617919
transform 1 0 16468 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_179
timestamp 1619617919
transform 1 0 17572 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_191
timestamp 1619617919
transform 1 0 18676 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _383_
timestamp 1619617919
transform 1 0 19596 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1619617919
transform -1 0 21804 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1619617919
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_199
timestamp 1619617919
transform 1 0 19412 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_221
timestamp 1619617919
transform 1 0 21436 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _390_
timestamp 1619617919
transform 1 0 2484 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1619617919
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1619617919
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1619617919
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_6
timestamp 1619617919
transform 1 0 1656 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_14
timestamp 1619617919
transform 1 0 2392 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1619617919
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1619617919
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _241_
timestamp 1619617919
transform 1 0 5244 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1619617919
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_35
timestamp 1619617919
transform 1 0 4324 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_43
timestamp 1619617919
transform 1 0 5060 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_48
timestamp 1619617919
transform 1 0 5520 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1619617919
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_30
timestamp 1619617919
transform 1 0 3864 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_42
timestamp 1619617919
transform 1 0 4968 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_1  _268_
timestamp 1619617919
transform 1 0 7176 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1619617919
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_56
timestamp 1619617919
transform 1 0 6256 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_58
timestamp 1619617919
transform 1 0 6440 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_70
timestamp 1619617919
transform 1 0 7544 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_54
timestamp 1619617919
transform 1 0 6072 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_74
timestamp 1619617919
transform 1 0 7912 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1619617919
transform 1 0 8188 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _398_
timestamp 1619617919
transform 1 0 9568 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1619617919
transform 1 0 9016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_82
timestamp 1619617919
transform 1 0 8648 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_90
timestamp 1619617919
transform 1 0 9384 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_80
timestamp 1619617919
transform 1 0 8464 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_87
timestamp 1619617919
transform 1 0 9108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_99
timestamp 1619617919
transform 1 0 10212 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _202_
timestamp 1619617919
transform -1 0 12420 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _233_
timestamp 1619617919
transform 1 0 11776 0 1 20128
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1619617919
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_112
timestamp 1619617919
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_115
timestamp 1619617919
transform 1 0 11684 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_111
timestamp 1619617919
transform 1 0 11316 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_115
timestamp 1619617919
transform 1 0 11684 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_123
timestamp 1619617919
transform 1 0 12420 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _195_
timestamp 1619617919
transform -1 0 15272 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1619617919
transform 1 0 14260 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_126
timestamp 1619617919
transform 1 0 12696 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_138
timestamp 1619617919
transform 1 0 13800 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_135
timestamp 1619617919
transform 1 0 13524 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_144
timestamp 1619617919
transform 1 0 14352 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1619617919
transform -1 0 15180 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _388_
timestamp 1619617919
transform 1 0 16192 0 -1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1619617919
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_153
timestamp 1619617919
transform 1 0 15180 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_165
timestamp 1619617919
transform 1 0 16284 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_172
timestamp 1619617919
transform 1 0 16928 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_154
timestamp 1619617919
transform 1 0 15272 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_162
timestamp 1619617919
transform 1 0 16008 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1619617919
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_196
timestamp 1619617919
transform 1 0 19136 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_185
timestamp 1619617919
transform 1 0 18124 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_197
timestamp 1619617919
transform 1 0 19228 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _193_
timestamp 1619617919
transform -1 0 21528 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1619617919
transform -1 0 21804 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1619617919
transform -1 0 21804 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1619617919
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output42
timestamp 1619617919
transform 1 0 21160 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_204
timestamp 1619617919
transform 1 0 19872 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_201
timestamp 1619617919
transform 1 0 19596 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_213
timestamp 1619617919
transform 1 0 20700 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_217
timestamp 1619617919
transform 1 0 21068 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _349_
timestamp 1619617919
transform 1 0 1748 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1619617919
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1619617919
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_10
timestamp 1619617919
transform 1 0 2024 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_22
timestamp 1619617919
transform 1 0 3128 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _389_
timestamp 1619617919
transform 1 0 3864 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1619617919
transform 1 0 5704 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _393_
timestamp 1619617919
transform 1 0 6624 0 1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1619617919
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_53
timestamp 1619617919
transform 1 0 5980 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_58
timestamp 1619617919
transform 1 0 6440 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _396_
timestamp 1619617919
transform 1 0 9016 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_35_81
timestamp 1619617919
transform 1 0 8556 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_85
timestamp 1619617919
transform 1 0 8924 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _204_
timestamp 1619617919
transform -1 0 11316 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _397_
timestamp 1619617919
transform 1 0 11776 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1619617919
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_111
timestamp 1619617919
transform 1 0 11316 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_115
timestamp 1619617919
transform 1 0 11684 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _403_
timestamp 1619617919
transform 1 0 14260 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_35_136
timestamp 1619617919
transform 1 0 13616 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_142
timestamp 1619617919
transform 1 0 14168 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1619617919
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_163
timestamp 1619617919
transform 1 0 16100 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_172
timestamp 1619617919
transform 1 0 16928 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _339_
timestamp 1619617919
transform -1 0 17388 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _381_
timestamp 1619617919
transform 1 0 17388 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _382_
timestamp 1619617919
transform 1 0 19228 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1619617919
transform -1 0 21804 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_217
timestamp 1619617919
transform 1 0 21068 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_221
timestamp 1619617919
transform 1 0 21436 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1619617919
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1619617919
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1619617919
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _278_
timestamp 1619617919
transform 1 0 4784 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _338_
timestamp 1619617919
transform 1 0 5428 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1619617919
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1619617919
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_30
timestamp 1619617919
transform 1 0 3864 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_38
timestamp 1619617919
transform 1 0 4600 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1619617919
transform -1 0 7820 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_50
timestamp 1619617919
transform 1 0 5704 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_62
timestamp 1619617919
transform 1 0 6808 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_73
timestamp 1619617919
transform 1 0 7820 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 1619617919
transform -1 0 10120 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1619617919
transform 1 0 9016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_85
timestamp 1619617919
transform 1 0 8924 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_87
timestamp 1619617919
transform 1 0 9108 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_98
timestamp 1619617919
transform 1 0 10120 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _203_
timestamp 1619617919
transform 1 0 11684 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_36_110
timestamp 1619617919
transform 1 0 11224 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_114
timestamp 1619617919
transform 1 0 11592 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_122
timestamp 1619617919
transform 1 0 12328 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1619617919
transform -1 0 12972 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1619617919
transform 1 0 14260 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1619617919
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1619617919
transform 1 0 14076 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_144
timestamp 1619617919
transform 1 0 14352 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp 1619617919
transform -1 0 15456 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_152
timestamp 1619617919
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_156
timestamp 1619617919
transform 1 0 15456 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1619617919
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp 1619617919
transform -1 0 18584 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_180
timestamp 1619617919
transform 1 0 17664 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_186
timestamp 1619617919
transform 1 0 18216 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_190
timestamp 1619617919
transform 1 0 18584 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_198
timestamp 1619617919
transform 1 0 19320 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _345_
timestamp 1619617919
transform -1 0 20240 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1619617919
transform -1 0 21804 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1619617919
transform 1 0 19504 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_201
timestamp 1619617919
transform 1 0 19596 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_208
timestamp 1619617919
transform 1 0 20240 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_220
timestamp 1619617919
transform 1 0 21344 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1619617919
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1619617919
transform 1 0 2760 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1619617919
transform -1 0 2024 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output44
timestamp 1619617919
transform -1 0 1748 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_10
timestamp 1619617919
transform 1 0 2024 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_21
timestamp 1619617919
transform 1 0 3036 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1619617919
transform 1 0 3772 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1619617919
transform 1 0 4600 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_30
timestamp 1619617919
transform 1 0 3864 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_41
timestamp 1619617919
transform 1 0 4876 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1619617919
transform 1 0 6440 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1619617919
transform 1 0 7820 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1619617919
transform 1 0 5980 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_56
timestamp 1619617919
transform 1 0 6256 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_59
timestamp 1619617919
transform 1 0 6532 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_71
timestamp 1619617919
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1619617919
transform 1 0 9108 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1619617919
transform 1 0 9660 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_76
timestamp 1619617919
transform 1 0 8096 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_84
timestamp 1619617919
transform 1 0 8832 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_88
timestamp 1619617919
transform 1 0 9200 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_92
timestamp 1619617919
transform 1 0 9568 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_96
timestamp 1619617919
transform 1 0 9936 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1619617919
transform 1 0 11776 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1619617919
transform 1 0 11500 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1619617919
transform 1 0 11040 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_112
timestamp 1619617919
transform 1 0 11408 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_117
timestamp 1619617919
transform 1 0 11868 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1619617919
transform 1 0 14444 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1619617919
transform -1 0 14996 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1619617919
transform 1 0 12880 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_125
timestamp 1619617919
transform 1 0 12604 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_131
timestamp 1619617919
transform 1 0 13156 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_143
timestamp 1619617919
transform 1 0 14260 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_146
timestamp 1619617919
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1619617919
transform -1 0 16836 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_151
timestamp 1619617919
transform 1 0 14996 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_163
timestamp 1619617919
transform 1 0 16100 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1619617919
transform 1 0 16468 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_171
timestamp 1619617919
transform 1 0 16836 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1619617919
transform 1 0 17112 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1619617919
transform 1 0 17940 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_175
timestamp 1619617919
transform 1 0 17204 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_186
timestamp 1619617919
transform 1 0 18216 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_198
timestamp 1619617919
transform 1 0 19320 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1619617919
transform -1 0 21804 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1619617919
transform 1 0 19780 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1619617919
transform -1 0 20148 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1619617919
transform -1 0 21160 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 21528 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_202
timestamp 1619617919
transform 1 0 19688 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_207
timestamp 1619617919
transform 1 0 20148 0 1 22304
box -38 -48 774 592
<< labels >>
rlabel metal3 s 0 10208 800 10328 6 clockc
port 0 nsew signal tristate
rlabel metal3 s 0 12928 800 13048 6 clockd[0]
port 1 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 clockd[1]
port 2 nsew signal tristate
rlabel metal3 s 22179 20408 22979 20528 6 clockd[2]
port 3 nsew signal tristate
rlabel metal2 s 20718 0 20774 800 6 clockd[3]
port 4 nsew signal tristate
rlabel metal3 s 0 23128 800 23248 6 clockp[0]
port 5 nsew signal tristate
rlabel metal2 s 1858 0 1914 800 6 clockp[1]
port 6 nsew signal tristate
rlabel metal2 s 15658 0 15714 800 6 dco
port 7 nsew signal input
rlabel metal3 s 22179 15648 22979 15768 6 div[0]
port 8 nsew signal input
rlabel metal2 s 19798 24323 19854 25123 6 div[1]
port 9 nsew signal input
rlabel metal2 s 7838 24323 7894 25123 6 div[2]
port 10 nsew signal input
rlabel metal2 s 478 0 534 800 6 div[3]
port 11 nsew signal input
rlabel metal2 s 14738 24323 14794 25123 6 div[4]
port 12 nsew signal input
rlabel metal2 s 16578 24323 16634 25123 6 ext_trim[0]
port 13 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 ext_trim[10]
port 14 nsew signal input
rlabel metal2 s 2778 24323 2834 25123 6 ext_trim[11]
port 15 nsew signal input
rlabel metal3 s 22179 5448 22979 5568 6 ext_trim[12]
port 16 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 ext_trim[13]
port 17 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 ext_trim[14]
port 18 nsew signal input
rlabel metal3 s 22179 17688 22979 17808 6 ext_trim[15]
port 19 nsew signal input
rlabel metal2 s 4618 24323 4674 25123 6 ext_trim[16]
port 20 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 ext_trim[17]
port 21 nsew signal input
rlabel metal2 s 5998 24323 6054 25123 6 ext_trim[18]
port 22 nsew signal input
rlabel metal3 s 22179 10208 22979 10328 6 ext_trim[19]
port 23 nsew signal input
rlabel metal2 s 12898 24323 12954 25123 6 ext_trim[1]
port 24 nsew signal input
rlabel metal2 s 11518 24323 11574 25123 6 ext_trim[20]
port 25 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 ext_trim[21]
port 26 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 ext_trim[22]
port 27 nsew signal input
rlabel metal3 s 22179 23128 22979 23248 6 ext_trim[23]
port 28 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 ext_trim[24]
port 29 nsew signal input
rlabel metal2 s 9678 24323 9734 25123 6 ext_trim[25]
port 30 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 ext_trim[2]
port 31 nsew signal input
rlabel metal3 s 22179 8168 22979 8288 6 ext_trim[3]
port 32 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 ext_trim[4]
port 33 nsew signal input
rlabel metal3 s 22179 12928 22979 13048 6 ext_trim[5]
port 34 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 ext_trim[6]
port 35 nsew signal input
rlabel metal2 s 938 24323 994 25123 6 ext_trim[7]
port 36 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 ext_trim[8]
port 37 nsew signal input
rlabel metal3 s 22179 2728 22979 2848 6 ext_trim[9]
port 38 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 extclk_sel
port 39 nsew signal input
rlabel metal2 s 17958 24323 18014 25123 6 osc
port 40 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 reset
port 41 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 sel[0]
port 42 nsew signal input
rlabel metal2 s 21638 24323 21694 25123 6 sel[1]
port 43 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 sel[2]
port 44 nsew signal input
rlabel metal4 s 18194 2128 18514 22896 6 VPWR
port 45 nsew power bidirectional
rlabel metal4 s 11294 2128 11614 22896 6 VPWR
port 46 nsew power bidirectional
rlabel metal4 s 4394 2128 4714 22896 6 VPWR
port 47 nsew power bidirectional
rlabel metal5 s 1104 19195 21804 19515 6 VPWR
port 48 nsew power bidirectional
rlabel metal5 s 1104 12304 21804 12624 6 VPWR
port 49 nsew power bidirectional
rlabel metal5 s 1104 5413 21804 5733 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 14744 2128 15064 22896 6 VGND
port 51 nsew ground bidirectional
rlabel metal4 s 7844 2128 8164 22896 6 VGND
port 52 nsew ground bidirectional
rlabel metal5 s 1104 15749 21804 16069 6 VGND
port 53 nsew ground bidirectional
rlabel metal5 s 1104 8859 21804 9179 6 VGND
port 54 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 22979 25123
<< end >>
