magic
tech sky130A
magscale 1 2
timestamp 1619613117
<< locali >>
rect 7113 20791 7147 20893
rect 8953 11135 8987 11305
rect 9413 8483 9447 8585
<< viali >>
rect 1501 22729 1535 22763
rect 2973 22661 3007 22695
rect 8033 22661 8067 22695
rect 2329 22525 2363 22559
rect 2789 22525 2823 22559
rect 4721 22525 4755 22559
rect 5365 22525 5399 22559
rect 7113 22525 7147 22559
rect 7849 22525 7883 22559
rect 9689 22525 9723 22559
rect 12449 22525 12483 22559
rect 12909 22525 12943 22559
rect 15117 22525 15151 22559
rect 16681 22525 16715 22559
rect 18153 22525 18187 22559
rect 19349 22525 19383 22559
rect 21097 22525 21131 22559
rect 1593 22457 1627 22491
rect 2145 22389 2179 22423
rect 4905 22389 4939 22423
rect 5549 22389 5583 22423
rect 6929 22389 6963 22423
rect 9873 22389 9907 22423
rect 12265 22389 12299 22423
rect 13093 22389 13127 22423
rect 14933 22389 14967 22423
rect 16497 22389 16531 22423
rect 17969 22389 18003 22423
rect 19165 22389 19199 22423
rect 20913 22389 20947 22423
rect 10885 22117 10919 22151
rect 11897 22117 11931 22151
rect 4997 22049 5031 22083
rect 5089 22049 5123 22083
rect 5365 22049 5399 22083
rect 7573 22049 7607 22083
rect 9873 22049 9907 22083
rect 11069 22049 11103 22083
rect 11713 22049 11747 22083
rect 11989 22049 12023 22083
rect 12127 22049 12161 22083
rect 12909 22049 12943 22083
rect 15393 22049 15427 22083
rect 18337 22049 18371 22083
rect 19993 22049 20027 22083
rect 21097 22049 21131 22083
rect 20913 21913 20947 21947
rect 4813 21845 4847 21879
rect 5273 21845 5307 21879
rect 7757 21845 7791 21879
rect 10057 21845 10091 21879
rect 10701 21845 10735 21879
rect 12265 21845 12299 21879
rect 12725 21845 12759 21879
rect 15209 21845 15243 21879
rect 18521 21845 18555 21879
rect 20177 21845 20211 21879
rect 1777 21641 1811 21675
rect 10885 21641 10919 21675
rect 8585 21573 8619 21607
rect 4169 21505 4203 21539
rect 9137 21505 9171 21539
rect 9413 21505 9447 21539
rect 13553 21505 13587 21539
rect 16037 21505 16071 21539
rect 17417 21505 17451 21539
rect 21005 21505 21039 21539
rect 1961 21437 1995 21471
rect 3893 21437 3927 21471
rect 6837 21437 6871 21471
rect 13829 21437 13863 21471
rect 20177 21437 20211 21471
rect 20361 21437 20395 21471
rect 20913 21437 20947 21471
rect 7113 21369 7147 21403
rect 15761 21369 15795 21403
rect 17693 21369 17727 21403
rect 19809 21369 19843 21403
rect 5641 21301 5675 21335
rect 12081 21301 12115 21335
rect 14289 21301 14323 21335
rect 19165 21301 19199 21335
rect 5273 21097 5307 21131
rect 7205 21097 7239 21131
rect 15301 21097 15335 21131
rect 7481 21029 7515 21063
rect 7711 21029 7745 21063
rect 12081 21029 12115 21063
rect 15025 21029 15059 21063
rect 5365 20961 5399 20995
rect 7389 20961 7423 20995
rect 7573 20961 7607 20995
rect 8309 20961 8343 20995
rect 11989 20961 12023 20995
rect 12173 20961 12207 20995
rect 12357 20961 12391 20995
rect 14749 20961 14783 20995
rect 14933 20961 14967 20995
rect 15117 20961 15151 20995
rect 16221 20961 16255 20995
rect 20913 20961 20947 20995
rect 7113 20893 7147 20927
rect 7849 20893 7883 20927
rect 16497 20893 16531 20927
rect 7113 20757 7147 20791
rect 8401 20757 8435 20791
rect 11805 20757 11839 20791
rect 17969 20757 18003 20791
rect 21005 20757 21039 20791
rect 7757 20553 7791 20587
rect 17325 20553 17359 20587
rect 11161 20485 11195 20519
rect 12541 20485 12575 20519
rect 2513 20417 2547 20451
rect 9413 20417 9447 20451
rect 9689 20417 9723 20451
rect 14197 20417 14231 20451
rect 15853 20417 15887 20451
rect 19349 20417 19383 20451
rect 1409 20349 1443 20383
rect 5273 20349 5307 20383
rect 5457 20349 5491 20383
rect 7665 20349 7699 20383
rect 7849 20349 7883 20383
rect 12081 20349 12115 20383
rect 12265 20349 12299 20383
rect 12633 20349 12667 20383
rect 12909 20349 12943 20383
rect 14289 20349 14323 20383
rect 14749 20349 14783 20383
rect 15117 20349 15151 20383
rect 15945 20349 15979 20383
rect 17509 20349 17543 20383
rect 19073 20349 19107 20383
rect 2789 20281 2823 20315
rect 14933 20281 14967 20315
rect 15025 20281 15059 20315
rect 1593 20213 1627 20247
rect 4261 20213 4295 20247
rect 5365 20213 5399 20247
rect 15301 20213 15335 20247
rect 20821 20213 20855 20247
rect 3341 20009 3375 20043
rect 4721 20009 4755 20043
rect 6193 20009 6227 20043
rect 8125 20009 8159 20043
rect 10517 20009 10551 20043
rect 16221 20009 16255 20043
rect 4997 19941 5031 19975
rect 6009 19941 6043 19975
rect 16405 19941 16439 19975
rect 3157 19873 3191 19907
rect 4905 19873 4939 19907
rect 5089 19873 5123 19907
rect 5207 19873 5241 19907
rect 5825 19873 5859 19907
rect 7757 19873 7791 19907
rect 7941 19873 7975 19907
rect 10333 19873 10367 19907
rect 14933 19873 14967 19907
rect 16129 19873 16163 19907
rect 20637 19873 20671 19907
rect 5365 19805 5399 19839
rect 15025 19805 15059 19839
rect 15393 19805 15427 19839
rect 16405 19737 16439 19771
rect 14749 19669 14783 19703
rect 20453 19669 20487 19703
rect 5181 19465 5215 19499
rect 15761 19465 15795 19499
rect 21097 19465 21131 19499
rect 5641 19329 5675 19363
rect 14657 19329 14691 19363
rect 19625 19329 19659 19363
rect 4537 19261 4571 19295
rect 5365 19261 5399 19295
rect 5457 19261 5491 19295
rect 5733 19261 5767 19295
rect 7389 19261 7423 19295
rect 7757 19261 7791 19295
rect 8493 19261 8527 19295
rect 8586 19261 8620 19295
rect 8958 19261 8992 19295
rect 9597 19261 9631 19295
rect 12725 19261 12759 19295
rect 13553 19261 13587 19295
rect 13737 19261 13771 19295
rect 14398 19261 14432 19295
rect 14565 19261 14599 19295
rect 14749 19261 14783 19295
rect 14933 19261 14967 19295
rect 15577 19261 15611 19295
rect 17601 19261 17635 19295
rect 19349 19261 19383 19295
rect 4629 19193 4663 19227
rect 7573 19193 7607 19227
rect 7665 19193 7699 19227
rect 8769 19193 8803 19227
rect 8861 19193 8895 19227
rect 9689 19193 9723 19227
rect 14197 19193 14231 19227
rect 15393 19193 15427 19227
rect 7941 19125 7975 19159
rect 9137 19125 9171 19159
rect 12633 19125 12667 19159
rect 13553 19125 13587 19159
rect 17785 19125 17819 19159
rect 6653 18921 6687 18955
rect 9597 18921 9631 18955
rect 20269 18921 20303 18955
rect 8125 18853 8159 18887
rect 13001 18853 13035 18887
rect 16221 18853 16255 18887
rect 16957 18853 16991 18887
rect 5641 18785 5675 18819
rect 6561 18785 6595 18819
rect 7849 18785 7883 18819
rect 9505 18785 9539 18819
rect 12541 18785 12575 18819
rect 12633 18785 12667 18819
rect 12909 18785 12943 18819
rect 13737 18785 13771 18819
rect 15485 18785 15519 18819
rect 15669 18785 15703 18819
rect 16037 18785 16071 18819
rect 16681 18785 16715 18819
rect 20361 18785 20395 18819
rect 20453 18785 20487 18819
rect 20913 18785 20947 18819
rect 21097 18785 21131 18819
rect 5365 18717 5399 18751
rect 5549 18717 5583 18751
rect 8125 18717 8159 18751
rect 12817 18717 12851 18751
rect 13461 18717 13495 18751
rect 15761 18717 15795 18751
rect 15853 18717 15887 18751
rect 18429 18717 18463 18751
rect 19993 18717 20027 18751
rect 5457 18649 5491 18683
rect 12357 18649 12391 18683
rect 7941 18581 7975 18615
rect 13553 18581 13587 18615
rect 13645 18581 13679 18615
rect 21005 18581 21039 18615
rect 8953 18377 8987 18411
rect 17417 18377 17451 18411
rect 19073 18377 19107 18411
rect 18521 18309 18555 18343
rect 4537 18241 4571 18275
rect 9505 18241 9539 18275
rect 12173 18241 12207 18275
rect 19441 18241 19475 18275
rect 19533 18241 19567 18275
rect 5457 18173 5491 18207
rect 8677 18173 8711 18207
rect 8769 18173 8803 18207
rect 9045 18173 9079 18207
rect 9689 18173 9723 18207
rect 9781 18173 9815 18207
rect 10333 18173 10367 18207
rect 12633 18173 12667 18207
rect 12817 18173 12851 18207
rect 13001 18173 13035 18207
rect 13185 18173 13219 18207
rect 13553 18173 13587 18207
rect 17325 18173 17359 18207
rect 17509 18173 17543 18207
rect 18613 18173 18647 18207
rect 19257 18173 19291 18207
rect 19625 18173 19659 18207
rect 19809 18173 19843 18207
rect 21097 18173 21131 18207
rect 4261 18105 4295 18139
rect 5641 18105 5675 18139
rect 2789 18037 2823 18071
rect 5273 18037 5307 18071
rect 8493 18037 8527 18071
rect 9505 18037 9539 18071
rect 10517 18037 10551 18071
rect 20913 18037 20947 18071
rect 3341 17833 3375 17867
rect 4629 17833 4663 17867
rect 12633 17833 12667 17867
rect 4905 17765 4939 17799
rect 6009 17765 6043 17799
rect 6193 17765 6227 17799
rect 6929 17765 6963 17799
rect 9781 17765 9815 17799
rect 14933 17765 14967 17799
rect 15025 17765 15059 17799
rect 1409 17697 1443 17731
rect 3157 17697 3191 17731
rect 4813 17697 4847 17731
rect 4997 17697 5031 17731
rect 5115 17697 5149 17731
rect 6377 17697 6411 17731
rect 6837 17697 6871 17731
rect 8033 17697 8067 17731
rect 8493 17697 8527 17731
rect 9505 17697 9539 17731
rect 12265 17697 12299 17731
rect 13093 17697 13127 17731
rect 14749 17697 14783 17731
rect 15117 17697 15151 17731
rect 20913 17697 20947 17731
rect 5273 17629 5307 17663
rect 8217 17629 8251 17663
rect 8309 17629 8343 17663
rect 12357 17629 12391 17663
rect 8125 17561 8159 17595
rect 13185 17561 13219 17595
rect 1593 17493 1627 17527
rect 7849 17493 7883 17527
rect 11253 17493 11287 17527
rect 12449 17493 12483 17527
rect 15301 17493 15335 17527
rect 20729 17493 20763 17527
rect 7481 17289 7515 17323
rect 10241 17289 10275 17323
rect 14473 17289 14507 17323
rect 12173 17221 12207 17255
rect 5825 17153 5859 17187
rect 7113 17153 7147 17187
rect 12633 17153 12667 17187
rect 12817 17153 12851 17187
rect 15945 17153 15979 17187
rect 16221 17153 16255 17187
rect 19349 17153 19383 17187
rect 5549 17085 5583 17119
rect 5641 17085 5675 17119
rect 5917 17085 5951 17119
rect 6837 17085 6871 17119
rect 7021 17085 7055 17119
rect 7205 17085 7239 17119
rect 7297 17085 7331 17119
rect 8309 17085 8343 17119
rect 10149 17085 10183 17119
rect 12081 17085 12115 17119
rect 12541 17085 12575 17119
rect 12909 17085 12943 17119
rect 19625 17017 19659 17051
rect 5365 16949 5399 16983
rect 8217 16949 8251 16983
rect 21097 16949 21131 16983
rect 6653 16745 6687 16779
rect 12265 16745 12299 16779
rect 20545 16745 20579 16779
rect 6101 16677 6135 16711
rect 17233 16677 17267 16711
rect 18981 16677 19015 16711
rect 20269 16677 20303 16711
rect 5825 16609 5859 16643
rect 5917 16609 5951 16643
rect 6561 16609 6595 16643
rect 8125 16609 8159 16643
rect 8217 16609 8251 16643
rect 12173 16609 12207 16643
rect 14933 16609 14967 16643
rect 15117 16609 15151 16643
rect 15209 16609 15243 16643
rect 16865 16609 16899 16643
rect 16957 16609 16991 16643
rect 17141 16609 17175 16643
rect 17325 16609 17359 16643
rect 17969 16609 18003 16643
rect 19073 16609 19107 16643
rect 19993 16609 20027 16643
rect 20177 16609 20211 16643
rect 20361 16609 20395 16643
rect 6101 16541 6135 16575
rect 14749 16405 14783 16439
rect 17509 16405 17543 16439
rect 18153 16405 18187 16439
rect 9781 16201 9815 16235
rect 12173 16201 12207 16235
rect 15577 16201 15611 16235
rect 19993 16201 20027 16235
rect 9137 16133 9171 16167
rect 15117 16133 15151 16167
rect 19073 16133 19107 16167
rect 9597 16065 9631 16099
rect 12817 16065 12851 16099
rect 14473 16065 14507 16099
rect 17325 16065 17359 16099
rect 17601 16065 17635 16099
rect 1593 15997 1627 16031
rect 2145 15997 2179 16031
rect 5917 15997 5951 16031
rect 6975 15997 7009 16031
rect 7205 15997 7239 16031
rect 7333 15997 7367 16031
rect 7481 15997 7515 16031
rect 8493 15997 8527 16031
rect 8586 15997 8620 16031
rect 8861 15997 8895 16031
rect 8958 15997 8992 16031
rect 9873 15997 9907 16031
rect 10977 15997 11011 16031
rect 12357 15997 12391 16031
rect 12449 15997 12483 16031
rect 14565 15997 14599 16031
rect 14936 15997 14970 16031
rect 15577 15997 15611 16031
rect 15761 15997 15795 16031
rect 19533 15997 19567 16031
rect 19809 15997 19843 16031
rect 20453 15997 20487 16031
rect 20637 15997 20671 16031
rect 2053 15929 2087 15963
rect 5825 15929 5859 15963
rect 7113 15929 7147 15963
rect 8769 15929 8803 15963
rect 6837 15861 6871 15895
rect 9597 15861 9631 15895
rect 11161 15861 11195 15895
rect 14933 15861 14967 15895
rect 19625 15861 19659 15895
rect 20545 15861 20579 15895
rect 7113 15657 7147 15691
rect 8585 15657 8619 15691
rect 13185 15657 13219 15691
rect 13369 15657 13403 15691
rect 17141 15657 17175 15691
rect 17233 15657 17267 15691
rect 20269 15657 20303 15691
rect 10241 15589 10275 15623
rect 12357 15589 12391 15623
rect 12725 15589 12759 15623
rect 1409 15521 1443 15555
rect 2605 15521 2639 15555
rect 3065 15521 3099 15555
rect 3249 15521 3283 15555
rect 4445 15521 4479 15555
rect 6561 15521 6595 15555
rect 7021 15521 7055 15555
rect 8033 15521 8067 15555
rect 8309 15521 8343 15555
rect 8401 15521 8435 15555
rect 12541 15521 12575 15555
rect 13366 15521 13400 15555
rect 13737 15521 13771 15555
rect 16957 15521 16991 15555
rect 17325 15521 17359 15555
rect 19993 15521 20027 15555
rect 20177 15521 20211 15555
rect 20453 15521 20487 15555
rect 20545 15521 20579 15555
rect 2053 15453 2087 15487
rect 6285 15453 6319 15487
rect 8125 15453 8159 15487
rect 9965 15453 9999 15487
rect 13829 15453 13863 15487
rect 2513 15385 2547 15419
rect 6469 15385 6503 15419
rect 1593 15317 1627 15351
rect 4261 15317 4295 15351
rect 6377 15317 6411 15351
rect 11713 15317 11747 15351
rect 17509 15317 17543 15351
rect 1593 15113 1627 15147
rect 6837 15113 6871 15147
rect 7297 15113 7331 15147
rect 10701 15113 10735 15147
rect 13093 15113 13127 15147
rect 18981 15113 19015 15147
rect 20913 15113 20947 15147
rect 4261 15045 4295 15079
rect 9505 15045 9539 15079
rect 14289 15045 14323 15079
rect 2053 14977 2087 15011
rect 2145 14977 2179 15011
rect 3893 14977 3927 15011
rect 9965 14977 9999 15011
rect 13645 14977 13679 15011
rect 13737 14977 13771 15011
rect 2881 14909 2915 14943
rect 3433 14909 3467 14943
rect 5089 14909 5123 14943
rect 7021 14909 7055 14943
rect 7113 14909 7147 14943
rect 7389 14909 7423 14943
rect 10609 14909 10643 14943
rect 13277 14909 13311 14943
rect 13369 14909 13403 14943
rect 14565 14909 14599 14943
rect 15025 14909 15059 14943
rect 15209 14909 15243 14943
rect 18889 14909 18923 14943
rect 19809 14909 19843 14943
rect 19993 14909 20027 14943
rect 20177 14909 20211 14943
rect 21097 14909 21131 14943
rect 2973 14841 3007 14875
rect 10057 14841 10091 14875
rect 14289 14841 14323 14875
rect 15117 14841 15151 14875
rect 19901 14841 19935 14875
rect 1961 14773 1995 14807
rect 4261 14773 4295 14807
rect 4905 14773 4939 14807
rect 9965 14773 9999 14807
rect 14473 14773 14507 14807
rect 19625 14773 19659 14807
rect 14749 14569 14783 14603
rect 14933 14569 14967 14603
rect 18061 14569 18095 14603
rect 20177 14569 20211 14603
rect 20361 14569 20395 14603
rect 5825 14501 5859 14535
rect 12909 14501 12943 14535
rect 6561 14433 6595 14467
rect 7389 14433 7423 14467
rect 12817 14433 12851 14467
rect 14930 14433 14964 14467
rect 15393 14433 15427 14467
rect 16037 14433 16071 14467
rect 17325 14433 17359 14467
rect 18153 14433 18187 14467
rect 18981 14433 19015 14467
rect 20358 14433 20392 14467
rect 20821 14433 20855 14467
rect 4353 14365 4387 14399
rect 6101 14365 6135 14399
rect 6653 14229 6687 14263
rect 7481 14229 7515 14263
rect 15301 14229 15335 14263
rect 15945 14229 15979 14263
rect 17417 14229 17451 14263
rect 18889 14229 18923 14263
rect 20729 14229 20763 14263
rect 6837 14025 6871 14059
rect 8769 14025 8803 14059
rect 9689 14025 9723 14059
rect 10241 14025 10275 14059
rect 20913 14025 20947 14059
rect 3157 13957 3191 13991
rect 7297 13889 7331 13923
rect 17601 13889 17635 13923
rect 18981 13889 19015 13923
rect 7021 13821 7055 13855
rect 7113 13821 7147 13855
rect 7205 13821 7239 13855
rect 8033 13821 8067 13855
rect 8217 13821 8251 13855
rect 8677 13821 8711 13855
rect 9505 13821 9539 13855
rect 9781 13821 9815 13855
rect 9873 13821 9907 13855
rect 9965 13821 9999 13855
rect 12173 13821 12207 13855
rect 12265 13821 12299 13855
rect 14289 13821 14323 13855
rect 14381 13821 14415 13855
rect 14657 13821 14691 13855
rect 17509 13821 17543 13855
rect 17693 13821 17727 13855
rect 17785 13821 17819 13855
rect 18705 13821 18739 13855
rect 18889 13821 18923 13855
rect 19073 13821 19107 13855
rect 19257 13821 19291 13855
rect 21097 13821 21131 13855
rect 3341 13753 3375 13787
rect 7849 13753 7883 13787
rect 14473 13753 14507 13787
rect 12449 13685 12483 13719
rect 14105 13685 14139 13719
rect 17325 13685 17359 13719
rect 18521 13685 18555 13719
rect 1869 13481 1903 13515
rect 7389 13481 7423 13515
rect 8309 13481 8343 13515
rect 18153 13481 18187 13515
rect 6101 13413 6135 13447
rect 6469 13413 6503 13447
rect 11253 13413 11287 13447
rect 12081 13413 12115 13447
rect 12173 13413 12207 13447
rect 12357 13413 12391 13447
rect 15669 13413 15703 13447
rect 17417 13413 17451 13447
rect 1961 13345 1995 13379
rect 6285 13345 6319 13379
rect 7297 13345 7331 13379
rect 8217 13345 8251 13379
rect 9505 13345 9539 13379
rect 9689 13345 9723 13379
rect 11069 13345 11103 13379
rect 18337 13345 18371 13379
rect 18521 13345 18555 13379
rect 20131 13345 20165 13379
rect 20269 13345 20303 13379
rect 20361 13345 20395 13379
rect 20545 13345 20579 13379
rect 1777 13277 1811 13311
rect 17693 13277 17727 13311
rect 2329 13141 2363 13175
rect 9505 13141 9539 13175
rect 9873 13141 9907 13175
rect 11437 13141 11471 13175
rect 12633 13141 12667 13175
rect 18521 13141 18555 13175
rect 19993 13141 20027 13175
rect 1501 12937 1535 12971
rect 2697 12937 2731 12971
rect 3525 12937 3559 12971
rect 4905 12937 4939 12971
rect 5273 12937 5307 12971
rect 9965 12937 9999 12971
rect 10057 12937 10091 12971
rect 10977 12937 11011 12971
rect 15577 12937 15611 12971
rect 16405 12937 16439 12971
rect 17417 12937 17451 12971
rect 21097 12937 21131 12971
rect 3157 12801 3191 12835
rect 13185 12801 13219 12835
rect 13829 12801 13863 12835
rect 14105 12801 14139 12835
rect 17325 12801 17359 12835
rect 17509 12801 17543 12835
rect 19349 12801 19383 12835
rect 19625 12801 19659 12835
rect 2145 12733 2179 12767
rect 2697 12733 2731 12767
rect 3525 12733 3559 12767
rect 5181 12733 5215 12767
rect 5273 12733 5307 12767
rect 7757 12733 7791 12767
rect 8677 12733 8711 12767
rect 8953 12733 8987 12767
rect 9689 12733 9723 12767
rect 9873 12733 9907 12767
rect 10149 12733 10183 12767
rect 10885 12733 10919 12767
rect 11069 12733 11103 12767
rect 13093 12733 13127 12767
rect 16221 12733 16255 12767
rect 17601 12733 17635 12767
rect 18521 12733 18555 12767
rect 1593 12665 1627 12699
rect 7573 12665 7607 12699
rect 10425 12665 10459 12699
rect 18705 12665 18739 12699
rect 7849 12597 7883 12631
rect 8861 12597 8895 12631
rect 12633 12597 12667 12631
rect 13001 12597 13035 12631
rect 18889 12597 18923 12631
rect 5549 12393 5583 12427
rect 11897 12393 11931 12427
rect 12265 12393 12299 12427
rect 13093 12393 13127 12427
rect 14933 12393 14967 12427
rect 20637 12393 20671 12427
rect 3341 12325 3375 12359
rect 11805 12325 11839 12359
rect 12725 12325 12759 12359
rect 3157 12257 3191 12291
rect 5641 12257 5675 12291
rect 6377 12257 6411 12291
rect 7573 12257 7607 12291
rect 12909 12257 12943 12291
rect 14749 12257 14783 12291
rect 20821 12257 20855 12291
rect 5549 12189 5583 12223
rect 6469 12189 6503 12223
rect 6561 12189 6595 12223
rect 6653 12189 6687 12223
rect 7849 12189 7883 12223
rect 11621 12189 11655 12223
rect 6193 12121 6227 12155
rect 7757 12121 7791 12155
rect 5089 12053 5123 12087
rect 7665 12053 7699 12087
rect 2973 11849 3007 11883
rect 8401 11849 8435 11883
rect 9413 11781 9447 11815
rect 5549 11713 5583 11747
rect 5733 11713 5767 11747
rect 6837 11713 6871 11747
rect 7941 11713 7975 11747
rect 8217 11713 8251 11747
rect 10517 11713 10551 11747
rect 2973 11645 3007 11679
rect 3525 11645 3559 11679
rect 5641 11645 5675 11679
rect 5825 11645 5859 11679
rect 7021 11645 7055 11679
rect 7205 11645 7239 11679
rect 8033 11645 8067 11679
rect 8125 11645 8159 11679
rect 9321 11645 9355 11679
rect 9597 11645 9631 11679
rect 10609 11645 10643 11679
rect 10793 11645 10827 11679
rect 5365 11509 5399 11543
rect 9781 11509 9815 11543
rect 10977 11509 11011 11543
rect 2053 11305 2087 11339
rect 2973 11305 3007 11339
rect 8953 11305 8987 11339
rect 10262 11305 10296 11339
rect 12909 11305 12943 11339
rect 18521 11305 18555 11339
rect 7021 11237 7055 11271
rect 1961 11169 1995 11203
rect 4445 11169 4479 11203
rect 6182 11169 6216 11203
rect 6285 11169 6319 11203
rect 6929 11169 6963 11203
rect 7573 11169 7607 11203
rect 7757 11169 7791 11203
rect 8125 11169 8159 11203
rect 10057 11237 10091 11271
rect 11621 11237 11655 11271
rect 11805 11237 11839 11271
rect 13001 11169 13035 11203
rect 15025 11169 15059 11203
rect 16957 11169 16991 11203
rect 17417 11169 17451 11203
rect 18429 11169 18463 11203
rect 20085 11169 20119 11203
rect 2237 11101 2271 11135
rect 2973 11101 3007 11135
rect 3341 11101 3375 11135
rect 6101 11101 6135 11135
rect 6377 11101 6411 11135
rect 8953 11101 8987 11135
rect 11897 11101 11931 11135
rect 12725 11101 12759 11135
rect 18613 11101 18647 11135
rect 4261 11033 4295 11067
rect 7757 11033 7791 11067
rect 10425 11033 10459 11067
rect 11345 11033 11379 11067
rect 13369 11033 13403 11067
rect 15209 11033 15243 11067
rect 17601 11033 17635 11067
rect 18061 11033 18095 11067
rect 20269 11033 20303 11067
rect 1593 10965 1627 10999
rect 5917 10965 5951 10999
rect 10241 10965 10275 10999
rect 16865 10965 16899 10999
rect 4629 10761 4663 10795
rect 4997 10761 5031 10795
rect 7573 10761 7607 10795
rect 13461 10761 13495 10795
rect 20913 10761 20947 10795
rect 16221 10693 16255 10727
rect 5089 10625 5123 10659
rect 7389 10625 7423 10659
rect 13093 10625 13127 10659
rect 15853 10625 15887 10659
rect 18337 10625 18371 10659
rect 19441 10625 19475 10659
rect 2697 10557 2731 10591
rect 4813 10557 4847 10591
rect 7665 10557 7699 10591
rect 9045 10557 9079 10591
rect 9597 10557 9631 10591
rect 13461 10557 13495 10591
rect 14841 10557 14875 10591
rect 15393 10557 15427 10591
rect 18061 10557 18095 10591
rect 19165 10557 19199 10591
rect 1593 10489 1627 10523
rect 2881 10489 2915 10523
rect 8493 10489 8527 10523
rect 15301 10489 15335 10523
rect 1501 10421 1535 10455
rect 7389 10421 7423 10455
rect 9689 10421 9723 10455
rect 16221 10421 16255 10455
rect 17693 10421 17727 10455
rect 18153 10421 18187 10455
rect 2237 10217 2271 10251
rect 5273 10217 5307 10251
rect 6745 10217 6779 10251
rect 7573 10217 7607 10251
rect 11897 10217 11931 10251
rect 18245 10217 18279 10251
rect 20913 10217 20947 10251
rect 5457 10149 5491 10183
rect 6653 10149 6687 10183
rect 13369 10149 13403 10183
rect 17325 10149 17359 10183
rect 1869 10081 1903 10115
rect 7665 10081 7699 10115
rect 8309 10081 8343 10115
rect 8585 10081 8619 10115
rect 9689 10081 9723 10115
rect 9965 10081 9999 10115
rect 12909 10081 12943 10115
rect 13461 10081 13495 10115
rect 17233 10081 17267 10115
rect 17785 10081 17819 10115
rect 18613 10081 18647 10115
rect 21097 10081 21131 10115
rect 5181 10013 5215 10047
rect 6837 10013 6871 10047
rect 8493 10013 8527 10047
rect 9781 10013 9815 10047
rect 11529 10013 11563 10047
rect 18245 10013 18279 10047
rect 2237 9945 2271 9979
rect 5733 9945 5767 9979
rect 11897 9945 11931 9979
rect 6285 9877 6319 9911
rect 8125 9877 8159 9911
rect 10149 9877 10183 9911
rect 2329 9673 2363 9707
rect 13185 9673 13219 9707
rect 2789 9605 2823 9639
rect 5273 9605 5307 9639
rect 7389 9537 7423 9571
rect 9597 9537 9631 9571
rect 9689 9537 9723 9571
rect 12449 9537 12483 9571
rect 1777 9469 1811 9503
rect 2329 9469 2363 9503
rect 2973 9469 3007 9503
rect 4997 9469 5031 9503
rect 7573 9469 7607 9503
rect 8309 9469 8343 9503
rect 12081 9469 12115 9503
rect 12633 9469 12667 9503
rect 13093 9469 13127 9503
rect 14289 9469 14323 9503
rect 4721 9401 4755 9435
rect 4813 9333 4847 9367
rect 9781 9333 9815 9367
rect 10149 9333 10183 9367
rect 14473 9333 14507 9367
rect 2697 9129 2731 9163
rect 9965 9129 9999 9163
rect 12173 9129 12207 9163
rect 15209 9129 15243 9163
rect 15301 9129 15335 9163
rect 18613 9129 18647 9163
rect 5825 9061 5859 9095
rect 6009 9061 6043 9095
rect 17325 9061 17359 9095
rect 4721 8993 4755 9027
rect 4905 8993 4939 9027
rect 4997 8993 5031 9027
rect 6837 8993 6871 9027
rect 7021 8993 7055 9027
rect 8125 8993 8159 9027
rect 9597 8993 9631 9027
rect 9781 8993 9815 9027
rect 11529 8993 11563 9027
rect 11713 8993 11747 9027
rect 12357 8993 12391 9027
rect 16221 8993 16255 9027
rect 16773 8993 16807 9027
rect 17509 8993 17543 9027
rect 18245 8993 18279 9027
rect 5733 8925 5767 8959
rect 7389 8925 7423 8959
rect 9505 8925 9539 8959
rect 15393 8925 15427 8959
rect 16589 8925 16623 8959
rect 4537 8857 4571 8891
rect 18613 8857 18647 8891
rect 2789 8789 2823 8823
rect 6285 8789 6319 8823
rect 7941 8789 7975 8823
rect 14841 8789 14875 8823
rect 2145 8585 2179 8619
rect 9413 8585 9447 8619
rect 9597 8585 9631 8619
rect 17693 8585 17727 8619
rect 18705 8585 18739 8619
rect 19165 8585 19199 8619
rect 1593 8517 1627 8551
rect 14565 8517 14599 8551
rect 15025 8517 15059 8551
rect 2605 8449 2639 8483
rect 2697 8449 2731 8483
rect 3341 8449 3375 8483
rect 3893 8449 3927 8483
rect 7113 8449 7147 8483
rect 9413 8449 9447 8483
rect 9597 8449 9631 8483
rect 14197 8449 14231 8483
rect 17325 8449 17359 8483
rect 1409 8381 1443 8415
rect 2513 8381 2547 8415
rect 7573 8381 7607 8415
rect 8309 8381 8343 8415
rect 9505 8381 9539 8415
rect 12081 8381 12115 8415
rect 15209 8381 15243 8415
rect 17693 8381 17727 8415
rect 18153 8381 18187 8415
rect 18705 8381 18739 8415
rect 19349 8381 19383 8415
rect 21097 8381 21131 8415
rect 3801 8313 3835 8347
rect 8217 8313 8251 8347
rect 12265 8313 12299 8347
rect 9873 8245 9907 8279
rect 12449 8245 12483 8279
rect 14565 8245 14599 8279
rect 20913 8245 20947 8279
rect 12817 8041 12851 8075
rect 18429 8041 18463 8075
rect 8033 7973 8067 8007
rect 15209 7973 15243 8007
rect 16405 7973 16439 8007
rect 18245 7973 18279 8007
rect 2145 7905 2179 7939
rect 2697 7905 2731 7939
rect 7757 7905 7791 7939
rect 9873 7905 9907 7939
rect 14749 7905 14783 7939
rect 15301 7905 15335 7939
rect 16221 7905 16255 7939
rect 12633 7837 12667 7871
rect 12725 7837 12759 7871
rect 2697 7701 2731 7735
rect 9781 7701 9815 7735
rect 13185 7701 13219 7735
rect 3801 7497 3835 7531
rect 12817 7497 12851 7531
rect 13645 7497 13679 7531
rect 4721 7361 4755 7395
rect 8125 7361 8159 7395
rect 13277 7361 13311 7395
rect 7757 7293 7791 7327
rect 8585 7293 8619 7327
rect 9505 7293 9539 7327
rect 9965 7293 9999 7327
rect 10701 7293 10735 7327
rect 12265 7293 12299 7327
rect 12817 7293 12851 7327
rect 13645 7293 13679 7327
rect 14105 7293 14139 7327
rect 14289 7293 14323 7327
rect 3893 7225 3927 7259
rect 5181 7225 5215 7259
rect 5273 7225 5307 7259
rect 5733 7225 5767 7259
rect 7941 7225 7975 7259
rect 9229 7225 9263 7259
rect 10885 7225 10919 7259
rect 5917 7157 5951 7191
rect 7849 6953 7883 6987
rect 10885 6953 10919 6987
rect 17785 6953 17819 6987
rect 4905 6885 4939 6919
rect 5733 6885 5767 6919
rect 8217 6885 8251 6919
rect 10333 6885 10367 6919
rect 4261 6817 4295 6851
rect 5181 6817 5215 6851
rect 5641 6817 5675 6851
rect 6193 6817 6227 6851
rect 8309 6817 8343 6851
rect 9873 6817 9907 6851
rect 10425 6817 10459 6851
rect 11069 6817 11103 6851
rect 15945 6817 15979 6851
rect 16037 6817 16071 6851
rect 17785 6817 17819 6851
rect 17969 6817 18003 6851
rect 8493 6749 8527 6783
rect 16221 6749 16255 6783
rect 17601 6749 17635 6783
rect 15577 6613 15611 6647
rect 5917 6341 5951 6375
rect 6837 6341 6871 6375
rect 10241 6341 10275 6375
rect 5549 6273 5583 6307
rect 9873 6273 9907 6307
rect 14657 6273 14691 6307
rect 17325 6273 17359 6307
rect 3490 6205 3524 6239
rect 7021 6205 7055 6239
rect 15025 6205 15059 6239
rect 17509 6205 17543 6239
rect 17693 6205 17727 6239
rect 17877 6205 17911 6239
rect 18429 6205 18463 6239
rect 18705 6205 18739 6239
rect 18889 6205 18923 6239
rect 3387 6069 3421 6103
rect 5917 6069 5951 6103
rect 10241 6069 10275 6103
rect 15025 6069 15059 6103
rect 18705 6069 18739 6103
rect 6929 5865 6963 5899
rect 16129 5865 16163 5899
rect 18613 5865 18647 5899
rect 20913 5865 20947 5899
rect 1593 5797 1627 5831
rect 13461 5797 13495 5831
rect 15209 5797 15243 5831
rect 2789 5729 2823 5763
rect 7021 5729 7055 5763
rect 12725 5729 12759 5763
rect 14749 5729 14783 5763
rect 15301 5729 15335 5763
rect 16497 5729 16531 5763
rect 17785 5729 17819 5763
rect 17969 5729 18003 5763
rect 18705 5729 18739 5763
rect 21097 5729 21131 5763
rect 16589 5661 16623 5695
rect 16773 5661 16807 5695
rect 17417 5661 17451 5695
rect 17601 5661 17635 5695
rect 13277 5593 13311 5627
rect 1501 5525 1535 5559
rect 2697 5525 2731 5559
rect 12633 5525 12667 5559
rect 8125 5321 8159 5355
rect 13001 5321 13035 5355
rect 13829 5321 13863 5355
rect 15117 5321 15151 5355
rect 17325 5321 17359 5355
rect 18613 5321 18647 5355
rect 3249 5185 3283 5219
rect 13461 5185 13495 5219
rect 17877 5185 17911 5219
rect 2973 5117 3007 5151
rect 4997 5117 5031 5151
rect 7573 5117 7607 5151
rect 8125 5117 8159 5151
rect 10241 5117 10275 5151
rect 12449 5117 12483 5151
rect 13001 5117 13035 5151
rect 13829 5117 13863 5151
rect 14473 5117 14507 5151
rect 14657 5117 14691 5151
rect 15301 5117 15335 5151
rect 18521 5117 18555 5151
rect 10977 5049 11011 5083
rect 11161 5049 11195 5083
rect 17693 4981 17727 5015
rect 17785 4981 17819 5015
rect 7849 4777 7883 4811
rect 17969 4777 18003 4811
rect 18429 4777 18463 4811
rect 8217 4709 8251 4743
rect 11161 4709 11195 4743
rect 4997 4641 5031 4675
rect 7021 4641 7055 4675
rect 10517 4641 10551 4675
rect 11437 4641 11471 4675
rect 18337 4641 18371 4675
rect 6745 4573 6779 4607
rect 8309 4573 8343 4607
rect 8493 4573 8527 4607
rect 18613 4573 18647 4607
rect 8309 4233 8343 4267
rect 12173 4233 12207 4267
rect 18416 4233 18450 4267
rect 15393 4165 15427 4199
rect 7941 4097 7975 4131
rect 9597 4097 9631 4131
rect 18153 4097 18187 4131
rect 8309 4029 8343 4063
rect 8769 4029 8803 4063
rect 9873 4029 9907 4063
rect 15577 3961 15611 3995
rect 8953 3893 8987 3927
rect 9781 3893 9815 3927
rect 10241 3893 10275 3927
rect 12081 3893 12115 3927
rect 14749 3893 14783 3927
rect 14841 3893 14875 3927
rect 20177 3893 20211 3927
rect 8585 3689 8619 3723
rect 11253 3689 11287 3723
rect 11345 3689 11379 3723
rect 12725 3689 12759 3723
rect 15945 3689 15979 3723
rect 4353 3621 4387 3655
rect 15025 3621 15059 3655
rect 1409 3553 1443 3587
rect 6929 3553 6963 3587
rect 9689 3553 9723 3587
rect 12265 3553 12299 3587
rect 12909 3553 12943 3587
rect 14933 3553 14967 3587
rect 15485 3553 15519 3587
rect 15945 3553 15979 3587
rect 21097 3553 21131 3587
rect 8217 3485 8251 3519
rect 11437 3485 11471 3519
rect 16313 3485 16347 3519
rect 8585 3417 8619 3451
rect 9505 3417 9539 3451
rect 1593 3349 1627 3383
rect 4445 3349 4479 3383
rect 6745 3349 6779 3383
rect 10885 3349 10919 3383
rect 12081 3349 12115 3383
rect 20913 3349 20947 3383
rect 9045 3145 9079 3179
rect 10057 3145 10091 3179
rect 11161 3145 11195 3179
rect 12173 3145 12207 3179
rect 14657 3145 14691 3179
rect 15577 3145 15611 3179
rect 20913 3145 20947 3179
rect 8493 3009 8527 3043
rect 13185 3009 13219 3043
rect 16037 3009 16071 3043
rect 16129 3009 16163 3043
rect 17325 3009 17359 3043
rect 17601 3009 17635 3043
rect 1409 2941 1443 2975
rect 8585 2941 8619 2975
rect 8677 2941 8711 2975
rect 9505 2941 9539 2975
rect 10057 2941 10091 2975
rect 10609 2941 10643 2975
rect 11161 2941 11195 2975
rect 12081 2941 12115 2975
rect 14289 2941 14323 2975
rect 14657 2941 14691 2975
rect 19349 2941 19383 2975
rect 21097 2941 21131 2975
rect 15945 2873 15979 2907
rect 1593 2805 1627 2839
rect 13369 2805 13403 2839
rect 13461 2805 13495 2839
rect 13829 2805 13863 2839
rect 4445 2601 4479 2635
rect 5733 2601 5767 2635
rect 7021 2601 7055 2635
rect 9781 2601 9815 2635
rect 11345 2601 11379 2635
rect 12909 2601 12943 2635
rect 14933 2601 14967 2635
rect 18889 2601 18923 2635
rect 2053 2533 2087 2567
rect 17877 2533 17911 2567
rect 20913 2533 20947 2567
rect 4261 2465 4295 2499
rect 5549 2465 5583 2499
rect 7113 2465 7147 2499
rect 9597 2465 9631 2499
rect 10333 2465 10367 2499
rect 10977 2465 11011 2499
rect 11345 2465 11379 2499
rect 12725 2465 12759 2499
rect 13369 2465 13403 2499
rect 13921 2465 13955 2499
rect 15117 2465 15151 2499
rect 15669 2465 15703 2499
rect 17693 2465 17727 2499
rect 19073 2465 19107 2499
rect 16129 2397 16163 2431
rect 1869 2329 1903 2363
rect 10517 2329 10551 2363
rect 20729 2329 20763 2363
rect 13921 2261 13955 2295
<< metal1 >>
rect 1104 22874 21804 22896
rect 1104 22822 4432 22874
rect 4484 22822 4496 22874
rect 4548 22822 4560 22874
rect 4612 22822 4624 22874
rect 4676 22822 11332 22874
rect 11384 22822 11396 22874
rect 11448 22822 11460 22874
rect 11512 22822 11524 22874
rect 11576 22822 18232 22874
rect 18284 22822 18296 22874
rect 18348 22822 18360 22874
rect 18412 22822 18424 22874
rect 18476 22822 21804 22874
rect 1104 22800 21804 22822
rect 1486 22760 1492 22772
rect 1447 22732 1492 22760
rect 1486 22720 1492 22732
rect 1544 22720 1550 22772
rect 2961 22695 3019 22701
rect 2961 22661 2973 22695
rect 3007 22692 3019 22695
rect 5442 22692 5448 22704
rect 3007 22664 5448 22692
rect 3007 22661 3019 22664
rect 2961 22655 3019 22661
rect 5442 22652 5448 22664
rect 5500 22652 5506 22704
rect 8021 22695 8079 22701
rect 8021 22661 8033 22695
rect 8067 22692 8079 22695
rect 11054 22692 11060 22704
rect 8067 22664 11060 22692
rect 8067 22661 8079 22664
rect 8021 22655 8079 22661
rect 11054 22652 11060 22664
rect 11112 22652 11118 22704
rect 934 22516 940 22568
rect 992 22556 998 22568
rect 2317 22559 2375 22565
rect 2317 22556 2329 22559
rect 992 22528 2329 22556
rect 992 22516 998 22528
rect 2317 22525 2329 22528
rect 2363 22525 2375 22559
rect 2317 22519 2375 22525
rect 2774 22516 2780 22568
rect 2832 22556 2838 22568
rect 4706 22556 4712 22568
rect 2832 22528 2877 22556
rect 4667 22528 4712 22556
rect 2832 22516 2838 22528
rect 4706 22516 4712 22528
rect 4764 22516 4770 22568
rect 4798 22516 4804 22568
rect 4856 22556 4862 22568
rect 5353 22559 5411 22565
rect 5353 22556 5365 22559
rect 4856 22528 5365 22556
rect 4856 22516 4862 22528
rect 5353 22525 5365 22528
rect 5399 22525 5411 22559
rect 5353 22519 5411 22525
rect 5994 22516 6000 22568
rect 6052 22556 6058 22568
rect 7101 22559 7159 22565
rect 7101 22556 7113 22559
rect 6052 22528 7113 22556
rect 6052 22516 6058 22528
rect 7101 22525 7113 22528
rect 7147 22525 7159 22559
rect 7834 22556 7840 22568
rect 7795 22528 7840 22556
rect 7101 22519 7159 22525
rect 7834 22516 7840 22528
rect 7892 22516 7898 22568
rect 9674 22556 9680 22568
rect 9635 22528 9680 22556
rect 9674 22516 9680 22528
rect 9732 22516 9738 22568
rect 11698 22516 11704 22568
rect 11756 22556 11762 22568
rect 12437 22559 12495 22565
rect 12437 22556 12449 22559
rect 11756 22528 12449 22556
rect 11756 22516 11762 22528
rect 12437 22525 12449 22528
rect 12483 22525 12495 22559
rect 12894 22556 12900 22568
rect 12855 22528 12900 22556
rect 12437 22519 12495 22525
rect 12894 22516 12900 22528
rect 12952 22516 12958 22568
rect 14734 22516 14740 22568
rect 14792 22556 14798 22568
rect 15105 22559 15163 22565
rect 15105 22556 15117 22559
rect 14792 22528 15117 22556
rect 14792 22516 14798 22528
rect 15105 22525 15117 22528
rect 15151 22525 15163 22559
rect 15105 22519 15163 22525
rect 16574 22516 16580 22568
rect 16632 22556 16638 22568
rect 16669 22559 16727 22565
rect 16669 22556 16681 22559
rect 16632 22528 16681 22556
rect 16632 22516 16638 22528
rect 16669 22525 16681 22528
rect 16715 22525 16727 22559
rect 16669 22519 16727 22525
rect 17954 22516 17960 22568
rect 18012 22556 18018 22568
rect 18141 22559 18199 22565
rect 18141 22556 18153 22559
rect 18012 22528 18153 22556
rect 18012 22516 18018 22528
rect 18141 22525 18153 22528
rect 18187 22525 18199 22559
rect 18141 22519 18199 22525
rect 19337 22559 19395 22565
rect 19337 22525 19349 22559
rect 19383 22556 19395 22559
rect 19794 22556 19800 22568
rect 19383 22528 19800 22556
rect 19383 22525 19395 22528
rect 19337 22519 19395 22525
rect 19794 22516 19800 22528
rect 19852 22516 19858 22568
rect 21085 22559 21143 22565
rect 21085 22525 21097 22559
rect 21131 22556 21143 22559
rect 21634 22556 21640 22568
rect 21131 22528 21640 22556
rect 21131 22525 21143 22528
rect 21085 22519 21143 22525
rect 21634 22516 21640 22528
rect 21692 22516 21698 22568
rect 1578 22488 1584 22500
rect 1539 22460 1584 22488
rect 1578 22448 1584 22460
rect 1636 22448 1642 22500
rect 2038 22380 2044 22432
rect 2096 22420 2102 22432
rect 2133 22423 2191 22429
rect 2133 22420 2145 22423
rect 2096 22392 2145 22420
rect 2096 22380 2102 22392
rect 2133 22389 2145 22392
rect 2179 22389 2191 22423
rect 4890 22420 4896 22432
rect 4851 22392 4896 22420
rect 2133 22383 2191 22389
rect 4890 22380 4896 22392
rect 4948 22380 4954 22432
rect 5537 22423 5595 22429
rect 5537 22389 5549 22423
rect 5583 22420 5595 22423
rect 6178 22420 6184 22432
rect 5583 22392 6184 22420
rect 5583 22389 5595 22392
rect 5537 22383 5595 22389
rect 6178 22380 6184 22392
rect 6236 22380 6242 22432
rect 6917 22423 6975 22429
rect 6917 22389 6929 22423
rect 6963 22420 6975 22423
rect 7006 22420 7012 22432
rect 6963 22392 7012 22420
rect 6963 22389 6975 22392
rect 6917 22383 6975 22389
rect 7006 22380 7012 22392
rect 7064 22380 7070 22432
rect 9861 22423 9919 22429
rect 9861 22389 9873 22423
rect 9907 22420 9919 22423
rect 10594 22420 10600 22432
rect 9907 22392 10600 22420
rect 9907 22389 9919 22392
rect 9861 22383 9919 22389
rect 10594 22380 10600 22392
rect 10652 22380 10658 22432
rect 12253 22423 12311 22429
rect 12253 22389 12265 22423
rect 12299 22420 12311 22423
rect 12342 22420 12348 22432
rect 12299 22392 12348 22420
rect 12299 22389 12311 22392
rect 12253 22383 12311 22389
rect 12342 22380 12348 22392
rect 12400 22380 12406 22432
rect 12710 22380 12716 22432
rect 12768 22420 12774 22432
rect 13081 22423 13139 22429
rect 13081 22420 13093 22423
rect 12768 22392 13093 22420
rect 12768 22380 12774 22392
rect 13081 22389 13093 22392
rect 13127 22389 13139 22423
rect 13081 22383 13139 22389
rect 14642 22380 14648 22432
rect 14700 22420 14706 22432
rect 14921 22423 14979 22429
rect 14921 22420 14933 22423
rect 14700 22392 14933 22420
rect 14700 22380 14706 22392
rect 14921 22389 14933 22392
rect 14967 22389 14979 22423
rect 14921 22383 14979 22389
rect 16298 22380 16304 22432
rect 16356 22420 16362 22432
rect 16485 22423 16543 22429
rect 16485 22420 16497 22423
rect 16356 22392 16497 22420
rect 16356 22380 16362 22392
rect 16485 22389 16497 22392
rect 16531 22389 16543 22423
rect 17954 22420 17960 22432
rect 17915 22392 17960 22420
rect 16485 22383 16543 22389
rect 17954 22380 17960 22392
rect 18012 22380 18018 22432
rect 19150 22420 19156 22432
rect 19111 22392 19156 22420
rect 19150 22380 19156 22392
rect 19208 22380 19214 22432
rect 20901 22423 20959 22429
rect 20901 22389 20913 22423
rect 20947 22420 20959 22423
rect 21174 22420 21180 22432
rect 20947 22392 21180 22420
rect 20947 22389 20959 22392
rect 20901 22383 20959 22389
rect 21174 22380 21180 22392
rect 21232 22380 21238 22432
rect 1104 22330 21804 22352
rect 1104 22278 7882 22330
rect 7934 22278 7946 22330
rect 7998 22278 8010 22330
rect 8062 22278 8074 22330
rect 8126 22278 14782 22330
rect 14834 22278 14846 22330
rect 14898 22278 14910 22330
rect 14962 22278 14974 22330
rect 15026 22278 21804 22330
rect 1104 22256 21804 22278
rect 10870 22148 10876 22160
rect 10783 22120 10876 22148
rect 10870 22108 10876 22120
rect 10928 22148 10934 22160
rect 11882 22148 11888 22160
rect 10928 22120 11888 22148
rect 10928 22108 10934 22120
rect 11882 22108 11888 22120
rect 11940 22108 11946 22160
rect 4982 22080 4988 22092
rect 4943 22052 4988 22080
rect 4982 22040 4988 22052
rect 5040 22040 5046 22092
rect 5074 22040 5080 22092
rect 5132 22080 5138 22092
rect 5353 22083 5411 22089
rect 5132 22052 5177 22080
rect 5132 22040 5138 22052
rect 5353 22049 5365 22083
rect 5399 22080 5411 22083
rect 5534 22080 5540 22092
rect 5399 22052 5540 22080
rect 5399 22049 5411 22052
rect 5353 22043 5411 22049
rect 5534 22040 5540 22052
rect 5592 22040 5598 22092
rect 7561 22083 7619 22089
rect 7561 22049 7573 22083
rect 7607 22080 7619 22083
rect 9861 22083 9919 22089
rect 9861 22080 9873 22083
rect 7607 22052 9873 22080
rect 7607 22049 7619 22052
rect 7561 22043 7619 22049
rect 9861 22049 9873 22052
rect 9907 22080 9919 22083
rect 10318 22080 10324 22092
rect 9907 22052 10324 22080
rect 9907 22049 9919 22052
rect 9861 22043 9919 22049
rect 4706 21972 4712 22024
rect 4764 22012 4770 22024
rect 7576 22012 7604 22043
rect 10318 22040 10324 22052
rect 10376 22040 10382 22092
rect 11057 22083 11115 22089
rect 11057 22049 11069 22083
rect 11103 22080 11115 22083
rect 11698 22080 11704 22092
rect 11103 22052 11704 22080
rect 11103 22049 11115 22052
rect 11057 22043 11115 22049
rect 11698 22040 11704 22052
rect 11756 22040 11762 22092
rect 11974 22080 11980 22092
rect 11935 22052 11980 22080
rect 11974 22040 11980 22052
rect 12032 22040 12038 22092
rect 12158 22089 12164 22092
rect 12115 22083 12164 22089
rect 12115 22049 12127 22083
rect 12161 22049 12164 22083
rect 12115 22043 12164 22049
rect 12158 22040 12164 22043
rect 12216 22040 12222 22092
rect 12894 22080 12900 22092
rect 12807 22052 12900 22080
rect 12894 22040 12900 22052
rect 12952 22080 12958 22092
rect 15381 22083 15439 22089
rect 15381 22080 15393 22083
rect 12952 22052 15393 22080
rect 12952 22040 12958 22052
rect 15381 22049 15393 22052
rect 15427 22080 15439 22083
rect 17494 22080 17500 22092
rect 15427 22052 17500 22080
rect 15427 22049 15439 22052
rect 15381 22043 15439 22049
rect 17494 22040 17500 22052
rect 17552 22080 17558 22092
rect 18325 22083 18383 22089
rect 18325 22080 18337 22083
rect 17552 22052 18337 22080
rect 17552 22040 17558 22052
rect 18325 22049 18337 22052
rect 18371 22080 18383 22083
rect 19981 22083 20039 22089
rect 19981 22080 19993 22083
rect 18371 22052 19993 22080
rect 18371 22049 18383 22052
rect 18325 22043 18383 22049
rect 19981 22049 19993 22052
rect 20027 22080 20039 22083
rect 20530 22080 20536 22092
rect 20027 22052 20536 22080
rect 20027 22049 20039 22052
rect 19981 22043 20039 22049
rect 20530 22040 20536 22052
rect 20588 22040 20594 22092
rect 21082 22080 21088 22092
rect 21043 22052 21088 22080
rect 21082 22040 21088 22052
rect 21140 22040 21146 22092
rect 4764 21984 7604 22012
rect 4764 21972 4770 21984
rect 15286 21904 15292 21956
rect 15344 21944 15350 21956
rect 20901 21947 20959 21953
rect 20901 21944 20913 21947
rect 15344 21916 20913 21944
rect 15344 21904 15350 21916
rect 20901 21913 20913 21916
rect 20947 21913 20959 21947
rect 20901 21907 20959 21913
rect 4154 21836 4160 21888
rect 4212 21876 4218 21888
rect 4801 21879 4859 21885
rect 4801 21876 4813 21879
rect 4212 21848 4813 21876
rect 4212 21836 4218 21848
rect 4801 21845 4813 21848
rect 4847 21845 4859 21879
rect 5258 21876 5264 21888
rect 5219 21848 5264 21876
rect 4801 21839 4859 21845
rect 5258 21836 5264 21848
rect 5316 21836 5322 21888
rect 7742 21876 7748 21888
rect 7703 21848 7748 21876
rect 7742 21836 7748 21848
rect 7800 21836 7806 21888
rect 10042 21876 10048 21888
rect 10003 21848 10048 21876
rect 10042 21836 10048 21848
rect 10100 21836 10106 21888
rect 10686 21876 10692 21888
rect 10647 21848 10692 21876
rect 10686 21836 10692 21848
rect 10744 21836 10750 21888
rect 12250 21876 12256 21888
rect 12211 21848 12256 21876
rect 12250 21836 12256 21848
rect 12308 21836 12314 21888
rect 12713 21879 12771 21885
rect 12713 21845 12725 21879
rect 12759 21876 12771 21879
rect 12802 21876 12808 21888
rect 12759 21848 12808 21876
rect 12759 21845 12771 21848
rect 12713 21839 12771 21845
rect 12802 21836 12808 21848
rect 12860 21836 12866 21888
rect 15194 21876 15200 21888
rect 15155 21848 15200 21876
rect 15194 21836 15200 21848
rect 15252 21836 15258 21888
rect 18509 21879 18567 21885
rect 18509 21845 18521 21879
rect 18555 21876 18567 21879
rect 18690 21876 18696 21888
rect 18555 21848 18696 21876
rect 18555 21845 18567 21848
rect 18509 21839 18567 21845
rect 18690 21836 18696 21848
rect 18748 21836 18754 21888
rect 20070 21836 20076 21888
rect 20128 21876 20134 21888
rect 20165 21879 20223 21885
rect 20165 21876 20177 21879
rect 20128 21848 20177 21876
rect 20128 21836 20134 21848
rect 20165 21845 20177 21848
rect 20211 21845 20223 21879
rect 20165 21839 20223 21845
rect 1104 21786 21804 21808
rect 1104 21734 4432 21786
rect 4484 21734 4496 21786
rect 4548 21734 4560 21786
rect 4612 21734 4624 21786
rect 4676 21734 11332 21786
rect 11384 21734 11396 21786
rect 11448 21734 11460 21786
rect 11512 21734 11524 21786
rect 11576 21734 18232 21786
rect 18284 21734 18296 21786
rect 18348 21734 18360 21786
rect 18412 21734 18424 21786
rect 18476 21734 21804 21786
rect 1104 21712 21804 21734
rect 1578 21632 1584 21684
rect 1636 21672 1642 21684
rect 1765 21675 1823 21681
rect 1765 21672 1777 21675
rect 1636 21644 1777 21672
rect 1636 21632 1642 21644
rect 1765 21641 1777 21644
rect 1811 21641 1823 21675
rect 10870 21672 10876 21684
rect 10831 21644 10876 21672
rect 1765 21635 1823 21641
rect 10870 21632 10876 21644
rect 10928 21632 10934 21684
rect 8202 21564 8208 21616
rect 8260 21604 8266 21616
rect 8573 21607 8631 21613
rect 8573 21604 8585 21607
rect 8260 21576 8585 21604
rect 8260 21564 8266 21576
rect 8573 21573 8585 21576
rect 8619 21573 8631 21607
rect 8573 21567 8631 21573
rect 20162 21564 20168 21616
rect 20220 21604 20226 21616
rect 20220 21576 21036 21604
rect 20220 21564 20226 21576
rect 4154 21536 4160 21548
rect 4115 21508 4160 21536
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 9122 21536 9128 21548
rect 6840 21508 9128 21536
rect 1949 21471 2007 21477
rect 1949 21437 1961 21471
rect 1995 21468 2007 21471
rect 2498 21468 2504 21480
rect 1995 21440 2504 21468
rect 1995 21437 2007 21440
rect 1949 21431 2007 21437
rect 2498 21428 2504 21440
rect 2556 21468 2562 21480
rect 6840 21477 6868 21508
rect 9122 21496 9128 21508
rect 9180 21496 9186 21548
rect 9401 21539 9459 21545
rect 9401 21505 9413 21539
rect 9447 21536 9459 21539
rect 10686 21536 10692 21548
rect 9447 21508 10692 21536
rect 9447 21505 9459 21508
rect 9401 21499 9459 21505
rect 10686 21496 10692 21508
rect 10744 21496 10750 21548
rect 12250 21496 12256 21548
rect 12308 21536 12314 21548
rect 13541 21539 13599 21545
rect 13541 21536 13553 21539
rect 12308 21508 13553 21536
rect 12308 21496 12314 21508
rect 13541 21505 13553 21508
rect 13587 21505 13599 21539
rect 16025 21539 16083 21545
rect 16025 21536 16037 21539
rect 13541 21499 13599 21505
rect 13832 21508 16037 21536
rect 13832 21477 13860 21508
rect 16025 21505 16037 21508
rect 16071 21536 16083 21539
rect 16206 21536 16212 21548
rect 16071 21508 16212 21536
rect 16071 21505 16083 21508
rect 16025 21499 16083 21505
rect 16206 21496 16212 21508
rect 16264 21536 16270 21548
rect 17405 21539 17463 21545
rect 17405 21536 17417 21539
rect 16264 21508 17417 21536
rect 16264 21496 16270 21508
rect 17405 21505 17417 21508
rect 17451 21536 17463 21539
rect 19058 21536 19064 21548
rect 17451 21508 19064 21536
rect 17451 21505 17463 21508
rect 17405 21499 17463 21505
rect 19058 21496 19064 21508
rect 19116 21496 19122 21548
rect 21008 21545 21036 21576
rect 20993 21539 21051 21545
rect 20993 21505 21005 21539
rect 21039 21505 21051 21539
rect 20993 21499 21051 21505
rect 3881 21471 3939 21477
rect 3881 21468 3893 21471
rect 2556 21440 3893 21468
rect 2556 21428 2562 21440
rect 3881 21437 3893 21440
rect 3927 21437 3939 21471
rect 6825 21471 6883 21477
rect 6825 21468 6837 21471
rect 3881 21431 3939 21437
rect 5460 21440 6837 21468
rect 3896 21332 3924 21431
rect 4890 21360 4896 21412
rect 4948 21360 4954 21412
rect 5460 21332 5488 21440
rect 6825 21437 6837 21440
rect 6871 21437 6883 21471
rect 6825 21431 6883 21437
rect 13817 21471 13875 21477
rect 13817 21437 13829 21471
rect 13863 21437 13875 21471
rect 20162 21468 20168 21480
rect 20123 21440 20168 21468
rect 13817 21431 13875 21437
rect 7101 21403 7159 21409
rect 7101 21369 7113 21403
rect 7147 21400 7159 21403
rect 7190 21400 7196 21412
rect 7147 21372 7196 21400
rect 7147 21369 7159 21372
rect 7101 21363 7159 21369
rect 7190 21360 7196 21372
rect 7248 21360 7254 21412
rect 7742 21360 7748 21412
rect 7800 21360 7806 21412
rect 10042 21360 10048 21412
rect 10100 21360 10106 21412
rect 11900 21372 12204 21400
rect 3896 21304 5488 21332
rect 5534 21292 5540 21344
rect 5592 21332 5598 21344
rect 5629 21335 5687 21341
rect 5629 21332 5641 21335
rect 5592 21304 5641 21332
rect 5592 21292 5598 21304
rect 5629 21301 5641 21304
rect 5675 21301 5687 21335
rect 5629 21295 5687 21301
rect 9122 21292 9128 21344
rect 9180 21332 9186 21344
rect 11900 21332 11928 21372
rect 12066 21332 12072 21344
rect 9180 21304 11928 21332
rect 12027 21304 12072 21332
rect 9180 21292 9186 21304
rect 12066 21292 12072 21304
rect 12124 21292 12130 21344
rect 12176 21332 12204 21372
rect 12802 21360 12808 21412
rect 12860 21360 12866 21412
rect 13832 21332 13860 21431
rect 20162 21428 20168 21440
rect 20220 21428 20226 21480
rect 20349 21471 20407 21477
rect 20349 21437 20361 21471
rect 20395 21437 20407 21471
rect 20349 21431 20407 21437
rect 20901 21471 20959 21477
rect 20901 21437 20913 21471
rect 20947 21468 20959 21471
rect 21082 21468 21088 21480
rect 20947 21440 21088 21468
rect 20947 21437 20959 21440
rect 20901 21431 20959 21437
rect 15194 21360 15200 21412
rect 15252 21360 15258 21412
rect 15746 21400 15752 21412
rect 15707 21372 15752 21400
rect 15746 21360 15752 21372
rect 15804 21360 15810 21412
rect 17681 21403 17739 21409
rect 17681 21369 17693 21403
rect 17727 21400 17739 21403
rect 17954 21400 17960 21412
rect 17727 21372 17960 21400
rect 17727 21369 17739 21372
rect 17681 21363 17739 21369
rect 17954 21360 17960 21372
rect 18012 21360 18018 21412
rect 18690 21360 18696 21412
rect 18748 21360 18754 21412
rect 19797 21403 19855 21409
rect 19797 21400 19809 21403
rect 18984 21372 19809 21400
rect 14274 21332 14280 21344
rect 12176 21304 13860 21332
rect 14235 21304 14280 21332
rect 14274 21292 14280 21304
rect 14332 21292 14338 21344
rect 15470 21292 15476 21344
rect 15528 21332 15534 21344
rect 18984 21332 19012 21372
rect 19797 21369 19809 21372
rect 19843 21369 19855 21403
rect 20364 21400 20392 21431
rect 20916 21400 20944 21431
rect 21082 21428 21088 21440
rect 21140 21428 21146 21480
rect 20364 21372 20944 21400
rect 19797 21363 19855 21369
rect 15528 21304 19012 21332
rect 19153 21335 19211 21341
rect 15528 21292 15534 21304
rect 19153 21301 19165 21335
rect 19199 21332 19211 21335
rect 19334 21332 19340 21344
rect 19199 21304 19340 21332
rect 19199 21301 19211 21304
rect 19153 21295 19211 21301
rect 19334 21292 19340 21304
rect 19392 21292 19398 21344
rect 1104 21242 21804 21264
rect 1104 21190 7882 21242
rect 7934 21190 7946 21242
rect 7998 21190 8010 21242
rect 8062 21190 8074 21242
rect 8126 21190 14782 21242
rect 14834 21190 14846 21242
rect 14898 21190 14910 21242
rect 14962 21190 14974 21242
rect 15026 21190 21804 21242
rect 1104 21168 21804 21190
rect 4982 21088 4988 21140
rect 5040 21128 5046 21140
rect 5261 21131 5319 21137
rect 5261 21128 5273 21131
rect 5040 21100 5273 21128
rect 5040 21088 5046 21100
rect 5261 21097 5273 21100
rect 5307 21097 5319 21131
rect 7190 21128 7196 21140
rect 7151 21100 7196 21128
rect 5261 21091 5319 21097
rect 7190 21088 7196 21100
rect 7248 21088 7254 21140
rect 11698 21088 11704 21140
rect 11756 21128 11762 21140
rect 11974 21128 11980 21140
rect 11756 21100 11980 21128
rect 11756 21088 11762 21100
rect 11974 21088 11980 21100
rect 12032 21088 12038 21140
rect 12158 21088 12164 21140
rect 12216 21128 12222 21140
rect 15289 21131 15347 21137
rect 12216 21100 15148 21128
rect 12216 21088 12222 21100
rect 7466 21060 7472 21072
rect 7427 21032 7472 21060
rect 7466 21020 7472 21032
rect 7524 21020 7530 21072
rect 7650 21060 7656 21072
rect 7609 21032 7656 21060
rect 7650 21020 7656 21032
rect 7708 21069 7714 21072
rect 7708 21063 7757 21069
rect 7708 21029 7711 21063
rect 7745 21060 7757 21063
rect 8202 21060 8208 21072
rect 7745 21032 8208 21060
rect 7745 21029 7757 21032
rect 7708 21023 7757 21029
rect 7708 21020 7714 21023
rect 8202 21020 8208 21032
rect 8260 21020 8266 21072
rect 12066 21060 12072 21072
rect 12027 21032 12072 21060
rect 12066 21020 12072 21032
rect 12124 21020 12130 21072
rect 5353 20995 5411 21001
rect 5353 20961 5365 20995
rect 5399 20992 5411 20995
rect 5534 20992 5540 21004
rect 5399 20964 5540 20992
rect 5399 20961 5411 20964
rect 5353 20955 5411 20961
rect 5534 20952 5540 20964
rect 5592 20952 5598 21004
rect 7374 20992 7380 21004
rect 7335 20964 7380 20992
rect 7374 20952 7380 20964
rect 7432 20952 7438 21004
rect 7561 20995 7619 21001
rect 7561 20992 7573 20995
rect 7484 20964 7573 20992
rect 7101 20927 7159 20933
rect 7101 20893 7113 20927
rect 7147 20924 7159 20927
rect 7484 20924 7512 20964
rect 7561 20961 7573 20964
rect 7607 20961 7619 20995
rect 8297 20995 8355 21001
rect 8297 20992 8309 20995
rect 7561 20955 7619 20961
rect 7852 20964 8309 20992
rect 7852 20933 7880 20964
rect 8297 20961 8309 20964
rect 8343 20992 8355 20995
rect 8478 20992 8484 21004
rect 8343 20964 8484 20992
rect 8343 20961 8355 20964
rect 8297 20955 8355 20961
rect 8478 20952 8484 20964
rect 8536 20952 8542 21004
rect 11974 20952 11980 21004
rect 12032 20992 12038 21004
rect 12032 20964 12077 20992
rect 12032 20952 12038 20964
rect 12158 20952 12164 21004
rect 12216 20992 12222 21004
rect 12360 21001 12388 21100
rect 14274 21020 14280 21072
rect 14332 21060 14338 21072
rect 15013 21063 15071 21069
rect 15013 21060 15025 21063
rect 14332 21032 15025 21060
rect 14332 21020 14338 21032
rect 15013 21029 15025 21032
rect 15059 21029 15071 21063
rect 15013 21023 15071 21029
rect 15120 21001 15148 21100
rect 15289 21097 15301 21131
rect 15335 21128 15347 21131
rect 15746 21128 15752 21140
rect 15335 21100 15752 21128
rect 15335 21097 15347 21100
rect 15289 21091 15347 21097
rect 15746 21088 15752 21100
rect 15804 21088 15810 21140
rect 17218 21020 17224 21072
rect 17276 21020 17282 21072
rect 12345 20995 12403 21001
rect 12216 20964 12261 20992
rect 12216 20952 12222 20964
rect 12345 20961 12357 20995
rect 12391 20961 12403 20995
rect 12345 20955 12403 20961
rect 14737 20995 14795 21001
rect 14737 20961 14749 20995
rect 14783 20961 14795 20995
rect 14737 20955 14795 20961
rect 14921 20995 14979 21001
rect 14921 20961 14933 20995
rect 14967 20961 14979 20995
rect 14921 20955 14979 20961
rect 15105 20995 15163 21001
rect 15105 20961 15117 20995
rect 15151 20992 15163 20995
rect 15470 20992 15476 21004
rect 15151 20964 15476 20992
rect 15151 20961 15163 20964
rect 15105 20955 15163 20961
rect 7147 20896 7512 20924
rect 7837 20927 7895 20933
rect 7147 20893 7159 20896
rect 7101 20887 7159 20893
rect 7837 20893 7849 20927
rect 7883 20893 7895 20927
rect 7837 20887 7895 20893
rect 5074 20816 5080 20868
rect 5132 20856 5138 20868
rect 7852 20856 7880 20887
rect 5132 20828 7880 20856
rect 14752 20856 14780 20955
rect 14936 20924 14964 20955
rect 15470 20952 15476 20964
rect 15528 20952 15534 21004
rect 16206 20992 16212 21004
rect 16167 20964 16212 20992
rect 16206 20952 16212 20964
rect 16264 20952 16270 21004
rect 20806 20952 20812 21004
rect 20864 20992 20870 21004
rect 20901 20995 20959 21001
rect 20901 20992 20913 20995
rect 20864 20964 20913 20992
rect 20864 20952 20870 20964
rect 20901 20961 20913 20964
rect 20947 20961 20959 20995
rect 20901 20955 20959 20961
rect 15654 20924 15660 20936
rect 14936 20896 15660 20924
rect 15654 20884 15660 20896
rect 15712 20884 15718 20936
rect 16482 20924 16488 20936
rect 16443 20896 16488 20924
rect 16482 20884 16488 20896
rect 16540 20884 16546 20936
rect 15378 20856 15384 20868
rect 14752 20828 15384 20856
rect 5132 20816 5138 20828
rect 15378 20816 15384 20828
rect 15436 20816 15442 20868
rect 4982 20748 4988 20800
rect 5040 20788 5046 20800
rect 5258 20788 5264 20800
rect 5040 20760 5264 20788
rect 5040 20748 5046 20760
rect 5258 20748 5264 20760
rect 5316 20788 5322 20800
rect 7101 20791 7159 20797
rect 7101 20788 7113 20791
rect 5316 20760 7113 20788
rect 5316 20748 5322 20760
rect 7101 20757 7113 20760
rect 7147 20788 7159 20791
rect 8389 20791 8447 20797
rect 8389 20788 8401 20791
rect 7147 20760 8401 20788
rect 7147 20757 7159 20760
rect 7101 20751 7159 20757
rect 8389 20757 8401 20760
rect 8435 20757 8447 20791
rect 11790 20788 11796 20800
rect 11751 20760 11796 20788
rect 8389 20751 8447 20757
rect 11790 20748 11796 20760
rect 11848 20748 11854 20800
rect 15654 20748 15660 20800
rect 15712 20788 15718 20800
rect 17957 20791 18015 20797
rect 17957 20788 17969 20791
rect 15712 20760 17969 20788
rect 15712 20748 15718 20760
rect 17957 20757 17969 20760
rect 18003 20757 18015 20791
rect 17957 20751 18015 20757
rect 20622 20748 20628 20800
rect 20680 20788 20686 20800
rect 20993 20791 21051 20797
rect 20993 20788 21005 20791
rect 20680 20760 21005 20788
rect 20680 20748 20686 20760
rect 20993 20757 21005 20760
rect 21039 20757 21051 20791
rect 20993 20751 21051 20757
rect 1104 20698 21804 20720
rect 1104 20646 4432 20698
rect 4484 20646 4496 20698
rect 4548 20646 4560 20698
rect 4612 20646 4624 20698
rect 4676 20646 11332 20698
rect 11384 20646 11396 20698
rect 11448 20646 11460 20698
rect 11512 20646 11524 20698
rect 11576 20646 18232 20698
rect 18284 20646 18296 20698
rect 18348 20646 18360 20698
rect 18412 20646 18424 20698
rect 18476 20646 21804 20698
rect 1104 20624 21804 20646
rect 7374 20544 7380 20596
rect 7432 20584 7438 20596
rect 7745 20587 7803 20593
rect 7745 20584 7757 20587
rect 7432 20556 7757 20584
rect 7432 20544 7438 20556
rect 7745 20553 7757 20556
rect 7791 20553 7803 20587
rect 7745 20547 7803 20553
rect 12066 20544 12072 20596
rect 12124 20584 12130 20596
rect 12124 20556 12940 20584
rect 12124 20544 12130 20556
rect 11149 20519 11207 20525
rect 11149 20485 11161 20519
rect 11195 20516 11207 20519
rect 12158 20516 12164 20528
rect 11195 20488 12164 20516
rect 11195 20485 11207 20488
rect 11149 20479 11207 20485
rect 12158 20476 12164 20488
rect 12216 20516 12222 20528
rect 12526 20516 12532 20528
rect 12216 20488 12296 20516
rect 12487 20488 12532 20516
rect 12216 20476 12222 20488
rect 2498 20448 2504 20460
rect 2459 20420 2504 20448
rect 2498 20408 2504 20420
rect 2556 20408 2562 20460
rect 9122 20408 9128 20460
rect 9180 20448 9186 20460
rect 9401 20451 9459 20457
rect 9401 20448 9413 20451
rect 9180 20420 9413 20448
rect 9180 20408 9186 20420
rect 9401 20417 9413 20420
rect 9447 20417 9459 20451
rect 9401 20411 9459 20417
rect 9677 20451 9735 20457
rect 9677 20417 9689 20451
rect 9723 20448 9735 20451
rect 11790 20448 11796 20460
rect 9723 20420 11796 20448
rect 9723 20417 9735 20420
rect 9677 20411 9735 20417
rect 11790 20408 11796 20420
rect 11848 20408 11854 20460
rect 1394 20380 1400 20392
rect 1355 20352 1400 20380
rect 1394 20340 1400 20352
rect 1452 20340 1458 20392
rect 5258 20380 5264 20392
rect 5219 20352 5264 20380
rect 5258 20340 5264 20352
rect 5316 20340 5322 20392
rect 5445 20383 5503 20389
rect 5445 20349 5457 20383
rect 5491 20380 5503 20383
rect 5534 20380 5540 20392
rect 5491 20352 5540 20380
rect 5491 20349 5503 20352
rect 5445 20343 5503 20349
rect 5534 20340 5540 20352
rect 5592 20380 5598 20392
rect 5994 20380 6000 20392
rect 5592 20352 6000 20380
rect 5592 20340 5598 20352
rect 5994 20340 6000 20352
rect 6052 20340 6058 20392
rect 7650 20380 7656 20392
rect 7611 20352 7656 20380
rect 7650 20340 7656 20352
rect 7708 20340 7714 20392
rect 7742 20340 7748 20392
rect 7800 20380 7806 20392
rect 7837 20383 7895 20389
rect 7837 20380 7849 20383
rect 7800 20352 7849 20380
rect 7800 20340 7806 20352
rect 7837 20349 7849 20352
rect 7883 20349 7895 20383
rect 7837 20343 7895 20349
rect 11882 20340 11888 20392
rect 11940 20380 11946 20392
rect 12268 20389 12296 20488
rect 12526 20476 12532 20488
rect 12584 20476 12590 20528
rect 12912 20389 12940 20556
rect 17218 20544 17224 20596
rect 17276 20584 17282 20596
rect 17313 20587 17371 20593
rect 17313 20584 17325 20587
rect 17276 20556 17325 20584
rect 17276 20544 17282 20556
rect 17313 20553 17325 20556
rect 17359 20553 17371 20587
rect 17313 20547 17371 20553
rect 14274 20476 14280 20528
rect 14332 20516 14338 20528
rect 14332 20488 14872 20516
rect 14332 20476 14338 20488
rect 14185 20451 14243 20457
rect 14185 20417 14197 20451
rect 14231 20448 14243 20451
rect 14550 20448 14556 20460
rect 14231 20420 14556 20448
rect 14231 20417 14243 20420
rect 14185 20411 14243 20417
rect 14550 20408 14556 20420
rect 14608 20448 14614 20460
rect 14608 20420 14780 20448
rect 14608 20408 14614 20420
rect 12069 20383 12127 20389
rect 12069 20380 12081 20383
rect 11940 20352 12081 20380
rect 11940 20340 11946 20352
rect 12069 20349 12081 20352
rect 12115 20349 12127 20383
rect 12069 20343 12127 20349
rect 12253 20383 12311 20389
rect 12253 20349 12265 20383
rect 12299 20349 12311 20383
rect 12253 20343 12311 20349
rect 12621 20383 12679 20389
rect 12621 20349 12633 20383
rect 12667 20349 12679 20383
rect 12621 20343 12679 20349
rect 12897 20383 12955 20389
rect 12897 20349 12909 20383
rect 12943 20349 12955 20383
rect 14274 20380 14280 20392
rect 14235 20352 14280 20380
rect 12897 20343 12955 20349
rect 2777 20315 2835 20321
rect 2777 20281 2789 20315
rect 2823 20281 2835 20315
rect 2777 20275 2835 20281
rect 1486 20204 1492 20256
rect 1544 20244 1550 20256
rect 1581 20247 1639 20253
rect 1581 20244 1593 20247
rect 1544 20216 1593 20244
rect 1544 20204 1550 20216
rect 1581 20213 1593 20216
rect 1627 20213 1639 20247
rect 2792 20244 2820 20275
rect 3326 20272 3332 20324
rect 3384 20272 3390 20324
rect 10410 20272 10416 20324
rect 10468 20272 10474 20324
rect 11974 20272 11980 20324
rect 12032 20312 12038 20324
rect 12636 20312 12664 20343
rect 14274 20340 14280 20352
rect 14332 20340 14338 20392
rect 14752 20389 14780 20420
rect 14737 20383 14795 20389
rect 14737 20349 14749 20383
rect 14783 20349 14795 20383
rect 14844 20380 14872 20488
rect 14918 20408 14924 20460
rect 14976 20448 14982 20460
rect 15841 20451 15899 20457
rect 15841 20448 15853 20451
rect 14976 20420 15853 20448
rect 14976 20408 14982 20420
rect 15841 20417 15853 20420
rect 15887 20448 15899 20451
rect 16206 20448 16212 20460
rect 15887 20420 16212 20448
rect 15887 20417 15899 20420
rect 15841 20411 15899 20417
rect 16206 20408 16212 20420
rect 16264 20408 16270 20460
rect 19334 20448 19340 20460
rect 19295 20420 19340 20448
rect 19334 20408 19340 20420
rect 19392 20408 19398 20460
rect 15105 20383 15163 20389
rect 15105 20380 15117 20383
rect 14844 20352 15117 20380
rect 14737 20343 14795 20349
rect 15105 20349 15117 20352
rect 15151 20349 15163 20383
rect 15105 20343 15163 20349
rect 15654 20340 15660 20392
rect 15712 20380 15718 20392
rect 15933 20383 15991 20389
rect 15933 20380 15945 20383
rect 15712 20352 15945 20380
rect 15712 20340 15718 20352
rect 15933 20349 15945 20352
rect 15979 20349 15991 20383
rect 17494 20380 17500 20392
rect 17455 20352 17500 20380
rect 15933 20343 15991 20349
rect 17494 20340 17500 20352
rect 17552 20340 17558 20392
rect 19058 20380 19064 20392
rect 19019 20352 19064 20380
rect 19058 20340 19064 20352
rect 19116 20340 19122 20392
rect 14458 20312 14464 20324
rect 12032 20284 14464 20312
rect 12032 20272 12038 20284
rect 14458 20272 14464 20284
rect 14516 20272 14522 20324
rect 14918 20312 14924 20324
rect 14831 20284 14924 20312
rect 14918 20272 14924 20284
rect 14976 20272 14982 20324
rect 15013 20315 15071 20321
rect 15013 20281 15025 20315
rect 15059 20312 15071 20315
rect 15672 20312 15700 20340
rect 15059 20284 15700 20312
rect 15059 20281 15071 20284
rect 15013 20275 15071 20281
rect 20070 20272 20076 20324
rect 20128 20272 20134 20324
rect 4154 20244 4160 20256
rect 2792 20216 4160 20244
rect 1581 20207 1639 20213
rect 4154 20204 4160 20216
rect 4212 20204 4218 20256
rect 4249 20247 4307 20253
rect 4249 20213 4261 20247
rect 4295 20244 4307 20247
rect 5166 20244 5172 20256
rect 4295 20216 5172 20244
rect 4295 20213 4307 20216
rect 4249 20207 4307 20213
rect 5166 20204 5172 20216
rect 5224 20204 5230 20256
rect 5350 20244 5356 20256
rect 5311 20216 5356 20244
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 14274 20204 14280 20256
rect 14332 20244 14338 20256
rect 14936 20244 14964 20272
rect 14332 20216 14964 20244
rect 14332 20204 14338 20216
rect 15194 20204 15200 20256
rect 15252 20244 15258 20256
rect 15289 20247 15347 20253
rect 15289 20244 15301 20247
rect 15252 20216 15301 20244
rect 15252 20204 15258 20216
rect 15289 20213 15301 20216
rect 15335 20213 15347 20247
rect 15289 20207 15347 20213
rect 19610 20204 19616 20256
rect 19668 20244 19674 20256
rect 20162 20244 20168 20256
rect 19668 20216 20168 20244
rect 19668 20204 19674 20216
rect 20162 20204 20168 20216
rect 20220 20244 20226 20256
rect 20809 20247 20867 20253
rect 20809 20244 20821 20247
rect 20220 20216 20821 20244
rect 20220 20204 20226 20216
rect 20809 20213 20821 20216
rect 20855 20213 20867 20247
rect 20809 20207 20867 20213
rect 1104 20154 21804 20176
rect 1104 20102 7882 20154
rect 7934 20102 7946 20154
rect 7998 20102 8010 20154
rect 8062 20102 8074 20154
rect 8126 20102 14782 20154
rect 14834 20102 14846 20154
rect 14898 20102 14910 20154
rect 14962 20102 14974 20154
rect 15026 20102 21804 20154
rect 1104 20080 21804 20102
rect 3326 20040 3332 20052
rect 3287 20012 3332 20040
rect 3326 20000 3332 20012
rect 3384 20000 3390 20052
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 4709 20043 4767 20049
rect 4709 20040 4721 20043
rect 4212 20012 4721 20040
rect 4212 20000 4218 20012
rect 4709 20009 4721 20012
rect 4755 20009 4767 20043
rect 6181 20043 6239 20049
rect 6181 20040 6193 20043
rect 4709 20003 4767 20009
rect 4908 20012 6193 20040
rect 3145 19907 3203 19913
rect 3145 19873 3157 19907
rect 3191 19904 3203 19907
rect 4798 19904 4804 19916
rect 3191 19876 4804 19904
rect 3191 19873 3203 19876
rect 3145 19867 3203 19873
rect 4798 19864 4804 19876
rect 4856 19864 4862 19916
rect 4908 19913 4936 20012
rect 6181 20009 6193 20012
rect 6227 20009 6239 20043
rect 6181 20003 6239 20009
rect 7466 20000 7472 20052
rect 7524 20040 7530 20052
rect 8113 20043 8171 20049
rect 8113 20040 8125 20043
rect 7524 20012 8125 20040
rect 7524 20000 7530 20012
rect 8113 20009 8125 20012
rect 8159 20040 8171 20043
rect 8202 20040 8208 20052
rect 8159 20012 8208 20040
rect 8159 20009 8171 20012
rect 8113 20003 8171 20009
rect 8202 20000 8208 20012
rect 8260 20000 8266 20052
rect 10410 20000 10416 20052
rect 10468 20040 10474 20052
rect 10505 20043 10563 20049
rect 10505 20040 10517 20043
rect 10468 20012 10517 20040
rect 10468 20000 10474 20012
rect 10505 20009 10517 20012
rect 10551 20009 10563 20043
rect 16206 20040 16212 20052
rect 16167 20012 16212 20040
rect 10505 20003 10563 20009
rect 16206 20000 16212 20012
rect 16264 20000 16270 20052
rect 4985 19975 5043 19981
rect 4985 19941 4997 19975
rect 5031 19972 5043 19975
rect 5350 19972 5356 19984
rect 5031 19944 5356 19972
rect 5031 19941 5043 19944
rect 4985 19935 5043 19941
rect 5350 19932 5356 19944
rect 5408 19932 5414 19984
rect 5994 19972 6000 19984
rect 5955 19944 6000 19972
rect 5994 19932 6000 19944
rect 6052 19932 6058 19984
rect 14458 19932 14464 19984
rect 14516 19972 14522 19984
rect 15378 19972 15384 19984
rect 14516 19944 15384 19972
rect 14516 19932 14522 19944
rect 15378 19932 15384 19944
rect 15436 19972 15442 19984
rect 16393 19975 16451 19981
rect 16393 19972 16405 19975
rect 15436 19944 16405 19972
rect 15436 19932 15442 19944
rect 16393 19941 16405 19944
rect 16439 19941 16451 19975
rect 16393 19935 16451 19941
rect 4893 19907 4951 19913
rect 4893 19873 4905 19907
rect 4939 19873 4951 19907
rect 4893 19867 4951 19873
rect 5077 19907 5135 19913
rect 5077 19873 5089 19907
rect 5123 19873 5135 19907
rect 5077 19867 5135 19873
rect 4982 19796 4988 19848
rect 5040 19836 5046 19848
rect 5092 19836 5120 19867
rect 5166 19864 5172 19916
rect 5224 19913 5230 19916
rect 5224 19907 5253 19913
rect 5241 19873 5253 19907
rect 5224 19867 5253 19873
rect 5813 19907 5871 19913
rect 5813 19873 5825 19907
rect 5859 19873 5871 19907
rect 7742 19904 7748 19916
rect 7703 19876 7748 19904
rect 5813 19867 5871 19873
rect 5224 19864 5230 19867
rect 5353 19839 5411 19845
rect 5353 19836 5365 19839
rect 5040 19808 5120 19836
rect 5184 19808 5365 19836
rect 5040 19796 5046 19808
rect 5074 19728 5080 19780
rect 5132 19768 5138 19780
rect 5184 19768 5212 19808
rect 5353 19805 5365 19808
rect 5399 19805 5411 19839
rect 5353 19799 5411 19805
rect 5132 19740 5212 19768
rect 5132 19728 5138 19740
rect 5258 19728 5264 19780
rect 5316 19768 5322 19780
rect 5828 19768 5856 19867
rect 7742 19864 7748 19876
rect 7800 19864 7806 19916
rect 7929 19907 7987 19913
rect 7929 19873 7941 19907
rect 7975 19873 7987 19907
rect 10318 19904 10324 19916
rect 10231 19876 10324 19904
rect 7929 19867 7987 19873
rect 7466 19796 7472 19848
rect 7524 19836 7530 19848
rect 7650 19836 7656 19848
rect 7524 19808 7656 19836
rect 7524 19796 7530 19808
rect 7650 19796 7656 19808
rect 7708 19836 7714 19848
rect 7944 19836 7972 19867
rect 10318 19864 10324 19876
rect 10376 19904 10382 19916
rect 12894 19904 12900 19916
rect 10376 19876 12900 19904
rect 10376 19864 10382 19876
rect 12894 19864 12900 19876
rect 12952 19864 12958 19916
rect 14921 19907 14979 19913
rect 14921 19873 14933 19907
rect 14967 19904 14979 19907
rect 15102 19904 15108 19916
rect 14967 19876 15108 19904
rect 14967 19873 14979 19876
rect 14921 19867 14979 19873
rect 15102 19864 15108 19876
rect 15160 19864 15166 19916
rect 15746 19864 15752 19916
rect 15804 19904 15810 19916
rect 16117 19907 16175 19913
rect 16117 19904 16129 19907
rect 15804 19876 16129 19904
rect 15804 19864 15810 19876
rect 16117 19873 16129 19876
rect 16163 19873 16175 19907
rect 16117 19867 16175 19873
rect 20530 19864 20536 19916
rect 20588 19904 20594 19916
rect 20625 19907 20683 19913
rect 20625 19904 20637 19907
rect 20588 19876 20637 19904
rect 20588 19864 20594 19876
rect 20625 19873 20637 19876
rect 20671 19873 20683 19907
rect 20625 19867 20683 19873
rect 7708 19808 7972 19836
rect 15013 19839 15071 19845
rect 7708 19796 7714 19808
rect 15013 19805 15025 19839
rect 15059 19836 15071 19839
rect 15194 19836 15200 19848
rect 15059 19808 15200 19836
rect 15059 19805 15071 19808
rect 15013 19799 15071 19805
rect 15194 19796 15200 19808
rect 15252 19796 15258 19848
rect 15378 19836 15384 19848
rect 15339 19808 15384 19836
rect 15378 19796 15384 19808
rect 15436 19796 15442 19848
rect 5316 19740 5856 19768
rect 16393 19771 16451 19777
rect 5316 19728 5322 19740
rect 16393 19737 16405 19771
rect 16439 19768 16451 19771
rect 16482 19768 16488 19780
rect 16439 19740 16488 19768
rect 16439 19737 16451 19740
rect 16393 19731 16451 19737
rect 16482 19728 16488 19740
rect 16540 19728 16546 19780
rect 14642 19660 14648 19712
rect 14700 19700 14706 19712
rect 14737 19703 14795 19709
rect 14737 19700 14749 19703
rect 14700 19672 14749 19700
rect 14700 19660 14706 19672
rect 14737 19669 14749 19672
rect 14783 19669 14795 19703
rect 14737 19663 14795 19669
rect 20346 19660 20352 19712
rect 20404 19700 20410 19712
rect 20441 19703 20499 19709
rect 20441 19700 20453 19703
rect 20404 19672 20453 19700
rect 20404 19660 20410 19672
rect 20441 19669 20453 19672
rect 20487 19669 20499 19703
rect 20441 19663 20499 19669
rect 1104 19610 21804 19632
rect 1104 19558 4432 19610
rect 4484 19558 4496 19610
rect 4548 19558 4560 19610
rect 4612 19558 4624 19610
rect 4676 19558 11332 19610
rect 11384 19558 11396 19610
rect 11448 19558 11460 19610
rect 11512 19558 11524 19610
rect 11576 19558 18232 19610
rect 18284 19558 18296 19610
rect 18348 19558 18360 19610
rect 18412 19558 18424 19610
rect 18476 19558 21804 19610
rect 1104 19536 21804 19558
rect 5169 19499 5227 19505
rect 5169 19465 5181 19499
rect 5215 19496 5227 19499
rect 5258 19496 5264 19508
rect 5215 19468 5264 19496
rect 5215 19465 5227 19468
rect 5169 19459 5227 19465
rect 5258 19456 5264 19468
rect 5316 19456 5322 19508
rect 15378 19456 15384 19508
rect 15436 19496 15442 19508
rect 15749 19499 15807 19505
rect 15749 19496 15761 19499
rect 15436 19468 15761 19496
rect 15436 19456 15442 19468
rect 15749 19465 15761 19468
rect 15795 19465 15807 19499
rect 21082 19496 21088 19508
rect 21043 19468 21088 19496
rect 15749 19459 15807 19465
rect 21082 19456 21088 19468
rect 21140 19456 21146 19508
rect 5629 19363 5687 19369
rect 5629 19329 5641 19363
rect 5675 19360 5687 19363
rect 14642 19360 14648 19372
rect 5675 19332 5856 19360
rect 5675 19329 5687 19332
rect 5629 19323 5687 19329
rect 4525 19295 4583 19301
rect 4525 19261 4537 19295
rect 4571 19292 4583 19295
rect 5166 19292 5172 19304
rect 4571 19264 5172 19292
rect 4571 19261 4583 19264
rect 4525 19255 4583 19261
rect 5166 19252 5172 19264
rect 5224 19292 5230 19304
rect 5353 19295 5411 19301
rect 5353 19292 5365 19295
rect 5224 19264 5365 19292
rect 5224 19252 5230 19264
rect 5353 19261 5365 19264
rect 5399 19261 5411 19295
rect 5353 19255 5411 19261
rect 5445 19295 5503 19301
rect 5445 19261 5457 19295
rect 5491 19292 5503 19295
rect 5534 19292 5540 19304
rect 5491 19264 5540 19292
rect 5491 19261 5503 19264
rect 5445 19255 5503 19261
rect 5534 19252 5540 19264
rect 5592 19252 5598 19304
rect 5721 19295 5779 19301
rect 5721 19261 5733 19295
rect 5767 19261 5779 19295
rect 5828 19292 5856 19332
rect 14200 19332 14648 19360
rect 5902 19292 5908 19304
rect 5828 19264 5908 19292
rect 5721 19255 5779 19261
rect 4617 19227 4675 19233
rect 4617 19193 4629 19227
rect 4663 19224 4675 19227
rect 5626 19224 5632 19236
rect 4663 19196 5632 19224
rect 4663 19193 4675 19196
rect 4617 19187 4675 19193
rect 5626 19184 5632 19196
rect 5684 19224 5690 19236
rect 5736 19224 5764 19255
rect 5902 19252 5908 19264
rect 5960 19252 5966 19304
rect 7374 19292 7380 19304
rect 7335 19264 7380 19292
rect 7374 19252 7380 19264
rect 7432 19252 7438 19304
rect 7745 19295 7803 19301
rect 7745 19292 7757 19295
rect 7484 19264 7757 19292
rect 5684 19196 5764 19224
rect 5684 19184 5690 19196
rect 6638 19184 6644 19236
rect 6696 19224 6702 19236
rect 7484 19224 7512 19264
rect 7745 19261 7757 19264
rect 7791 19261 7803 19295
rect 8478 19292 8484 19304
rect 8439 19264 8484 19292
rect 7745 19255 7803 19261
rect 8478 19252 8484 19264
rect 8536 19252 8542 19304
rect 8574 19295 8632 19301
rect 8574 19261 8586 19295
rect 8620 19261 8632 19295
rect 8574 19255 8632 19261
rect 6696 19196 7512 19224
rect 7561 19227 7619 19233
rect 6696 19184 6702 19196
rect 7561 19193 7573 19227
rect 7607 19193 7619 19227
rect 7561 19187 7619 19193
rect 7282 19116 7288 19168
rect 7340 19156 7346 19168
rect 7576 19156 7604 19187
rect 7650 19184 7656 19236
rect 7708 19224 7714 19236
rect 7708 19196 7753 19224
rect 7708 19184 7714 19196
rect 7340 19128 7604 19156
rect 7340 19116 7346 19128
rect 7742 19116 7748 19168
rect 7800 19156 7806 19168
rect 7929 19159 7987 19165
rect 7929 19156 7941 19159
rect 7800 19128 7941 19156
rect 7800 19116 7806 19128
rect 7929 19125 7941 19128
rect 7975 19125 7987 19159
rect 8588 19156 8616 19255
rect 8938 19252 8944 19304
rect 8996 19301 9002 19304
rect 8996 19292 9004 19301
rect 9585 19295 9643 19301
rect 9585 19292 9597 19295
rect 8996 19264 9597 19292
rect 8996 19255 9004 19264
rect 9585 19261 9597 19264
rect 9631 19261 9643 19295
rect 9585 19255 9643 19261
rect 12713 19295 12771 19301
rect 12713 19261 12725 19295
rect 12759 19261 12771 19295
rect 12713 19255 12771 19261
rect 13541 19295 13599 19301
rect 13541 19261 13553 19295
rect 13587 19292 13599 19295
rect 13630 19292 13636 19304
rect 13587 19264 13636 19292
rect 13587 19261 13599 19264
rect 13541 19255 13599 19261
rect 8996 19252 9002 19255
rect 8754 19224 8760 19236
rect 8715 19196 8760 19224
rect 8754 19184 8760 19196
rect 8812 19184 8818 19236
rect 8846 19184 8852 19236
rect 8904 19224 8910 19236
rect 9677 19227 9735 19233
rect 9677 19224 9689 19227
rect 8904 19196 8949 19224
rect 9048 19196 9689 19224
rect 8904 19184 8910 19196
rect 9048 19156 9076 19196
rect 9677 19193 9689 19196
rect 9723 19193 9735 19227
rect 12728 19224 12756 19255
rect 13630 19252 13636 19264
rect 13688 19252 13694 19304
rect 13725 19295 13783 19301
rect 13725 19261 13737 19295
rect 13771 19292 13783 19295
rect 14200 19292 14228 19332
rect 14642 19320 14648 19332
rect 14700 19320 14706 19372
rect 15396 19360 15424 19456
rect 19610 19360 19616 19372
rect 15120 19332 15424 19360
rect 19571 19332 19616 19360
rect 13771 19264 14228 19292
rect 13771 19261 13783 19264
rect 13725 19255 13783 19261
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 14386 19295 14444 19301
rect 14386 19292 14398 19295
rect 14332 19264 14398 19292
rect 14332 19252 14338 19264
rect 14386 19261 14398 19264
rect 14432 19261 14444 19295
rect 14550 19292 14556 19304
rect 14511 19264 14556 19292
rect 14386 19255 14444 19261
rect 14550 19252 14556 19264
rect 14608 19252 14614 19304
rect 14734 19292 14740 19304
rect 14695 19264 14740 19292
rect 14734 19252 14740 19264
rect 14792 19252 14798 19304
rect 14921 19295 14979 19301
rect 14921 19261 14933 19295
rect 14967 19292 14979 19295
rect 15120 19292 15148 19332
rect 19610 19320 19616 19332
rect 19668 19320 19674 19372
rect 14967 19264 15148 19292
rect 14967 19261 14979 19264
rect 14921 19255 14979 19261
rect 15194 19252 15200 19304
rect 15252 19292 15258 19304
rect 15565 19295 15623 19301
rect 15565 19292 15577 19295
rect 15252 19264 15577 19292
rect 15252 19252 15258 19264
rect 15565 19261 15577 19264
rect 15611 19261 15623 19295
rect 15565 19255 15623 19261
rect 17494 19252 17500 19304
rect 17552 19292 17558 19304
rect 17589 19295 17647 19301
rect 17589 19292 17601 19295
rect 17552 19264 17601 19292
rect 17552 19252 17558 19264
rect 17589 19261 17601 19264
rect 17635 19261 17647 19295
rect 17589 19255 17647 19261
rect 17770 19252 17776 19304
rect 17828 19292 17834 19304
rect 19058 19292 19064 19304
rect 17828 19264 19064 19292
rect 17828 19252 17834 19264
rect 19058 19252 19064 19264
rect 19116 19292 19122 19304
rect 19337 19295 19395 19301
rect 19337 19292 19349 19295
rect 19116 19264 19349 19292
rect 19116 19252 19122 19264
rect 19337 19261 19349 19264
rect 19383 19261 19395 19295
rect 19337 19255 19395 19261
rect 12802 19224 12808 19236
rect 12715 19196 12808 19224
rect 9677 19187 9735 19193
rect 12802 19184 12808 19196
rect 12860 19224 12866 19236
rect 14185 19227 14243 19233
rect 14185 19224 14197 19227
rect 12860 19196 14197 19224
rect 12860 19184 12866 19196
rect 14185 19193 14197 19196
rect 14231 19193 14243 19227
rect 14185 19187 14243 19193
rect 8588 19128 9076 19156
rect 9125 19159 9183 19165
rect 7929 19119 7987 19125
rect 9125 19125 9137 19159
rect 9171 19156 9183 19159
rect 9490 19156 9496 19168
rect 9171 19128 9496 19156
rect 9171 19125 9183 19128
rect 9125 19119 9183 19125
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 12618 19156 12624 19168
rect 12579 19128 12624 19156
rect 12618 19116 12624 19128
rect 12676 19116 12682 19168
rect 12986 19116 12992 19168
rect 13044 19156 13050 19168
rect 13541 19159 13599 19165
rect 13541 19156 13553 19159
rect 13044 19128 13553 19156
rect 13044 19116 13050 19128
rect 13541 19125 13553 19128
rect 13587 19125 13599 19159
rect 13541 19119 13599 19125
rect 13630 19116 13636 19168
rect 13688 19156 13694 19168
rect 14752 19156 14780 19252
rect 15102 19184 15108 19236
rect 15160 19224 15166 19236
rect 15381 19227 15439 19233
rect 15381 19224 15393 19227
rect 15160 19196 15393 19224
rect 15160 19184 15166 19196
rect 15381 19193 15393 19196
rect 15427 19193 15439 19227
rect 15381 19187 15439 19193
rect 20346 19184 20352 19236
rect 20404 19184 20410 19236
rect 13688 19128 14780 19156
rect 13688 19116 13694 19128
rect 17678 19116 17684 19168
rect 17736 19156 17742 19168
rect 17773 19159 17831 19165
rect 17773 19156 17785 19159
rect 17736 19128 17785 19156
rect 17736 19116 17742 19128
rect 17773 19125 17785 19128
rect 17819 19125 17831 19159
rect 17773 19119 17831 19125
rect 1104 19066 21804 19088
rect 1104 19014 7882 19066
rect 7934 19014 7946 19066
rect 7998 19014 8010 19066
rect 8062 19014 8074 19066
rect 8126 19014 14782 19066
rect 14834 19014 14846 19066
rect 14898 19014 14910 19066
rect 14962 19014 14974 19066
rect 15026 19014 21804 19066
rect 1104 18992 21804 19014
rect 5534 18912 5540 18964
rect 5592 18952 5598 18964
rect 5810 18952 5816 18964
rect 5592 18924 5816 18952
rect 5592 18912 5598 18924
rect 5810 18912 5816 18924
rect 5868 18952 5874 18964
rect 6638 18952 6644 18964
rect 5868 18924 6644 18952
rect 5868 18912 5874 18924
rect 6638 18912 6644 18924
rect 6696 18912 6702 18964
rect 8846 18912 8852 18964
rect 8904 18952 8910 18964
rect 9585 18955 9643 18961
rect 9585 18952 9597 18955
rect 8904 18924 9597 18952
rect 8904 18912 8910 18924
rect 9585 18921 9597 18924
rect 9631 18921 9643 18955
rect 20257 18955 20315 18961
rect 20257 18952 20269 18955
rect 9585 18915 9643 18921
rect 16132 18924 20269 18952
rect 7282 18844 7288 18896
rect 7340 18884 7346 18896
rect 8113 18887 8171 18893
rect 7340 18856 7880 18884
rect 7340 18844 7346 18856
rect 5626 18816 5632 18828
rect 5587 18788 5632 18816
rect 5626 18776 5632 18788
rect 5684 18776 5690 18828
rect 6549 18819 6607 18825
rect 6549 18785 6561 18819
rect 6595 18816 6607 18819
rect 6730 18816 6736 18828
rect 6595 18788 6736 18816
rect 6595 18785 6607 18788
rect 6549 18779 6607 18785
rect 5350 18748 5356 18760
rect 5311 18720 5356 18748
rect 5350 18708 5356 18720
rect 5408 18708 5414 18760
rect 5537 18751 5595 18757
rect 5537 18717 5549 18751
rect 5583 18748 5595 18751
rect 5902 18748 5908 18760
rect 5583 18720 5908 18748
rect 5583 18717 5595 18720
rect 5537 18711 5595 18717
rect 5902 18708 5908 18720
rect 5960 18748 5966 18760
rect 6564 18748 6592 18779
rect 6730 18776 6736 18788
rect 6788 18816 6794 18828
rect 7374 18816 7380 18828
rect 6788 18788 7380 18816
rect 6788 18776 6794 18788
rect 7374 18776 7380 18788
rect 7432 18776 7438 18828
rect 7852 18825 7880 18856
rect 8113 18853 8125 18887
rect 8159 18884 8171 18887
rect 8938 18884 8944 18896
rect 8159 18856 8944 18884
rect 8159 18853 8171 18856
rect 8113 18847 8171 18853
rect 8938 18844 8944 18856
rect 8996 18844 9002 18896
rect 12802 18844 12808 18896
rect 12860 18844 12866 18896
rect 12986 18884 12992 18896
rect 12947 18856 12992 18884
rect 12986 18844 12992 18856
rect 13044 18844 13050 18896
rect 16132 18884 16160 18924
rect 20257 18921 20269 18924
rect 20303 18921 20315 18955
rect 20257 18915 20315 18921
rect 13648 18856 16160 18884
rect 16209 18887 16267 18893
rect 7837 18819 7895 18825
rect 7837 18785 7849 18819
rect 7883 18816 7895 18819
rect 8662 18816 8668 18828
rect 7883 18788 8668 18816
rect 7883 18785 7895 18788
rect 7837 18779 7895 18785
rect 8662 18776 8668 18788
rect 8720 18776 8726 18828
rect 8754 18776 8760 18828
rect 8812 18816 8818 18828
rect 9493 18819 9551 18825
rect 9493 18816 9505 18819
rect 8812 18788 9505 18816
rect 8812 18776 8818 18788
rect 9493 18785 9505 18788
rect 9539 18785 9551 18819
rect 12526 18816 12532 18828
rect 12487 18788 12532 18816
rect 9493 18779 9551 18785
rect 12526 18776 12532 18788
rect 12584 18776 12590 18828
rect 12621 18819 12679 18825
rect 12621 18785 12633 18819
rect 12667 18816 12679 18819
rect 12820 18816 12848 18844
rect 12667 18788 12848 18816
rect 12897 18819 12955 18825
rect 12667 18785 12679 18788
rect 12621 18779 12679 18785
rect 12897 18785 12909 18819
rect 12943 18816 12955 18819
rect 13648 18816 13676 18856
rect 16209 18853 16221 18887
rect 16255 18884 16267 18887
rect 16945 18887 17003 18893
rect 16945 18884 16957 18887
rect 16255 18856 16957 18884
rect 16255 18853 16267 18856
rect 16209 18847 16267 18853
rect 16945 18853 16957 18856
rect 16991 18853 17003 18887
rect 16945 18847 17003 18853
rect 17678 18844 17684 18896
rect 17736 18844 17742 18896
rect 19978 18844 19984 18896
rect 20036 18884 20042 18896
rect 20036 18856 20484 18884
rect 20036 18844 20042 18856
rect 12943 18788 13676 18816
rect 12943 18785 12955 18788
rect 12897 18779 12955 18785
rect 13722 18776 13728 18828
rect 13780 18816 13786 18828
rect 15470 18816 15476 18828
rect 13780 18788 13825 18816
rect 15431 18788 15476 18816
rect 13780 18776 13786 18788
rect 15470 18776 15476 18788
rect 15528 18776 15534 18828
rect 15654 18816 15660 18828
rect 15615 18788 15660 18816
rect 15654 18776 15660 18788
rect 15712 18776 15718 18828
rect 16025 18819 16083 18825
rect 16025 18785 16037 18819
rect 16071 18816 16083 18819
rect 16482 18816 16488 18828
rect 16071 18788 16488 18816
rect 16071 18785 16083 18788
rect 16025 18779 16083 18785
rect 16482 18776 16488 18788
rect 16540 18776 16546 18828
rect 16669 18819 16727 18825
rect 16669 18785 16681 18819
rect 16715 18785 16727 18819
rect 20346 18816 20352 18828
rect 20307 18788 20352 18816
rect 16669 18779 16727 18785
rect 5960 18720 6592 18748
rect 8113 18751 8171 18757
rect 5960 18708 5966 18720
rect 8113 18717 8125 18751
rect 8159 18748 8171 18751
rect 8202 18748 8208 18760
rect 8159 18720 8208 18748
rect 8159 18717 8171 18720
rect 8113 18711 8171 18717
rect 8202 18708 8208 18720
rect 8260 18708 8266 18760
rect 12805 18751 12863 18757
rect 12805 18748 12817 18751
rect 12544 18720 12817 18748
rect 12544 18692 12572 18720
rect 12805 18717 12817 18720
rect 12851 18748 12863 18751
rect 13449 18751 13507 18757
rect 13449 18748 13461 18751
rect 12851 18720 13461 18748
rect 12851 18717 12863 18720
rect 12805 18711 12863 18717
rect 13449 18717 13461 18720
rect 13495 18717 13507 18751
rect 15746 18748 15752 18760
rect 15707 18720 15752 18748
rect 13449 18711 13507 18717
rect 15746 18708 15752 18720
rect 15804 18708 15810 18760
rect 15841 18751 15899 18757
rect 15841 18717 15853 18751
rect 15887 18748 15899 18751
rect 16574 18748 16580 18760
rect 15887 18720 16580 18748
rect 15887 18717 15899 18720
rect 15841 18711 15899 18717
rect 16574 18708 16580 18720
rect 16632 18708 16638 18760
rect 16684 18692 16712 18779
rect 20346 18776 20352 18788
rect 20404 18776 20410 18828
rect 20456 18825 20484 18856
rect 20530 18844 20536 18896
rect 20588 18884 20594 18896
rect 20588 18856 21128 18884
rect 20588 18844 20594 18856
rect 21100 18825 21128 18856
rect 20441 18819 20499 18825
rect 20441 18785 20453 18819
rect 20487 18785 20499 18819
rect 20441 18779 20499 18785
rect 20901 18819 20959 18825
rect 20901 18785 20913 18819
rect 20947 18785 20959 18819
rect 20901 18779 20959 18785
rect 21085 18819 21143 18825
rect 21085 18785 21097 18819
rect 21131 18785 21143 18819
rect 21085 18779 21143 18785
rect 16942 18708 16948 18760
rect 17000 18748 17006 18760
rect 17310 18748 17316 18760
rect 17000 18720 17316 18748
rect 17000 18708 17006 18720
rect 17310 18708 17316 18720
rect 17368 18748 17374 18760
rect 18417 18751 18475 18757
rect 18417 18748 18429 18751
rect 17368 18720 18429 18748
rect 17368 18708 17374 18720
rect 18417 18717 18429 18720
rect 18463 18717 18475 18751
rect 19981 18751 20039 18757
rect 19981 18748 19993 18751
rect 18417 18711 18475 18717
rect 19076 18720 19993 18748
rect 5445 18683 5503 18689
rect 5445 18649 5457 18683
rect 5491 18680 5503 18683
rect 5718 18680 5724 18692
rect 5491 18652 5724 18680
rect 5491 18649 5503 18652
rect 5445 18643 5503 18649
rect 5718 18640 5724 18652
rect 5776 18640 5782 18692
rect 8478 18640 8484 18692
rect 8536 18680 8542 18692
rect 9030 18680 9036 18692
rect 8536 18652 9036 18680
rect 8536 18640 8542 18652
rect 9030 18640 9036 18652
rect 9088 18680 9094 18692
rect 12345 18683 12403 18689
rect 12345 18680 12357 18683
rect 9088 18652 12357 18680
rect 9088 18640 9094 18652
rect 12345 18649 12357 18652
rect 12391 18649 12403 18683
rect 12345 18643 12403 18649
rect 12526 18640 12532 18692
rect 12584 18640 12590 18692
rect 16666 18640 16672 18692
rect 16724 18640 16730 18692
rect 19076 18624 19104 18720
rect 19981 18717 19993 18720
rect 20027 18717 20039 18751
rect 19981 18711 20039 18717
rect 19150 18640 19156 18692
rect 19208 18680 19214 18692
rect 20916 18680 20944 18779
rect 19208 18652 20944 18680
rect 19208 18640 19214 18652
rect 7374 18572 7380 18624
rect 7432 18612 7438 18624
rect 7929 18615 7987 18621
rect 7929 18612 7941 18615
rect 7432 18584 7941 18612
rect 7432 18572 7438 18584
rect 7929 18581 7941 18584
rect 7975 18612 7987 18615
rect 8570 18612 8576 18624
rect 7975 18584 8576 18612
rect 7975 18581 7987 18584
rect 7929 18575 7987 18581
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 13538 18612 13544 18624
rect 13499 18584 13544 18612
rect 13538 18572 13544 18584
rect 13596 18572 13602 18624
rect 13633 18615 13691 18621
rect 13633 18581 13645 18615
rect 13679 18612 13691 18615
rect 19058 18612 19064 18624
rect 13679 18584 19064 18612
rect 13679 18581 13691 18584
rect 13633 18575 13691 18581
rect 19058 18572 19064 18584
rect 19116 18572 19122 18624
rect 20254 18572 20260 18624
rect 20312 18612 20318 18624
rect 20993 18615 21051 18621
rect 20993 18612 21005 18615
rect 20312 18584 21005 18612
rect 20312 18572 20318 18584
rect 20993 18581 21005 18584
rect 21039 18581 21051 18615
rect 20993 18575 21051 18581
rect 1104 18522 21804 18544
rect 1104 18470 4432 18522
rect 4484 18470 4496 18522
rect 4548 18470 4560 18522
rect 4612 18470 4624 18522
rect 4676 18470 11332 18522
rect 11384 18470 11396 18522
rect 11448 18470 11460 18522
rect 11512 18470 11524 18522
rect 11576 18470 18232 18522
rect 18284 18470 18296 18522
rect 18348 18470 18360 18522
rect 18412 18470 18424 18522
rect 18476 18470 21804 18522
rect 1104 18448 21804 18470
rect 6638 18368 6644 18420
rect 6696 18408 6702 18420
rect 8941 18411 8999 18417
rect 8941 18408 8953 18411
rect 6696 18380 8953 18408
rect 6696 18368 6702 18380
rect 8941 18377 8953 18380
rect 8987 18377 8999 18411
rect 8941 18371 8999 18377
rect 15746 18368 15752 18420
rect 15804 18408 15810 18420
rect 17405 18411 17463 18417
rect 17405 18408 17417 18411
rect 15804 18380 17417 18408
rect 15804 18368 15810 18380
rect 17405 18377 17417 18380
rect 17451 18377 17463 18411
rect 19058 18408 19064 18420
rect 19019 18380 19064 18408
rect 17405 18371 17463 18377
rect 19058 18368 19064 18380
rect 19116 18368 19122 18420
rect 8864 18312 12204 18340
rect 2498 18232 2504 18284
rect 2556 18272 2562 18284
rect 4525 18275 4583 18281
rect 4525 18272 4537 18275
rect 2556 18244 4537 18272
rect 2556 18232 2562 18244
rect 4525 18241 4537 18244
rect 4571 18241 4583 18275
rect 4525 18235 4583 18241
rect 8570 18232 8576 18284
rect 8628 18272 8634 18284
rect 8864 18272 8892 18312
rect 9490 18272 9496 18284
rect 8628 18244 8892 18272
rect 9451 18244 9496 18272
rect 8628 18232 8634 18244
rect 5445 18207 5503 18213
rect 5445 18173 5457 18207
rect 5491 18204 5503 18207
rect 5718 18204 5724 18216
rect 5491 18176 5724 18204
rect 5491 18173 5503 18176
rect 5445 18167 5503 18173
rect 5718 18164 5724 18176
rect 5776 18204 5782 18216
rect 6822 18204 6828 18216
rect 5776 18176 6828 18204
rect 5776 18164 5782 18176
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 8665 18207 8723 18213
rect 8665 18173 8677 18207
rect 8711 18173 8723 18207
rect 8665 18167 8723 18173
rect 8757 18207 8815 18213
rect 8757 18173 8769 18207
rect 8803 18204 8815 18207
rect 8864 18204 8892 18244
rect 9490 18232 9496 18244
rect 9548 18232 9554 18284
rect 12176 18281 12204 18312
rect 12986 18300 12992 18352
rect 13044 18300 13050 18352
rect 13722 18300 13728 18352
rect 13780 18340 13786 18352
rect 18509 18343 18567 18349
rect 18509 18340 18521 18343
rect 13780 18312 18521 18340
rect 13780 18300 13786 18312
rect 18509 18309 18521 18312
rect 18555 18309 18567 18343
rect 20530 18340 20536 18352
rect 18509 18303 18567 18309
rect 19444 18312 20536 18340
rect 12161 18275 12219 18281
rect 12161 18241 12173 18275
rect 12207 18241 12219 18275
rect 13004 18272 13032 18300
rect 12161 18235 12219 18241
rect 12820 18244 13032 18272
rect 8803 18176 8892 18204
rect 9033 18207 9091 18213
rect 8803 18173 8815 18176
rect 8757 18167 8815 18173
rect 9033 18173 9045 18207
rect 9079 18173 9091 18207
rect 9674 18204 9680 18216
rect 9635 18176 9680 18204
rect 9033 18167 9091 18173
rect 3234 18096 3240 18148
rect 3292 18096 3298 18148
rect 4246 18136 4252 18148
rect 4207 18108 4252 18136
rect 4246 18096 4252 18108
rect 4304 18096 4310 18148
rect 5074 18136 5080 18148
rect 4724 18108 5080 18136
rect 2777 18071 2835 18077
rect 2777 18037 2789 18071
rect 2823 18068 2835 18071
rect 4724 18068 4752 18108
rect 5074 18096 5080 18108
rect 5132 18096 5138 18148
rect 5626 18136 5632 18148
rect 5587 18108 5632 18136
rect 5626 18096 5632 18108
rect 5684 18096 5690 18148
rect 8680 18136 8708 18167
rect 8846 18136 8852 18148
rect 8680 18108 8852 18136
rect 8846 18096 8852 18108
rect 8904 18096 8910 18148
rect 9048 18136 9076 18167
rect 9674 18164 9680 18176
rect 9732 18164 9738 18216
rect 9769 18207 9827 18213
rect 9769 18173 9781 18207
rect 9815 18173 9827 18207
rect 10318 18204 10324 18216
rect 10279 18176 10324 18204
rect 9769 18167 9827 18173
rect 9784 18136 9812 18167
rect 10318 18164 10324 18176
rect 10376 18204 10382 18216
rect 10962 18204 10968 18216
rect 10376 18176 10968 18204
rect 10376 18164 10382 18176
rect 10962 18164 10968 18176
rect 11020 18164 11026 18216
rect 12618 18204 12624 18216
rect 12579 18176 12624 18204
rect 12618 18164 12624 18176
rect 12676 18164 12682 18216
rect 12820 18213 12848 18244
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 17218 18272 17224 18284
rect 16632 18244 17224 18272
rect 16632 18232 16638 18244
rect 17218 18232 17224 18244
rect 17276 18272 17282 18284
rect 19444 18281 19472 18312
rect 20530 18300 20536 18312
rect 20588 18300 20594 18352
rect 19429 18275 19487 18281
rect 17276 18244 17540 18272
rect 17276 18232 17282 18244
rect 12805 18207 12863 18213
rect 12805 18173 12817 18207
rect 12851 18173 12863 18207
rect 12986 18204 12992 18216
rect 12947 18176 12992 18204
rect 12805 18167 12863 18173
rect 12986 18164 12992 18176
rect 13044 18164 13050 18216
rect 13170 18204 13176 18216
rect 13131 18176 13176 18204
rect 13170 18164 13176 18176
rect 13228 18164 13234 18216
rect 13538 18204 13544 18216
rect 13499 18176 13544 18204
rect 13538 18164 13544 18176
rect 13596 18164 13602 18216
rect 17126 18164 17132 18216
rect 17184 18204 17190 18216
rect 17310 18204 17316 18216
rect 17184 18176 17316 18204
rect 17184 18164 17190 18176
rect 17310 18164 17316 18176
rect 17368 18164 17374 18216
rect 17512 18213 17540 18244
rect 19429 18241 19441 18275
rect 19475 18241 19487 18275
rect 19429 18235 19487 18241
rect 19521 18275 19579 18281
rect 19521 18241 19533 18275
rect 19567 18272 19579 18275
rect 19978 18272 19984 18284
rect 19567 18244 19984 18272
rect 19567 18241 19579 18244
rect 19521 18235 19579 18241
rect 19978 18232 19984 18244
rect 20036 18232 20042 18284
rect 17497 18207 17555 18213
rect 17497 18173 17509 18207
rect 17543 18173 17555 18207
rect 17497 18167 17555 18173
rect 18601 18207 18659 18213
rect 18601 18173 18613 18207
rect 18647 18173 18659 18207
rect 18601 18167 18659 18173
rect 10226 18136 10232 18148
rect 9048 18108 10232 18136
rect 10226 18096 10232 18108
rect 10284 18096 10290 18148
rect 18616 18136 18644 18167
rect 19150 18164 19156 18216
rect 19208 18204 19214 18216
rect 19245 18207 19303 18213
rect 19245 18204 19257 18207
rect 19208 18176 19257 18204
rect 19208 18164 19214 18176
rect 19245 18173 19257 18176
rect 19291 18173 19303 18207
rect 19610 18204 19616 18216
rect 19571 18176 19616 18204
rect 19245 18167 19303 18173
rect 19610 18164 19616 18176
rect 19668 18164 19674 18216
rect 19797 18207 19855 18213
rect 19797 18173 19809 18207
rect 19843 18204 19855 18207
rect 20254 18204 20260 18216
rect 19843 18176 20260 18204
rect 19843 18173 19855 18176
rect 19797 18167 19855 18173
rect 19812 18136 19840 18167
rect 20254 18164 20260 18176
rect 20312 18164 20318 18216
rect 20622 18164 20628 18216
rect 20680 18204 20686 18216
rect 21085 18207 21143 18213
rect 21085 18204 21097 18207
rect 20680 18176 21097 18204
rect 20680 18164 20686 18176
rect 21085 18173 21097 18176
rect 21131 18173 21143 18207
rect 21085 18167 21143 18173
rect 18616 18108 19840 18136
rect 2823 18040 4752 18068
rect 2823 18037 2835 18040
rect 2777 18031 2835 18037
rect 4798 18028 4804 18080
rect 4856 18068 4862 18080
rect 5261 18071 5319 18077
rect 5261 18068 5273 18071
rect 4856 18040 5273 18068
rect 4856 18028 4862 18040
rect 5261 18037 5273 18040
rect 5307 18037 5319 18071
rect 8478 18068 8484 18080
rect 8439 18040 8484 18068
rect 5261 18031 5319 18037
rect 8478 18028 8484 18040
rect 8536 18068 8542 18080
rect 8754 18068 8760 18080
rect 8536 18040 8760 18068
rect 8536 18028 8542 18040
rect 8754 18028 8760 18040
rect 8812 18028 8818 18080
rect 9493 18071 9551 18077
rect 9493 18037 9505 18071
rect 9539 18068 9551 18071
rect 9766 18068 9772 18080
rect 9539 18040 9772 18068
rect 9539 18037 9551 18040
rect 9493 18031 9551 18037
rect 9766 18028 9772 18040
rect 9824 18028 9830 18080
rect 10502 18068 10508 18080
rect 10463 18040 10508 18068
rect 10502 18028 10508 18040
rect 10560 18028 10566 18080
rect 15654 18028 15660 18080
rect 15712 18068 15718 18080
rect 17310 18068 17316 18080
rect 15712 18040 17316 18068
rect 15712 18028 15718 18040
rect 17310 18028 17316 18040
rect 17368 18028 17374 18080
rect 19610 18028 19616 18080
rect 19668 18068 19674 18080
rect 20346 18068 20352 18080
rect 19668 18040 20352 18068
rect 19668 18028 19674 18040
rect 20346 18028 20352 18040
rect 20404 18028 20410 18080
rect 20901 18071 20959 18077
rect 20901 18037 20913 18071
rect 20947 18068 20959 18071
rect 20990 18068 20996 18080
rect 20947 18040 20996 18068
rect 20947 18037 20959 18040
rect 20901 18031 20959 18037
rect 20990 18028 20996 18040
rect 21048 18028 21054 18080
rect 1104 17978 21804 18000
rect 1104 17926 7882 17978
rect 7934 17926 7946 17978
rect 7998 17926 8010 17978
rect 8062 17926 8074 17978
rect 8126 17926 14782 17978
rect 14834 17926 14846 17978
rect 14898 17926 14910 17978
rect 14962 17926 14974 17978
rect 15026 17926 21804 17978
rect 1104 17904 21804 17926
rect 3234 17824 3240 17876
rect 3292 17864 3298 17876
rect 3329 17867 3387 17873
rect 3329 17864 3341 17867
rect 3292 17836 3341 17864
rect 3292 17824 3298 17836
rect 3329 17833 3341 17836
rect 3375 17833 3387 17867
rect 3329 17827 3387 17833
rect 4246 17824 4252 17876
rect 4304 17864 4310 17876
rect 4617 17867 4675 17873
rect 4617 17864 4629 17867
rect 4304 17836 4629 17864
rect 4304 17824 4310 17836
rect 4617 17833 4629 17836
rect 4663 17833 4675 17867
rect 4617 17827 4675 17833
rect 12621 17867 12679 17873
rect 12621 17833 12633 17867
rect 12667 17864 12679 17867
rect 13170 17864 13176 17876
rect 12667 17836 13176 17864
rect 12667 17833 12679 17836
rect 12621 17827 12679 17833
rect 13170 17824 13176 17836
rect 13228 17824 13234 17876
rect 4893 17799 4951 17805
rect 4893 17765 4905 17799
rect 4939 17796 4951 17799
rect 5997 17799 6055 17805
rect 5997 17796 6009 17799
rect 4939 17768 6009 17796
rect 4939 17765 4951 17768
rect 4893 17759 4951 17765
rect 5997 17765 6009 17768
rect 6043 17796 6055 17799
rect 6086 17796 6092 17808
rect 6043 17768 6092 17796
rect 6043 17765 6055 17768
rect 5997 17759 6055 17765
rect 6086 17756 6092 17768
rect 6144 17756 6150 17808
rect 6181 17799 6239 17805
rect 6181 17765 6193 17799
rect 6227 17796 6239 17799
rect 6917 17799 6975 17805
rect 6917 17796 6929 17799
rect 6227 17768 6929 17796
rect 6227 17765 6239 17768
rect 6181 17759 6239 17765
rect 6917 17765 6929 17768
rect 6963 17796 6975 17799
rect 7098 17796 7104 17808
rect 6963 17768 7104 17796
rect 6963 17765 6975 17768
rect 6917 17759 6975 17765
rect 7098 17756 7104 17768
rect 7156 17756 7162 17808
rect 9766 17796 9772 17808
rect 9727 17768 9772 17796
rect 9766 17756 9772 17768
rect 9824 17756 9830 17808
rect 10502 17756 10508 17808
rect 10560 17756 10566 17808
rect 14642 17756 14648 17808
rect 14700 17796 14706 17808
rect 14921 17799 14979 17805
rect 14921 17796 14933 17799
rect 14700 17768 14933 17796
rect 14700 17756 14706 17768
rect 14921 17765 14933 17768
rect 14967 17765 14979 17799
rect 14921 17759 14979 17765
rect 15013 17799 15071 17805
rect 15013 17765 15025 17799
rect 15059 17796 15071 17799
rect 15194 17796 15200 17808
rect 15059 17768 15200 17796
rect 15059 17765 15071 17768
rect 15013 17759 15071 17765
rect 15194 17756 15200 17768
rect 15252 17756 15258 17808
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 3145 17731 3203 17737
rect 3145 17697 3157 17731
rect 3191 17697 3203 17731
rect 4798 17728 4804 17740
rect 4759 17700 4804 17728
rect 3145 17691 3203 17697
rect 3160 17660 3188 17691
rect 4798 17688 4804 17700
rect 4856 17688 4862 17740
rect 4982 17728 4988 17740
rect 4943 17700 4988 17728
rect 4982 17688 4988 17700
rect 5040 17688 5046 17740
rect 5074 17688 5080 17740
rect 5132 17737 5138 17740
rect 5132 17731 5161 17737
rect 5149 17728 5161 17731
rect 5534 17728 5540 17740
rect 5149 17700 5540 17728
rect 5149 17697 5161 17700
rect 5132 17691 5161 17697
rect 5132 17688 5138 17691
rect 5534 17688 5540 17700
rect 5592 17688 5598 17740
rect 6365 17731 6423 17737
rect 6365 17697 6377 17731
rect 6411 17728 6423 17731
rect 6638 17728 6644 17740
rect 6411 17700 6644 17728
rect 6411 17697 6423 17700
rect 6365 17691 6423 17697
rect 6638 17688 6644 17700
rect 6696 17688 6702 17740
rect 6822 17728 6828 17740
rect 6783 17700 6828 17728
rect 6822 17688 6828 17700
rect 6880 17688 6886 17740
rect 7742 17688 7748 17740
rect 7800 17728 7806 17740
rect 8021 17731 8079 17737
rect 8021 17728 8033 17731
rect 7800 17700 8033 17728
rect 7800 17688 7806 17700
rect 8021 17697 8033 17700
rect 8067 17697 8079 17731
rect 8021 17691 8079 17697
rect 8481 17731 8539 17737
rect 8481 17697 8493 17731
rect 8527 17728 8539 17731
rect 8570 17728 8576 17740
rect 8527 17700 8576 17728
rect 8527 17697 8539 17700
rect 8481 17691 8539 17697
rect 8570 17688 8576 17700
rect 8628 17728 8634 17740
rect 8938 17728 8944 17740
rect 8628 17700 8944 17728
rect 8628 17688 8634 17700
rect 8938 17688 8944 17700
rect 8996 17688 9002 17740
rect 9122 17688 9128 17740
rect 9180 17728 9186 17740
rect 9493 17731 9551 17737
rect 9493 17728 9505 17731
rect 9180 17700 9505 17728
rect 9180 17688 9186 17700
rect 9493 17697 9505 17700
rect 9539 17697 9551 17731
rect 9493 17691 9551 17697
rect 12158 17688 12164 17740
rect 12216 17728 12222 17740
rect 12253 17731 12311 17737
rect 12253 17728 12265 17731
rect 12216 17700 12265 17728
rect 12216 17688 12222 17700
rect 12253 17697 12265 17700
rect 12299 17697 12311 17731
rect 12253 17691 12311 17697
rect 12618 17688 12624 17740
rect 12676 17728 12682 17740
rect 13081 17731 13139 17737
rect 13081 17728 13093 17731
rect 12676 17700 13093 17728
rect 12676 17688 12682 17700
rect 13081 17697 13093 17700
rect 13127 17697 13139 17731
rect 13081 17691 13139 17697
rect 14458 17688 14464 17740
rect 14516 17728 14522 17740
rect 14737 17731 14795 17737
rect 14737 17728 14749 17731
rect 14516 17700 14749 17728
rect 14516 17688 14522 17700
rect 14737 17697 14749 17700
rect 14783 17697 14795 17731
rect 14737 17691 14795 17697
rect 15105 17731 15163 17737
rect 15105 17697 15117 17731
rect 15151 17728 15163 17731
rect 15470 17728 15476 17740
rect 15151 17700 15476 17728
rect 15151 17697 15163 17700
rect 15105 17691 15163 17697
rect 15470 17688 15476 17700
rect 15528 17688 15534 17740
rect 20898 17728 20904 17740
rect 20859 17700 20904 17728
rect 20898 17688 20904 17700
rect 20956 17688 20962 17740
rect 4890 17660 4896 17672
rect 3160 17632 4896 17660
rect 4890 17620 4896 17632
rect 4948 17620 4954 17672
rect 5258 17660 5264 17672
rect 5219 17632 5264 17660
rect 5258 17620 5264 17632
rect 5316 17620 5322 17672
rect 7466 17620 7472 17672
rect 7524 17660 7530 17672
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 7524 17632 8217 17660
rect 7524 17620 7530 17632
rect 8205 17629 8217 17632
rect 8251 17629 8263 17663
rect 8205 17623 8263 17629
rect 8297 17663 8355 17669
rect 8297 17629 8309 17663
rect 8343 17660 8355 17663
rect 8386 17660 8392 17672
rect 8343 17632 8392 17660
rect 8343 17629 8355 17632
rect 8297 17623 8355 17629
rect 8386 17620 8392 17632
rect 8444 17620 8450 17672
rect 12345 17663 12403 17669
rect 12345 17629 12357 17663
rect 12391 17660 12403 17663
rect 12434 17660 12440 17672
rect 12391 17632 12440 17660
rect 12391 17629 12403 17632
rect 12345 17623 12403 17629
rect 12434 17620 12440 17632
rect 12492 17620 12498 17672
rect 8113 17595 8171 17601
rect 8113 17561 8125 17595
rect 8159 17592 8171 17595
rect 8478 17592 8484 17604
rect 8159 17564 8484 17592
rect 8159 17561 8171 17564
rect 8113 17555 8171 17561
rect 8478 17552 8484 17564
rect 8536 17552 8542 17604
rect 12802 17592 12808 17604
rect 12452 17564 12808 17592
rect 1578 17524 1584 17536
rect 1539 17496 1584 17524
rect 1578 17484 1584 17496
rect 1636 17484 1642 17536
rect 7837 17527 7895 17533
rect 7837 17493 7849 17527
rect 7883 17524 7895 17527
rect 8294 17524 8300 17536
rect 7883 17496 8300 17524
rect 7883 17493 7895 17496
rect 7837 17487 7895 17493
rect 8294 17484 8300 17496
rect 8352 17484 8358 17536
rect 8846 17484 8852 17536
rect 8904 17524 8910 17536
rect 10134 17524 10140 17536
rect 8904 17496 10140 17524
rect 8904 17484 8910 17496
rect 10134 17484 10140 17496
rect 10192 17524 10198 17536
rect 12452 17533 12480 17564
rect 12802 17552 12808 17564
rect 12860 17592 12866 17604
rect 13173 17595 13231 17601
rect 13173 17592 13185 17595
rect 12860 17564 13185 17592
rect 12860 17552 12866 17564
rect 13173 17561 13185 17564
rect 13219 17561 13231 17595
rect 13173 17555 13231 17561
rect 11241 17527 11299 17533
rect 11241 17524 11253 17527
rect 10192 17496 11253 17524
rect 10192 17484 10198 17496
rect 11241 17493 11253 17496
rect 11287 17493 11299 17527
rect 11241 17487 11299 17493
rect 12437 17527 12495 17533
rect 12437 17493 12449 17527
rect 12483 17493 12495 17527
rect 12437 17487 12495 17493
rect 15289 17527 15347 17533
rect 15289 17493 15301 17527
rect 15335 17524 15347 17527
rect 15930 17524 15936 17536
rect 15335 17496 15936 17524
rect 15335 17493 15347 17496
rect 15289 17487 15347 17493
rect 15930 17484 15936 17496
rect 15988 17484 15994 17536
rect 20714 17524 20720 17536
rect 20675 17496 20720 17524
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 1104 17434 21804 17456
rect 1104 17382 4432 17434
rect 4484 17382 4496 17434
rect 4548 17382 4560 17434
rect 4612 17382 4624 17434
rect 4676 17382 11332 17434
rect 11384 17382 11396 17434
rect 11448 17382 11460 17434
rect 11512 17382 11524 17434
rect 11576 17382 18232 17434
rect 18284 17382 18296 17434
rect 18348 17382 18360 17434
rect 18412 17382 18424 17434
rect 18476 17382 21804 17434
rect 1104 17360 21804 17382
rect 5810 17280 5816 17332
rect 5868 17280 5874 17332
rect 7466 17320 7472 17332
rect 7427 17292 7472 17320
rect 7466 17280 7472 17292
rect 7524 17280 7530 17332
rect 10226 17320 10232 17332
rect 10187 17292 10232 17320
rect 10226 17280 10232 17292
rect 10284 17280 10290 17332
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 14461 17323 14519 17329
rect 12492 17292 12940 17320
rect 12492 17280 12498 17292
rect 5828 17252 5856 17280
rect 5644 17224 5856 17252
rect 5534 17116 5540 17128
rect 5495 17088 5540 17116
rect 5534 17076 5540 17088
rect 5592 17076 5598 17128
rect 5644 17125 5672 17224
rect 5902 17212 5908 17264
rect 5960 17212 5966 17264
rect 7374 17252 7380 17264
rect 6932 17224 7380 17252
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 5920 17184 5948 17212
rect 5859 17156 6776 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 6748 17128 6776 17156
rect 5629 17119 5687 17125
rect 5629 17085 5641 17119
rect 5675 17116 5687 17119
rect 5718 17116 5724 17128
rect 5675 17088 5724 17116
rect 5675 17085 5687 17088
rect 5629 17079 5687 17085
rect 5718 17076 5724 17088
rect 5776 17076 5782 17128
rect 5905 17119 5963 17125
rect 5905 17085 5917 17119
rect 5951 17085 5963 17119
rect 5905 17079 5963 17085
rect 5810 17008 5816 17060
rect 5868 17048 5874 17060
rect 5920 17048 5948 17079
rect 6730 17076 6736 17128
rect 6788 17116 6794 17128
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6788 17088 6837 17116
rect 6788 17076 6794 17088
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6932 17116 6960 17224
rect 7374 17212 7380 17224
rect 7432 17212 7438 17264
rect 12161 17255 12219 17261
rect 12161 17221 12173 17255
rect 12207 17252 12219 17255
rect 12526 17252 12532 17264
rect 12207 17224 12532 17252
rect 12207 17221 12219 17224
rect 12161 17215 12219 17221
rect 12526 17212 12532 17224
rect 12584 17212 12590 17264
rect 7098 17184 7104 17196
rect 7059 17156 7104 17184
rect 7098 17144 7104 17156
rect 7156 17144 7162 17196
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 12250 17184 12256 17196
rect 11112 17156 12256 17184
rect 11112 17144 11118 17156
rect 12250 17144 12256 17156
rect 12308 17184 12314 17196
rect 12618 17184 12624 17196
rect 12308 17156 12434 17184
rect 12579 17156 12624 17184
rect 12308 17144 12314 17156
rect 7009 17119 7067 17125
rect 7009 17116 7021 17119
rect 6932 17088 7021 17116
rect 6825 17079 6883 17085
rect 7009 17085 7021 17088
rect 7055 17085 7067 17119
rect 7190 17116 7196 17128
rect 7151 17088 7196 17116
rect 7009 17079 7067 17085
rect 7190 17076 7196 17088
rect 7248 17076 7254 17128
rect 7285 17119 7343 17125
rect 7285 17085 7297 17119
rect 7331 17085 7343 17119
rect 7285 17079 7343 17085
rect 8297 17119 8355 17125
rect 8297 17085 8309 17119
rect 8343 17116 8355 17119
rect 8478 17116 8484 17128
rect 8343 17088 8484 17116
rect 8343 17085 8355 17088
rect 8297 17079 8355 17085
rect 5868 17020 5948 17048
rect 5868 17008 5874 17020
rect 6638 17008 6644 17060
rect 6696 17048 6702 17060
rect 7300 17048 7328 17079
rect 8478 17076 8484 17088
rect 8536 17076 8542 17128
rect 10134 17116 10140 17128
rect 10095 17088 10140 17116
rect 10134 17076 10140 17088
rect 10192 17076 10198 17128
rect 12069 17119 12127 17125
rect 12069 17085 12081 17119
rect 12115 17116 12127 17119
rect 12158 17116 12164 17128
rect 12115 17088 12164 17116
rect 12115 17085 12127 17088
rect 12069 17079 12127 17085
rect 12158 17076 12164 17088
rect 12216 17076 12222 17128
rect 12406 17116 12434 17156
rect 12618 17144 12624 17156
rect 12676 17144 12682 17196
rect 12802 17184 12808 17196
rect 12763 17156 12808 17184
rect 12802 17144 12808 17156
rect 12860 17144 12866 17196
rect 12912 17125 12940 17292
rect 14461 17289 14473 17323
rect 14507 17320 14519 17323
rect 15194 17320 15200 17332
rect 14507 17292 15200 17320
rect 14507 17289 14519 17292
rect 14461 17283 14519 17289
rect 15194 17280 15200 17292
rect 15252 17280 15258 17332
rect 15930 17184 15936 17196
rect 15891 17156 15936 17184
rect 15930 17144 15936 17156
rect 15988 17144 15994 17196
rect 16209 17187 16267 17193
rect 16209 17153 16221 17187
rect 16255 17184 16267 17187
rect 16666 17184 16672 17196
rect 16255 17156 16672 17184
rect 16255 17153 16267 17156
rect 16209 17147 16267 17153
rect 16666 17144 16672 17156
rect 16724 17184 16730 17196
rect 17034 17184 17040 17196
rect 16724 17156 17040 17184
rect 16724 17144 16730 17156
rect 17034 17144 17040 17156
rect 17092 17184 17098 17196
rect 17770 17184 17776 17196
rect 17092 17156 17776 17184
rect 17092 17144 17098 17156
rect 17770 17144 17776 17156
rect 17828 17184 17834 17196
rect 19337 17187 19395 17193
rect 19337 17184 19349 17187
rect 17828 17156 19349 17184
rect 17828 17144 17834 17156
rect 19337 17153 19349 17156
rect 19383 17153 19395 17187
rect 19337 17147 19395 17153
rect 12529 17119 12587 17125
rect 12529 17116 12541 17119
rect 12406 17088 12541 17116
rect 12529 17085 12541 17088
rect 12575 17085 12587 17119
rect 12529 17079 12587 17085
rect 12897 17119 12955 17125
rect 12897 17085 12909 17119
rect 12943 17085 12955 17119
rect 12897 17079 12955 17085
rect 20714 17076 20720 17128
rect 20772 17076 20778 17128
rect 6696 17020 7328 17048
rect 6696 17008 6702 17020
rect 10962 17008 10968 17060
rect 11020 17048 11026 17060
rect 19610 17048 19616 17060
rect 11020 17034 14766 17048
rect 11020 17020 14780 17034
rect 19571 17020 19616 17048
rect 11020 17008 11026 17020
rect 5353 16983 5411 16989
rect 5353 16949 5365 16983
rect 5399 16980 5411 16983
rect 5626 16980 5632 16992
rect 5399 16952 5632 16980
rect 5399 16949 5411 16952
rect 5353 16943 5411 16949
rect 5626 16940 5632 16952
rect 5684 16980 5690 16992
rect 6546 16980 6552 16992
rect 5684 16952 6552 16980
rect 5684 16940 5690 16952
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 8205 16983 8263 16989
rect 8205 16949 8217 16983
rect 8251 16980 8263 16983
rect 8570 16980 8576 16992
rect 8251 16952 8576 16980
rect 8251 16949 8263 16952
rect 8205 16943 8263 16949
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 14752 16980 14780 17020
rect 19610 17008 19616 17020
rect 19668 17008 19674 17060
rect 16206 16980 16212 16992
rect 14752 16952 16212 16980
rect 16206 16940 16212 16952
rect 16264 16980 16270 16992
rect 17862 16980 17868 16992
rect 16264 16952 17868 16980
rect 16264 16940 16270 16952
rect 17862 16940 17868 16952
rect 17920 16940 17926 16992
rect 20254 16940 20260 16992
rect 20312 16980 20318 16992
rect 21085 16983 21143 16989
rect 21085 16980 21097 16983
rect 20312 16952 21097 16980
rect 20312 16940 20318 16952
rect 21085 16949 21097 16952
rect 21131 16949 21143 16983
rect 21085 16943 21143 16949
rect 1104 16890 21804 16912
rect 1104 16838 7882 16890
rect 7934 16838 7946 16890
rect 7998 16838 8010 16890
rect 8062 16838 8074 16890
rect 8126 16838 14782 16890
rect 14834 16838 14846 16890
rect 14898 16838 14910 16890
rect 14962 16838 14974 16890
rect 15026 16838 21804 16890
rect 1104 16816 21804 16838
rect 6638 16776 6644 16788
rect 6599 16748 6644 16776
rect 6638 16736 6644 16748
rect 6696 16736 6702 16788
rect 12253 16779 12311 16785
rect 12253 16745 12265 16779
rect 12299 16776 12311 16779
rect 12434 16776 12440 16788
rect 12299 16748 12440 16776
rect 12299 16745 12311 16748
rect 12253 16739 12311 16745
rect 12434 16736 12440 16748
rect 12492 16736 12498 16788
rect 14458 16736 14464 16788
rect 14516 16776 14522 16788
rect 19242 16776 19248 16788
rect 14516 16748 16896 16776
rect 14516 16736 14522 16748
rect 6089 16711 6147 16717
rect 6089 16677 6101 16711
rect 6135 16708 6147 16711
rect 6914 16708 6920 16720
rect 6135 16680 6920 16708
rect 6135 16677 6147 16680
rect 6089 16671 6147 16677
rect 6914 16668 6920 16680
rect 6972 16668 6978 16720
rect 8294 16708 8300 16720
rect 8128 16680 8300 16708
rect 5810 16640 5816 16652
rect 5771 16612 5816 16640
rect 5810 16600 5816 16612
rect 5868 16600 5874 16652
rect 5902 16600 5908 16652
rect 5960 16640 5966 16652
rect 6546 16640 6552 16652
rect 5960 16612 6005 16640
rect 6507 16612 6552 16640
rect 5960 16600 5966 16612
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 8128 16649 8156 16680
rect 8294 16668 8300 16680
rect 8352 16668 8358 16720
rect 14642 16668 14648 16720
rect 14700 16708 14706 16720
rect 14700 16680 15056 16708
rect 14700 16668 14706 16680
rect 15028 16652 15056 16680
rect 8113 16643 8171 16649
rect 8113 16609 8125 16643
rect 8159 16609 8171 16643
rect 8113 16603 8171 16609
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16640 8263 16643
rect 8846 16640 8852 16652
rect 8251 16612 8852 16640
rect 8251 16609 8263 16612
rect 8205 16603 8263 16609
rect 8846 16600 8852 16612
rect 8904 16600 8910 16652
rect 12161 16643 12219 16649
rect 12161 16609 12173 16643
rect 12207 16640 12219 16643
rect 12250 16640 12256 16652
rect 12207 16612 12256 16640
rect 12207 16609 12219 16612
rect 12161 16603 12219 16609
rect 12250 16600 12256 16612
rect 12308 16600 12314 16652
rect 14918 16640 14924 16652
rect 14879 16612 14924 16640
rect 14918 16600 14924 16612
rect 14976 16600 14982 16652
rect 15010 16600 15016 16652
rect 15068 16640 15074 16652
rect 15105 16643 15163 16649
rect 15105 16640 15117 16643
rect 15068 16612 15117 16640
rect 15068 16600 15074 16612
rect 15105 16609 15117 16612
rect 15151 16609 15163 16643
rect 15105 16603 15163 16609
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 16868 16649 16896 16748
rect 16960 16748 19248 16776
rect 16960 16649 16988 16748
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 19610 16736 19616 16788
rect 19668 16776 19674 16788
rect 20533 16779 20591 16785
rect 20533 16776 20545 16779
rect 19668 16748 20545 16776
rect 19668 16736 19674 16748
rect 20533 16745 20545 16748
rect 20579 16745 20591 16779
rect 20533 16739 20591 16745
rect 17218 16708 17224 16720
rect 17179 16680 17224 16708
rect 17218 16668 17224 16680
rect 17276 16668 17282 16720
rect 18969 16711 19027 16717
rect 17420 16680 18092 16708
rect 16853 16643 16911 16649
rect 15252 16612 15297 16640
rect 15252 16600 15258 16612
rect 16853 16609 16865 16643
rect 16899 16609 16911 16643
rect 16853 16603 16911 16609
rect 16945 16643 17003 16649
rect 16945 16609 16957 16643
rect 16991 16609 17003 16643
rect 17126 16640 17132 16652
rect 17087 16612 17132 16640
rect 16945 16603 17003 16609
rect 6086 16572 6092 16584
rect 6047 16544 6092 16572
rect 6086 16532 6092 16544
rect 6144 16532 6150 16584
rect 16868 16572 16896 16603
rect 17126 16600 17132 16612
rect 17184 16600 17190 16652
rect 17310 16640 17316 16652
rect 17271 16612 17316 16640
rect 17310 16600 17316 16612
rect 17368 16600 17374 16652
rect 17420 16572 17448 16680
rect 17862 16600 17868 16652
rect 17920 16640 17926 16652
rect 17957 16643 18015 16649
rect 17957 16640 17969 16643
rect 17920 16612 17969 16640
rect 17920 16600 17926 16612
rect 17957 16609 17969 16612
rect 18003 16609 18015 16643
rect 18064 16640 18092 16680
rect 18969 16677 18981 16711
rect 19015 16708 19027 16711
rect 19518 16708 19524 16720
rect 19015 16680 19524 16708
rect 19015 16677 19027 16680
rect 18969 16671 19027 16677
rect 19518 16668 19524 16680
rect 19576 16668 19582 16720
rect 20254 16708 20260 16720
rect 19904 16680 20260 16708
rect 19061 16643 19119 16649
rect 18064 16612 19012 16640
rect 17957 16603 18015 16609
rect 16868 16544 17448 16572
rect 18984 16572 19012 16612
rect 19061 16609 19073 16643
rect 19107 16640 19119 16643
rect 19904 16640 19932 16680
rect 20254 16668 20260 16680
rect 20312 16668 20318 16720
rect 19107 16612 19932 16640
rect 19981 16643 20039 16649
rect 19107 16609 19119 16612
rect 19061 16603 19119 16609
rect 19981 16609 19993 16643
rect 20027 16609 20039 16643
rect 20162 16640 20168 16652
rect 20123 16612 20168 16640
rect 19981 16603 20039 16609
rect 19886 16572 19892 16584
rect 18984 16544 19892 16572
rect 19886 16532 19892 16544
rect 19944 16572 19950 16584
rect 19996 16572 20024 16603
rect 20162 16600 20168 16612
rect 20220 16600 20226 16652
rect 20349 16643 20407 16649
rect 20349 16640 20361 16643
rect 20272 16612 20361 16640
rect 19944 16544 20024 16572
rect 19944 16532 19950 16544
rect 20070 16532 20076 16584
rect 20128 16572 20134 16584
rect 20272 16572 20300 16612
rect 20349 16609 20361 16612
rect 20395 16609 20407 16643
rect 20349 16603 20407 16609
rect 20128 16544 20300 16572
rect 20128 16532 20134 16544
rect 20806 16532 20812 16584
rect 20864 16572 20870 16584
rect 21174 16572 21180 16584
rect 20864 16544 21180 16572
rect 20864 16532 20870 16544
rect 21174 16532 21180 16544
rect 21232 16532 21238 16584
rect 13906 16396 13912 16448
rect 13964 16436 13970 16448
rect 14737 16439 14795 16445
rect 14737 16436 14749 16439
rect 13964 16408 14749 16436
rect 13964 16396 13970 16408
rect 14737 16405 14749 16408
rect 14783 16405 14795 16439
rect 14737 16399 14795 16405
rect 17497 16439 17555 16445
rect 17497 16405 17509 16439
rect 17543 16436 17555 16439
rect 17586 16436 17592 16448
rect 17543 16408 17592 16436
rect 17543 16405 17555 16408
rect 17497 16399 17555 16405
rect 17586 16396 17592 16408
rect 17644 16396 17650 16448
rect 18046 16396 18052 16448
rect 18104 16436 18110 16448
rect 18141 16439 18199 16445
rect 18141 16436 18153 16439
rect 18104 16408 18153 16436
rect 18104 16396 18110 16408
rect 18141 16405 18153 16408
rect 18187 16405 18199 16439
rect 18141 16399 18199 16405
rect 1104 16346 21804 16368
rect 1104 16294 4432 16346
rect 4484 16294 4496 16346
rect 4548 16294 4560 16346
rect 4612 16294 4624 16346
rect 4676 16294 11332 16346
rect 11384 16294 11396 16346
rect 11448 16294 11460 16346
rect 11512 16294 11524 16346
rect 11576 16294 18232 16346
rect 18284 16294 18296 16346
rect 18348 16294 18360 16346
rect 18412 16294 18424 16346
rect 18476 16294 21804 16346
rect 1104 16272 21804 16294
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 9769 16235 9827 16241
rect 9769 16232 9781 16235
rect 9732 16204 9781 16232
rect 9732 16192 9738 16204
rect 9769 16201 9781 16204
rect 9815 16201 9827 16235
rect 12158 16232 12164 16244
rect 12119 16204 12164 16232
rect 9769 16195 9827 16201
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 14918 16232 14924 16244
rect 14476 16204 14924 16232
rect 9125 16167 9183 16173
rect 9125 16133 9137 16167
rect 9171 16164 9183 16167
rect 9171 16136 9628 16164
rect 9171 16133 9183 16136
rect 9125 16127 9183 16133
rect 6822 16096 6828 16108
rect 5920 16068 6828 16096
rect 1581 16031 1639 16037
rect 1581 15997 1593 16031
rect 1627 16028 1639 16031
rect 1946 16028 1952 16040
rect 1627 16000 1952 16028
rect 1627 15997 1639 16000
rect 1581 15991 1639 15997
rect 1946 15988 1952 16000
rect 2004 15988 2010 16040
rect 2133 16031 2191 16037
rect 2133 15997 2145 16031
rect 2179 16028 2191 16031
rect 2866 16028 2872 16040
rect 2179 16000 2872 16028
rect 2179 15997 2191 16000
rect 2133 15991 2191 15997
rect 2866 15988 2872 16000
rect 2924 15988 2930 16040
rect 5920 16037 5948 16068
rect 6822 16056 6828 16068
rect 6880 16096 6886 16108
rect 9030 16096 9036 16108
rect 6880 16068 7236 16096
rect 6880 16056 6886 16068
rect 7208 16040 7236 16068
rect 8496 16068 9036 16096
rect 5905 16031 5963 16037
rect 5905 15997 5917 16031
rect 5951 15997 5963 16031
rect 5905 15991 5963 15997
rect 6914 15988 6920 16040
rect 6972 16037 6978 16040
rect 6972 16031 7021 16037
rect 6972 15997 6975 16031
rect 7009 15997 7021 16031
rect 7190 16028 7196 16040
rect 7151 16000 7196 16028
rect 6972 15991 7021 15997
rect 6972 15988 6978 15991
rect 7190 15988 7196 16000
rect 7248 15988 7254 16040
rect 7282 15988 7288 16040
rect 7340 16037 7346 16040
rect 8496 16037 8524 16068
rect 9030 16056 9036 16068
rect 9088 16056 9094 16108
rect 9600 16105 9628 16136
rect 9585 16099 9643 16105
rect 9585 16065 9597 16099
rect 9631 16065 9643 16099
rect 9585 16059 9643 16065
rect 12805 16099 12863 16105
rect 12805 16065 12817 16099
rect 12851 16096 12863 16099
rect 12986 16096 12992 16108
rect 12851 16068 12992 16096
rect 12851 16065 12863 16068
rect 12805 16059 12863 16065
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 14476 16105 14504 16204
rect 14918 16192 14924 16204
rect 14976 16232 14982 16244
rect 15565 16235 15623 16241
rect 15565 16232 15577 16235
rect 14976 16204 15577 16232
rect 14976 16192 14982 16204
rect 15565 16201 15577 16204
rect 15611 16201 15623 16235
rect 19978 16232 19984 16244
rect 19939 16204 19984 16232
rect 15565 16195 15623 16201
rect 19978 16192 19984 16204
rect 20036 16192 20042 16244
rect 15102 16164 15108 16176
rect 15063 16136 15108 16164
rect 15102 16124 15108 16136
rect 15160 16124 15166 16176
rect 19061 16167 19119 16173
rect 19061 16133 19073 16167
rect 19107 16164 19119 16167
rect 19334 16164 19340 16176
rect 19107 16136 19340 16164
rect 19107 16133 19119 16136
rect 19061 16127 19119 16133
rect 19334 16124 19340 16136
rect 19392 16164 19398 16176
rect 20162 16164 20168 16176
rect 19392 16136 20168 16164
rect 19392 16124 19398 16136
rect 20162 16124 20168 16136
rect 20220 16124 20226 16176
rect 14461 16099 14519 16105
rect 14461 16065 14473 16099
rect 14507 16065 14519 16099
rect 15010 16096 15016 16108
rect 14461 16059 14519 16065
rect 14936 16068 15016 16096
rect 7340 16031 7379 16037
rect 7367 15997 7379 16031
rect 7340 15991 7379 15997
rect 7469 16031 7527 16037
rect 7469 15997 7481 16031
rect 7515 16028 7527 16031
rect 8481 16031 8539 16037
rect 8481 16028 8493 16031
rect 7515 16000 8493 16028
rect 7515 15997 7527 16000
rect 7469 15991 7527 15997
rect 8481 15997 8493 16000
rect 8527 15997 8539 16031
rect 8481 15991 8539 15997
rect 7340 15988 7346 15991
rect 8570 15988 8576 16040
rect 8628 16028 8634 16040
rect 8846 16028 8852 16040
rect 8628 16000 8673 16028
rect 8807 16000 8852 16028
rect 8628 15988 8634 16000
rect 8846 15988 8852 16000
rect 8904 15988 8910 16040
rect 8946 16031 9004 16037
rect 8946 15997 8958 16031
rect 8992 15997 9004 16031
rect 8946 15991 9004 15997
rect 2041 15963 2099 15969
rect 2041 15929 2053 15963
rect 2087 15960 2099 15963
rect 2682 15960 2688 15972
rect 2087 15932 2688 15960
rect 2087 15929 2099 15932
rect 2041 15923 2099 15929
rect 2682 15920 2688 15932
rect 2740 15920 2746 15972
rect 5813 15963 5871 15969
rect 5813 15929 5825 15963
rect 5859 15960 5871 15963
rect 7101 15963 7159 15969
rect 7101 15960 7113 15963
rect 5859 15932 7113 15960
rect 5859 15929 5871 15932
rect 5813 15923 5871 15929
rect 7101 15929 7113 15932
rect 7147 15929 7159 15963
rect 7101 15923 7159 15929
rect 8294 15920 8300 15972
rect 8352 15960 8358 15972
rect 8757 15963 8815 15969
rect 8757 15960 8769 15963
rect 8352 15932 8769 15960
rect 8352 15920 8358 15932
rect 8757 15929 8769 15932
rect 8803 15929 8815 15963
rect 8757 15923 8815 15929
rect 6270 15852 6276 15904
rect 6328 15892 6334 15904
rect 6825 15895 6883 15901
rect 6825 15892 6837 15895
rect 6328 15864 6837 15892
rect 6328 15852 6334 15864
rect 6825 15861 6837 15864
rect 6871 15861 6883 15895
rect 6825 15855 6883 15861
rect 8478 15852 8484 15904
rect 8536 15892 8542 15904
rect 8956 15892 8984 15991
rect 9858 15988 9864 16040
rect 9916 16028 9922 16040
rect 10962 16028 10968 16040
rect 9916 16000 9961 16028
rect 10923 16000 10968 16028
rect 9916 15988 9922 16000
rect 10962 15988 10968 16000
rect 11020 15988 11026 16040
rect 12342 16028 12348 16040
rect 12303 16000 12348 16028
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 12437 16031 12495 16037
rect 12437 15997 12449 16031
rect 12483 16028 12495 16031
rect 12526 16028 12532 16040
rect 12483 16000 12532 16028
rect 12483 15997 12495 16000
rect 12437 15991 12495 15997
rect 12526 15988 12532 16000
rect 12584 15988 12590 16040
rect 14550 16028 14556 16040
rect 14511 16000 14556 16028
rect 14550 15988 14556 16000
rect 14608 15988 14614 16040
rect 14936 16037 14964 16068
rect 15010 16056 15016 16068
rect 15068 16096 15074 16108
rect 15068 16068 15792 16096
rect 15068 16056 15074 16068
rect 14924 16031 14982 16037
rect 14924 15997 14936 16031
rect 14970 15997 14982 16031
rect 14924 15991 14982 15997
rect 15194 15988 15200 16040
rect 15252 16028 15258 16040
rect 15764 16037 15792 16068
rect 17034 16056 17040 16108
rect 17092 16096 17098 16108
rect 17313 16099 17371 16105
rect 17313 16096 17325 16099
rect 17092 16068 17325 16096
rect 17092 16056 17098 16068
rect 17313 16065 17325 16068
rect 17359 16065 17371 16099
rect 17586 16096 17592 16108
rect 17547 16068 17592 16096
rect 17313 16059 17371 16065
rect 17586 16056 17592 16068
rect 17644 16056 17650 16108
rect 19242 16056 19248 16108
rect 19300 16096 19306 16108
rect 19300 16068 20484 16096
rect 19300 16056 19306 16068
rect 15565 16031 15623 16037
rect 15565 16028 15577 16031
rect 15252 16000 15577 16028
rect 15252 15988 15258 16000
rect 15565 15997 15577 16000
rect 15611 15997 15623 16031
rect 15565 15991 15623 15997
rect 15749 16031 15807 16037
rect 15749 15997 15761 16031
rect 15795 16028 15807 16031
rect 17126 16028 17132 16040
rect 15795 16000 17132 16028
rect 15795 15997 15807 16000
rect 15749 15991 15807 15997
rect 17126 15988 17132 16000
rect 17184 15988 17190 16040
rect 19518 16028 19524 16040
rect 19479 16000 19524 16028
rect 19518 15988 19524 16000
rect 19576 15988 19582 16040
rect 19794 16028 19800 16040
rect 19755 16000 19800 16028
rect 19794 15988 19800 16000
rect 19852 15988 19858 16040
rect 20456 16037 20484 16068
rect 20441 16031 20499 16037
rect 20441 15997 20453 16031
rect 20487 15997 20499 16031
rect 20441 15991 20499 15997
rect 20625 16031 20683 16037
rect 20625 15997 20637 16031
rect 20671 15997 20683 16031
rect 20625 15991 20683 15997
rect 18046 15920 18052 15972
rect 18104 15920 18110 15972
rect 19536 15960 19564 15988
rect 20640 15960 20668 15991
rect 19536 15932 20668 15960
rect 8536 15864 8984 15892
rect 9585 15895 9643 15901
rect 8536 15852 8542 15864
rect 9585 15861 9597 15895
rect 9631 15892 9643 15895
rect 10226 15892 10232 15904
rect 9631 15864 10232 15892
rect 9631 15861 9643 15864
rect 9585 15855 9643 15861
rect 10226 15852 10232 15864
rect 10284 15852 10290 15904
rect 11149 15895 11207 15901
rect 11149 15861 11161 15895
rect 11195 15892 11207 15895
rect 11238 15892 11244 15904
rect 11195 15864 11244 15892
rect 11195 15861 11207 15864
rect 11149 15855 11207 15861
rect 11238 15852 11244 15864
rect 11296 15852 11302 15904
rect 14921 15895 14979 15901
rect 14921 15861 14933 15895
rect 14967 15892 14979 15895
rect 15194 15892 15200 15904
rect 14967 15864 15200 15892
rect 14967 15861 14979 15864
rect 14921 15855 14979 15861
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 19242 15852 19248 15904
rect 19300 15892 19306 15904
rect 19613 15895 19671 15901
rect 19613 15892 19625 15895
rect 19300 15864 19625 15892
rect 19300 15852 19306 15864
rect 19613 15861 19625 15864
rect 19659 15861 19671 15895
rect 20530 15892 20536 15904
rect 20491 15864 20536 15892
rect 19613 15855 19671 15861
rect 20530 15852 20536 15864
rect 20588 15852 20594 15904
rect 1104 15802 21804 15824
rect 1104 15750 7882 15802
rect 7934 15750 7946 15802
rect 7998 15750 8010 15802
rect 8062 15750 8074 15802
rect 8126 15750 14782 15802
rect 14834 15750 14846 15802
rect 14898 15750 14910 15802
rect 14962 15750 14974 15802
rect 15026 15750 21804 15802
rect 1104 15728 21804 15750
rect 7101 15691 7159 15697
rect 7101 15657 7113 15691
rect 7147 15688 7159 15691
rect 7282 15688 7288 15700
rect 7147 15660 7288 15688
rect 7147 15657 7159 15660
rect 7101 15651 7159 15657
rect 7282 15648 7288 15660
rect 7340 15648 7346 15700
rect 8478 15648 8484 15700
rect 8536 15688 8542 15700
rect 8573 15691 8631 15697
rect 8573 15688 8585 15691
rect 8536 15660 8585 15688
rect 8536 15648 8542 15660
rect 8573 15657 8585 15660
rect 8619 15657 8631 15691
rect 13173 15691 13231 15697
rect 13173 15688 13185 15691
rect 8573 15651 8631 15657
rect 12406 15660 13185 15688
rect 12406 15632 12434 15660
rect 13173 15657 13185 15660
rect 13219 15657 13231 15691
rect 13173 15651 13231 15657
rect 13357 15691 13415 15697
rect 13357 15657 13369 15691
rect 13403 15688 13415 15691
rect 17129 15691 17187 15697
rect 13403 15660 13768 15688
rect 13403 15657 13415 15660
rect 13357 15651 13415 15657
rect 5718 15580 5724 15632
rect 5776 15620 5782 15632
rect 7190 15620 7196 15632
rect 5776 15592 7196 15620
rect 5776 15580 5782 15592
rect 7190 15580 7196 15592
rect 7248 15620 7254 15632
rect 8938 15620 8944 15632
rect 7248 15592 8156 15620
rect 7248 15580 7254 15592
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 2593 15555 2651 15561
rect 2593 15521 2605 15555
rect 2639 15552 2651 15555
rect 3053 15555 3111 15561
rect 3053 15552 3065 15555
rect 2639 15524 3065 15552
rect 2639 15521 2651 15524
rect 2593 15515 2651 15521
rect 3053 15521 3065 15524
rect 3099 15521 3111 15555
rect 3234 15552 3240 15564
rect 3195 15524 3240 15552
rect 3053 15515 3111 15521
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15521 4491 15555
rect 4433 15515 4491 15521
rect 6549 15555 6607 15561
rect 6549 15521 6561 15555
rect 6595 15521 6607 15555
rect 6549 15515 6607 15521
rect 1946 15444 1952 15496
rect 2004 15484 2010 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 2004 15456 2053 15484
rect 2004 15444 2010 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 2041 15447 2099 15453
rect 2866 15444 2872 15496
rect 2924 15484 2930 15496
rect 4448 15484 4476 15515
rect 6270 15484 6276 15496
rect 2924 15456 4476 15484
rect 6231 15456 6276 15484
rect 2924 15444 2930 15456
rect 6270 15444 6276 15456
rect 6328 15444 6334 15496
rect 6564 15484 6592 15515
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 7009 15555 7067 15561
rect 7009 15552 7021 15555
rect 6972 15524 7021 15552
rect 6972 15512 6978 15524
rect 7009 15521 7021 15524
rect 7055 15521 7067 15555
rect 7009 15515 7067 15521
rect 7282 15512 7288 15564
rect 7340 15552 7346 15564
rect 8021 15555 8079 15561
rect 8021 15552 8033 15555
rect 7340 15524 8033 15552
rect 7340 15512 7346 15524
rect 8021 15521 8033 15524
rect 8067 15521 8079 15555
rect 8021 15515 8079 15521
rect 7466 15484 7472 15496
rect 6564 15456 7472 15484
rect 7466 15444 7472 15456
rect 7524 15444 7530 15496
rect 8128 15493 8156 15592
rect 8312 15592 8944 15620
rect 8312 15564 8340 15592
rect 8938 15580 8944 15592
rect 8996 15580 9002 15632
rect 10226 15620 10232 15632
rect 10187 15592 10232 15620
rect 10226 15580 10232 15592
rect 10284 15580 10290 15632
rect 11238 15580 11244 15632
rect 11296 15580 11302 15632
rect 12342 15620 12348 15632
rect 12303 15592 12348 15620
rect 12342 15580 12348 15592
rect 12400 15592 12434 15632
rect 12713 15623 12771 15629
rect 12400 15580 12406 15592
rect 12713 15589 12725 15623
rect 12759 15620 12771 15623
rect 12986 15620 12992 15632
rect 12759 15592 12992 15620
rect 12759 15589 12771 15592
rect 12713 15583 12771 15589
rect 12986 15580 12992 15592
rect 13044 15580 13050 15632
rect 8294 15552 8300 15564
rect 8207 15524 8300 15552
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 8389 15555 8447 15561
rect 8389 15521 8401 15555
rect 8435 15552 8447 15555
rect 9858 15552 9864 15564
rect 8435 15524 9864 15552
rect 8435 15521 8447 15524
rect 8389 15515 8447 15521
rect 9858 15512 9864 15524
rect 9916 15512 9922 15564
rect 12526 15552 12532 15564
rect 12487 15524 12532 15552
rect 12526 15512 12532 15524
rect 12584 15512 12590 15564
rect 13740 15561 13768 15660
rect 17129 15657 17141 15691
rect 17175 15657 17187 15691
rect 17129 15651 17187 15657
rect 17221 15691 17279 15697
rect 17221 15657 17233 15691
rect 17267 15688 17279 15691
rect 17310 15688 17316 15700
rect 17267 15660 17316 15688
rect 17267 15657 17279 15660
rect 17221 15651 17279 15657
rect 17144 15620 17172 15651
rect 17310 15648 17316 15660
rect 17368 15648 17374 15700
rect 20257 15691 20315 15697
rect 20257 15657 20269 15691
rect 20303 15688 20315 15691
rect 20438 15688 20444 15700
rect 20303 15660 20444 15688
rect 20303 15657 20315 15660
rect 20257 15651 20315 15657
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 17144 15592 17264 15620
rect 17236 15564 17264 15592
rect 19794 15580 19800 15632
rect 19852 15620 19858 15632
rect 19852 15592 20576 15620
rect 19852 15580 19858 15592
rect 19996 15564 20024 15592
rect 20548 15564 20576 15592
rect 13354 15555 13412 15561
rect 13354 15521 13366 15555
rect 13400 15552 13412 15555
rect 13725 15555 13783 15561
rect 13400 15524 13676 15552
rect 13400 15521 13412 15524
rect 13354 15515 13412 15521
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15453 8171 15487
rect 8113 15447 8171 15453
rect 9122 15444 9128 15496
rect 9180 15484 9186 15496
rect 9953 15487 10011 15493
rect 9953 15484 9965 15487
rect 9180 15456 9965 15484
rect 9180 15444 9186 15456
rect 9953 15453 9965 15456
rect 9999 15453 10011 15487
rect 13648 15484 13676 15524
rect 13725 15521 13737 15555
rect 13771 15552 13783 15555
rect 13906 15552 13912 15564
rect 13771 15524 13912 15552
rect 13771 15521 13783 15524
rect 13725 15515 13783 15521
rect 13906 15512 13912 15524
rect 13964 15512 13970 15564
rect 16945 15555 17003 15561
rect 16945 15521 16957 15555
rect 16991 15552 17003 15555
rect 17126 15552 17132 15564
rect 16991 15524 17132 15552
rect 16991 15521 17003 15524
rect 16945 15515 17003 15521
rect 17126 15512 17132 15524
rect 17184 15512 17190 15564
rect 17218 15512 17224 15564
rect 17276 15512 17282 15564
rect 17313 15555 17371 15561
rect 17313 15521 17325 15555
rect 17359 15552 17371 15555
rect 17678 15552 17684 15564
rect 17359 15524 17684 15552
rect 17359 15521 17371 15524
rect 17313 15515 17371 15521
rect 17678 15512 17684 15524
rect 17736 15512 17742 15564
rect 19978 15552 19984 15564
rect 19891 15524 19984 15552
rect 19978 15512 19984 15524
rect 20036 15512 20042 15564
rect 20162 15552 20168 15564
rect 20075 15524 20168 15552
rect 20162 15512 20168 15524
rect 20220 15552 20226 15564
rect 20441 15555 20499 15561
rect 20441 15552 20453 15555
rect 20220 15524 20453 15552
rect 20220 15512 20226 15524
rect 20441 15521 20453 15524
rect 20487 15521 20499 15555
rect 20441 15515 20499 15521
rect 20530 15512 20536 15564
rect 20588 15552 20594 15564
rect 20588 15524 20633 15552
rect 20588 15512 20594 15524
rect 13817 15487 13875 15493
rect 13817 15484 13829 15487
rect 13648 15456 13829 15484
rect 9953 15447 10011 15453
rect 13817 15453 13829 15456
rect 13863 15484 13875 15487
rect 14550 15484 14556 15496
rect 13863 15456 14556 15484
rect 13863 15453 13875 15456
rect 13817 15447 13875 15453
rect 14550 15444 14556 15456
rect 14608 15444 14614 15496
rect 2501 15419 2559 15425
rect 2501 15385 2513 15419
rect 2547 15416 2559 15419
rect 2682 15416 2688 15428
rect 2547 15388 2688 15416
rect 2547 15385 2559 15388
rect 2501 15379 2559 15385
rect 2682 15376 2688 15388
rect 2740 15376 2746 15428
rect 4982 15376 4988 15428
rect 5040 15416 5046 15428
rect 6457 15419 6515 15425
rect 6457 15416 6469 15419
rect 5040 15388 6469 15416
rect 5040 15376 5046 15388
rect 6457 15385 6469 15388
rect 6503 15416 6515 15419
rect 9674 15416 9680 15428
rect 6503 15388 9680 15416
rect 6503 15385 6515 15388
rect 6457 15379 6515 15385
rect 9674 15376 9680 15388
rect 9732 15376 9738 15428
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15348 1639 15351
rect 1854 15348 1860 15360
rect 1627 15320 1860 15348
rect 1627 15317 1639 15320
rect 1581 15311 1639 15317
rect 1854 15308 1860 15320
rect 1912 15308 1918 15360
rect 4246 15348 4252 15360
rect 4207 15320 4252 15348
rect 4246 15308 4252 15320
rect 4304 15308 4310 15360
rect 6362 15348 6368 15360
rect 6323 15320 6368 15348
rect 6362 15308 6368 15320
rect 6420 15308 6426 15360
rect 10410 15308 10416 15360
rect 10468 15348 10474 15360
rect 11701 15351 11759 15357
rect 11701 15348 11713 15351
rect 10468 15320 11713 15348
rect 10468 15308 10474 15320
rect 11701 15317 11713 15320
rect 11747 15317 11759 15351
rect 11701 15311 11759 15317
rect 17497 15351 17555 15357
rect 17497 15317 17509 15351
rect 17543 15348 17555 15351
rect 17770 15348 17776 15360
rect 17543 15320 17776 15348
rect 17543 15317 17555 15320
rect 17497 15311 17555 15317
rect 17770 15308 17776 15320
rect 17828 15308 17834 15360
rect 1104 15258 21804 15280
rect 1104 15206 4432 15258
rect 4484 15206 4496 15258
rect 4548 15206 4560 15258
rect 4612 15206 4624 15258
rect 4676 15206 11332 15258
rect 11384 15206 11396 15258
rect 11448 15206 11460 15258
rect 11512 15206 11524 15258
rect 11576 15206 18232 15258
rect 18284 15206 18296 15258
rect 18348 15206 18360 15258
rect 18412 15206 18424 15258
rect 18476 15206 21804 15258
rect 1104 15184 21804 15206
rect 1581 15147 1639 15153
rect 1581 15113 1593 15147
rect 1627 15144 1639 15147
rect 1946 15144 1952 15156
rect 1627 15116 1952 15144
rect 1627 15113 1639 15116
rect 1581 15107 1639 15113
rect 1946 15104 1952 15116
rect 2004 15104 2010 15156
rect 6822 15144 6828 15156
rect 6783 15116 6828 15144
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 7190 15104 7196 15156
rect 7248 15144 7254 15156
rect 7285 15147 7343 15153
rect 7285 15144 7297 15147
rect 7248 15116 7297 15144
rect 7248 15104 7254 15116
rect 7285 15113 7297 15116
rect 7331 15113 7343 15147
rect 7285 15107 7343 15113
rect 9858 15104 9864 15156
rect 9916 15144 9922 15156
rect 10689 15147 10747 15153
rect 10689 15144 10701 15147
rect 9916 15116 10701 15144
rect 9916 15104 9922 15116
rect 10689 15113 10701 15116
rect 10735 15113 10747 15147
rect 10689 15107 10747 15113
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 13081 15147 13139 15153
rect 13081 15144 13093 15147
rect 12676 15116 13093 15144
rect 12676 15104 12682 15116
rect 13081 15113 13093 15116
rect 13127 15113 13139 15147
rect 13081 15107 13139 15113
rect 18874 15104 18880 15156
rect 18932 15144 18938 15156
rect 18969 15147 19027 15153
rect 18969 15144 18981 15147
rect 18932 15116 18981 15144
rect 18932 15104 18938 15116
rect 18969 15113 18981 15116
rect 19015 15144 19027 15147
rect 19242 15144 19248 15156
rect 19015 15116 19248 15144
rect 19015 15113 19027 15116
rect 18969 15107 19027 15113
rect 19242 15104 19248 15116
rect 19300 15104 19306 15156
rect 20346 15104 20352 15156
rect 20404 15144 20410 15156
rect 20901 15147 20959 15153
rect 20901 15144 20913 15147
rect 20404 15116 20913 15144
rect 20404 15104 20410 15116
rect 20901 15113 20913 15116
rect 20947 15113 20959 15147
rect 20901 15107 20959 15113
rect 4246 15076 4252 15088
rect 4207 15048 4252 15076
rect 4246 15036 4252 15048
rect 4304 15036 4310 15088
rect 9493 15079 9551 15085
rect 9493 15076 9505 15079
rect 5644 15048 9505 15076
rect 2038 15008 2044 15020
rect 1999 14980 2044 15008
rect 2038 14968 2044 14980
rect 2096 14968 2102 15020
rect 2130 14968 2136 15020
rect 2188 15008 2194 15020
rect 3881 15011 3939 15017
rect 3881 15008 3893 15011
rect 2188 14980 2233 15008
rect 3436 14980 3893 15008
rect 2188 14968 2194 14980
rect 2866 14940 2872 14952
rect 2827 14912 2872 14940
rect 2866 14900 2872 14912
rect 2924 14900 2930 14952
rect 3436 14949 3464 14980
rect 3881 14977 3893 14980
rect 3927 15008 3939 15011
rect 5644 15008 5672 15048
rect 9493 15045 9505 15048
rect 9539 15045 9551 15079
rect 14277 15079 14335 15085
rect 14277 15076 14289 15079
rect 9493 15039 9551 15045
rect 13648 15048 14289 15076
rect 8294 15008 8300 15020
rect 3927 14980 5672 15008
rect 7116 14980 8300 15008
rect 3927 14977 3939 14980
rect 3881 14971 3939 14977
rect 3421 14943 3479 14949
rect 3421 14909 3433 14943
rect 3467 14909 3479 14943
rect 3421 14903 3479 14909
rect 4890 14900 4896 14952
rect 4948 14940 4954 14952
rect 5077 14943 5135 14949
rect 5077 14940 5089 14943
rect 4948 14912 5089 14940
rect 4948 14900 4954 14912
rect 5077 14909 5089 14912
rect 5123 14909 5135 14943
rect 5077 14903 5135 14909
rect 2961 14875 3019 14881
rect 2961 14841 2973 14875
rect 3007 14841 3019 14875
rect 5092 14872 5120 14903
rect 6822 14900 6828 14952
rect 6880 14940 6886 14952
rect 7116 14949 7144 14980
rect 8294 14968 8300 14980
rect 8352 14968 8358 15020
rect 9953 15011 10011 15017
rect 9953 14977 9965 15011
rect 9999 15008 10011 15011
rect 10226 15008 10232 15020
rect 9999 14980 10232 15008
rect 9999 14977 10011 14980
rect 9953 14971 10011 14977
rect 10226 14968 10232 14980
rect 10284 14968 10290 15020
rect 13648 15017 13676 15048
rect 14277 15045 14289 15048
rect 14323 15045 14335 15079
rect 14277 15039 14335 15045
rect 14568 15048 16068 15076
rect 13633 15011 13691 15017
rect 13633 15008 13645 15011
rect 13372 14980 13645 15008
rect 7009 14943 7067 14949
rect 7009 14940 7021 14943
rect 6880 14912 7021 14940
rect 6880 14900 6886 14912
rect 7009 14909 7021 14912
rect 7055 14909 7067 14943
rect 7009 14903 7067 14909
rect 7101 14943 7159 14949
rect 7101 14909 7113 14943
rect 7147 14909 7159 14943
rect 7101 14903 7159 14909
rect 7377 14943 7435 14949
rect 7377 14909 7389 14943
rect 7423 14940 7435 14943
rect 7466 14940 7472 14952
rect 7423 14912 7472 14940
rect 7423 14909 7435 14912
rect 7377 14903 7435 14909
rect 7466 14900 7472 14912
rect 7524 14900 7530 14952
rect 10410 14900 10416 14952
rect 10468 14940 10474 14952
rect 13372 14949 13400 14980
rect 13633 14977 13645 14980
rect 13679 14977 13691 15011
rect 13633 14971 13691 14977
rect 13725 15011 13783 15017
rect 13725 14977 13737 15011
rect 13771 15008 13783 15011
rect 14568 15008 14596 15048
rect 13771 14980 14596 15008
rect 14660 14980 15240 15008
rect 13771 14977 13783 14980
rect 13725 14971 13783 14977
rect 10597 14943 10655 14949
rect 10597 14940 10609 14943
rect 10468 14912 10609 14940
rect 10468 14900 10474 14912
rect 10597 14909 10609 14912
rect 10643 14909 10655 14943
rect 10597 14903 10655 14909
rect 13265 14943 13323 14949
rect 13265 14909 13277 14943
rect 13311 14909 13323 14943
rect 13265 14903 13323 14909
rect 13357 14943 13415 14949
rect 13357 14909 13369 14943
rect 13403 14909 13415 14943
rect 13357 14903 13415 14909
rect 7558 14872 7564 14884
rect 5092 14844 7564 14872
rect 2961 14835 3019 14841
rect 1946 14804 1952 14816
rect 1907 14776 1952 14804
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 2976 14804 3004 14835
rect 7558 14832 7564 14844
rect 7616 14832 7622 14884
rect 10045 14875 10103 14881
rect 10045 14841 10057 14875
rect 10091 14872 10103 14875
rect 12066 14872 12072 14884
rect 10091 14844 12072 14872
rect 10091 14841 10103 14844
rect 10045 14835 10103 14841
rect 12066 14832 12072 14844
rect 12124 14832 12130 14884
rect 13280 14872 13308 14903
rect 13740 14872 13768 14971
rect 14660 14952 14688 14980
rect 14553 14943 14611 14949
rect 14553 14909 14565 14943
rect 14599 14940 14611 14943
rect 14642 14940 14648 14952
rect 14599 14912 14648 14940
rect 14599 14909 14611 14912
rect 14553 14903 14611 14909
rect 14642 14900 14648 14912
rect 14700 14900 14706 14952
rect 15010 14940 15016 14952
rect 14971 14912 15016 14940
rect 15010 14900 15016 14912
rect 15068 14900 15074 14952
rect 15212 14949 15240 14980
rect 15197 14943 15255 14949
rect 15197 14909 15209 14943
rect 15243 14909 15255 14943
rect 15197 14903 15255 14909
rect 13280 14844 13768 14872
rect 14277 14875 14335 14881
rect 14277 14841 14289 14875
rect 14323 14872 14335 14875
rect 15105 14875 15163 14881
rect 15105 14872 15117 14875
rect 14323 14844 15117 14872
rect 14323 14841 14335 14844
rect 14277 14835 14335 14841
rect 15105 14841 15117 14844
rect 15151 14872 15163 14875
rect 15378 14872 15384 14884
rect 15151 14844 15384 14872
rect 15151 14841 15163 14844
rect 15105 14835 15163 14841
rect 15378 14832 15384 14844
rect 15436 14832 15442 14884
rect 16040 14816 16068 15048
rect 20254 15008 20260 15020
rect 19812 14980 20260 15008
rect 18877 14943 18935 14949
rect 18877 14909 18889 14943
rect 18923 14940 18935 14943
rect 19334 14940 19340 14952
rect 18923 14912 19340 14940
rect 18923 14909 18935 14912
rect 18877 14903 18935 14909
rect 19334 14900 19340 14912
rect 19392 14900 19398 14952
rect 19812 14949 19840 14980
rect 20254 14968 20260 14980
rect 20312 14968 20318 15020
rect 19797 14943 19855 14949
rect 19797 14909 19809 14943
rect 19843 14909 19855 14943
rect 19978 14940 19984 14952
rect 19939 14912 19984 14940
rect 19797 14903 19855 14909
rect 19978 14900 19984 14912
rect 20036 14900 20042 14952
rect 20162 14940 20168 14952
rect 20123 14912 20168 14940
rect 20162 14900 20168 14912
rect 20220 14900 20226 14952
rect 21082 14940 21088 14952
rect 21043 14912 21088 14940
rect 21082 14900 21088 14912
rect 21140 14900 21146 14952
rect 19889 14875 19947 14881
rect 19889 14841 19901 14875
rect 19935 14872 19947 14875
rect 20438 14872 20444 14884
rect 19935 14844 20444 14872
rect 19935 14841 19947 14844
rect 19889 14835 19947 14841
rect 20438 14832 20444 14844
rect 20496 14832 20502 14884
rect 3234 14804 3240 14816
rect 2976 14776 3240 14804
rect 3234 14764 3240 14776
rect 3292 14804 3298 14816
rect 4249 14807 4307 14813
rect 4249 14804 4261 14807
rect 3292 14776 4261 14804
rect 3292 14764 3298 14776
rect 4249 14773 4261 14776
rect 4295 14773 4307 14807
rect 4249 14767 4307 14773
rect 4798 14764 4804 14816
rect 4856 14804 4862 14816
rect 4893 14807 4951 14813
rect 4893 14804 4905 14807
rect 4856 14776 4905 14804
rect 4856 14764 4862 14776
rect 4893 14773 4905 14776
rect 4939 14773 4951 14807
rect 4893 14767 4951 14773
rect 9953 14807 10011 14813
rect 9953 14773 9965 14807
rect 9999 14804 10011 14807
rect 12250 14804 12256 14816
rect 9999 14776 12256 14804
rect 9999 14773 10011 14776
rect 9953 14767 10011 14773
rect 12250 14764 12256 14776
rect 12308 14764 12314 14816
rect 14461 14807 14519 14813
rect 14461 14773 14473 14807
rect 14507 14804 14519 14807
rect 15194 14804 15200 14816
rect 14507 14776 15200 14804
rect 14507 14773 14519 14776
rect 14461 14767 14519 14773
rect 15194 14764 15200 14776
rect 15252 14764 15258 14816
rect 16022 14764 16028 14816
rect 16080 14804 16086 14816
rect 19613 14807 19671 14813
rect 19613 14804 19625 14807
rect 16080 14776 19625 14804
rect 16080 14764 16086 14776
rect 19613 14773 19625 14776
rect 19659 14773 19671 14807
rect 19613 14767 19671 14773
rect 1104 14714 21804 14736
rect 1104 14662 7882 14714
rect 7934 14662 7946 14714
rect 7998 14662 8010 14714
rect 8062 14662 8074 14714
rect 8126 14662 14782 14714
rect 14834 14662 14846 14714
rect 14898 14662 14910 14714
rect 14962 14662 14974 14714
rect 15026 14662 21804 14714
rect 1104 14640 21804 14662
rect 5534 14560 5540 14612
rect 5592 14600 5598 14612
rect 6086 14600 6092 14612
rect 5592 14572 6092 14600
rect 5592 14560 5598 14572
rect 6086 14560 6092 14572
rect 6144 14600 6150 14612
rect 6144 14572 6500 14600
rect 6144 14560 6150 14572
rect 4798 14492 4804 14544
rect 4856 14492 4862 14544
rect 5813 14535 5871 14541
rect 5813 14501 5825 14535
rect 5859 14532 5871 14535
rect 6362 14532 6368 14544
rect 5859 14504 6368 14532
rect 5859 14501 5871 14504
rect 5813 14495 5871 14501
rect 6362 14492 6368 14504
rect 6420 14492 6426 14544
rect 6472 14464 6500 14572
rect 14550 14560 14556 14612
rect 14608 14600 14614 14612
rect 14737 14603 14795 14609
rect 14737 14600 14749 14603
rect 14608 14572 14749 14600
rect 14608 14560 14614 14572
rect 14737 14569 14749 14572
rect 14783 14569 14795 14603
rect 14737 14563 14795 14569
rect 14921 14603 14979 14609
rect 14921 14569 14933 14603
rect 14967 14569 14979 14603
rect 14921 14563 14979 14569
rect 8294 14532 8300 14544
rect 6748 14504 8300 14532
rect 6549 14467 6607 14473
rect 6549 14464 6561 14467
rect 6472 14436 6561 14464
rect 6549 14433 6561 14436
rect 6595 14433 6607 14467
rect 6549 14427 6607 14433
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14396 4399 14399
rect 6089 14399 6147 14405
rect 4387 14368 6040 14396
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 6012 14328 6040 14368
rect 6089 14365 6101 14399
rect 6135 14396 6147 14399
rect 6748 14396 6776 14504
rect 8294 14492 8300 14504
rect 8352 14532 8358 14544
rect 9122 14532 9128 14544
rect 8352 14504 9128 14532
rect 8352 14492 8358 14504
rect 9122 14492 9128 14504
rect 9180 14492 9186 14544
rect 12897 14535 12955 14541
rect 12897 14501 12909 14535
rect 12943 14532 12955 14535
rect 14458 14532 14464 14544
rect 12943 14504 14464 14532
rect 12943 14501 12955 14504
rect 12897 14495 12955 14501
rect 14458 14492 14464 14504
rect 14516 14492 14522 14544
rect 14936 14532 14964 14563
rect 17218 14560 17224 14612
rect 17276 14600 17282 14612
rect 18049 14603 18107 14609
rect 18049 14600 18061 14603
rect 17276 14572 18061 14600
rect 17276 14560 17282 14572
rect 18049 14569 18061 14572
rect 18095 14569 18107 14603
rect 20162 14600 20168 14612
rect 20123 14572 20168 14600
rect 18049 14563 18107 14569
rect 20162 14560 20168 14572
rect 20220 14560 20226 14612
rect 20254 14560 20260 14612
rect 20312 14600 20318 14612
rect 20349 14603 20407 14609
rect 20349 14600 20361 14603
rect 20312 14572 20361 14600
rect 20312 14560 20318 14572
rect 20349 14569 20361 14572
rect 20395 14569 20407 14603
rect 20349 14563 20407 14569
rect 14568 14504 14964 14532
rect 14568 14476 14596 14504
rect 6822 14424 6828 14476
rect 6880 14464 6886 14476
rect 7377 14467 7435 14473
rect 7377 14464 7389 14467
rect 6880 14436 7389 14464
rect 6880 14424 6886 14436
rect 7377 14433 7389 14436
rect 7423 14433 7435 14467
rect 7377 14427 7435 14433
rect 12805 14467 12863 14473
rect 12805 14433 12817 14467
rect 12851 14433 12863 14467
rect 12805 14427 12863 14433
rect 6135 14368 6776 14396
rect 6135 14365 6147 14368
rect 6089 14359 6147 14365
rect 7190 14356 7196 14408
rect 7248 14396 7254 14408
rect 8754 14396 8760 14408
rect 7248 14368 8760 14396
rect 7248 14356 7254 14368
rect 8754 14356 8760 14368
rect 8812 14356 8818 14408
rect 6822 14328 6828 14340
rect 6012 14300 6828 14328
rect 6822 14288 6828 14300
rect 6880 14288 6886 14340
rect 10318 14328 10324 14340
rect 6932 14300 10324 14328
rect 5810 14220 5816 14272
rect 5868 14260 5874 14272
rect 6638 14260 6644 14272
rect 5868 14232 6644 14260
rect 5868 14220 5874 14232
rect 6638 14220 6644 14232
rect 6696 14220 6702 14272
rect 6730 14220 6736 14272
rect 6788 14260 6794 14272
rect 6932 14260 6960 14300
rect 10318 14288 10324 14300
rect 10376 14288 10382 14340
rect 12820 14328 12848 14427
rect 14550 14424 14556 14476
rect 14608 14424 14614 14476
rect 14918 14467 14976 14473
rect 14918 14433 14930 14467
rect 14964 14464 14976 14467
rect 15194 14464 15200 14476
rect 14964 14436 15200 14464
rect 14964 14433 14976 14436
rect 14918 14427 14976 14433
rect 15194 14424 15200 14436
rect 15252 14424 15258 14476
rect 15378 14464 15384 14476
rect 15339 14436 15384 14464
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 16022 14464 16028 14476
rect 15983 14436 16028 14464
rect 16022 14424 16028 14436
rect 16080 14424 16086 14476
rect 17313 14467 17371 14473
rect 17313 14433 17325 14467
rect 17359 14433 17371 14467
rect 17313 14427 17371 14433
rect 15212 14396 15240 14424
rect 17328 14396 17356 14427
rect 18046 14424 18052 14476
rect 18104 14464 18110 14476
rect 18141 14467 18199 14473
rect 18141 14464 18153 14467
rect 18104 14436 18153 14464
rect 18104 14424 18110 14436
rect 18141 14433 18153 14436
rect 18187 14433 18199 14467
rect 18141 14427 18199 14433
rect 18969 14467 19027 14473
rect 18969 14433 18981 14467
rect 19015 14464 19027 14467
rect 20346 14467 20404 14473
rect 20346 14464 20358 14467
rect 19015 14436 20358 14464
rect 19015 14433 19027 14436
rect 18969 14427 19027 14433
rect 20346 14433 20358 14436
rect 20392 14464 20404 14467
rect 20438 14464 20444 14476
rect 20392 14436 20444 14464
rect 20392 14433 20404 14436
rect 20346 14427 20404 14433
rect 20438 14424 20444 14436
rect 20496 14464 20502 14476
rect 20809 14467 20867 14473
rect 20809 14464 20821 14467
rect 20496 14436 20821 14464
rect 20496 14424 20502 14436
rect 20809 14433 20821 14436
rect 20855 14433 20867 14467
rect 20809 14427 20867 14433
rect 15212 14368 17356 14396
rect 14274 14328 14280 14340
rect 12820 14300 14280 14328
rect 14274 14288 14280 14300
rect 14332 14328 14338 14340
rect 15470 14328 15476 14340
rect 14332 14300 15476 14328
rect 14332 14288 14338 14300
rect 15470 14288 15476 14300
rect 15528 14328 15534 14340
rect 17678 14328 17684 14340
rect 15528 14300 17684 14328
rect 15528 14288 15534 14300
rect 17678 14288 17684 14300
rect 17736 14288 17742 14340
rect 7466 14260 7472 14272
rect 6788 14232 6960 14260
rect 7427 14232 7472 14260
rect 6788 14220 6794 14232
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 15289 14263 15347 14269
rect 15289 14229 15301 14263
rect 15335 14260 15347 14263
rect 15933 14263 15991 14269
rect 15933 14260 15945 14263
rect 15335 14232 15945 14260
rect 15335 14229 15347 14232
rect 15289 14223 15347 14229
rect 15933 14229 15945 14232
rect 15979 14229 15991 14263
rect 17402 14260 17408 14272
rect 17363 14232 17408 14260
rect 15933 14223 15991 14229
rect 17402 14220 17408 14232
rect 17460 14220 17466 14272
rect 18690 14220 18696 14272
rect 18748 14260 18754 14272
rect 18877 14263 18935 14269
rect 18877 14260 18889 14263
rect 18748 14232 18889 14260
rect 18748 14220 18754 14232
rect 18877 14229 18889 14232
rect 18923 14229 18935 14263
rect 18877 14223 18935 14229
rect 20254 14220 20260 14272
rect 20312 14260 20318 14272
rect 20717 14263 20775 14269
rect 20717 14260 20729 14263
rect 20312 14232 20729 14260
rect 20312 14220 20318 14232
rect 20717 14229 20729 14232
rect 20763 14229 20775 14263
rect 20717 14223 20775 14229
rect 1104 14170 21804 14192
rect 1104 14118 4432 14170
rect 4484 14118 4496 14170
rect 4548 14118 4560 14170
rect 4612 14118 4624 14170
rect 4676 14118 11332 14170
rect 11384 14118 11396 14170
rect 11448 14118 11460 14170
rect 11512 14118 11524 14170
rect 11576 14118 18232 14170
rect 18284 14118 18296 14170
rect 18348 14118 18360 14170
rect 18412 14118 18424 14170
rect 18476 14118 21804 14170
rect 1104 14096 21804 14118
rect 1946 14016 1952 14068
rect 2004 14056 2010 14068
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 2004 14028 6837 14056
rect 2004 14016 2010 14028
rect 6825 14025 6837 14028
rect 6871 14025 6883 14059
rect 6825 14019 6883 14025
rect 8662 14016 8668 14068
rect 8720 14056 8726 14068
rect 8757 14059 8815 14065
rect 8757 14056 8769 14059
rect 8720 14028 8769 14056
rect 8720 14016 8726 14028
rect 8757 14025 8769 14028
rect 8803 14025 8815 14059
rect 9677 14059 9735 14065
rect 9677 14056 9689 14059
rect 8757 14019 8815 14025
rect 8864 14028 9689 14056
rect 2866 13948 2872 14000
rect 2924 13988 2930 14000
rect 3145 13991 3203 13997
rect 3145 13988 3157 13991
rect 2924 13960 3157 13988
rect 2924 13948 2930 13960
rect 3145 13957 3157 13960
rect 3191 13957 3203 13991
rect 3145 13951 3203 13957
rect 6638 13948 6644 14000
rect 6696 13988 6702 14000
rect 6696 13960 7420 13988
rect 6696 13948 6702 13960
rect 7282 13920 7288 13932
rect 7243 13892 7288 13920
rect 7282 13880 7288 13892
rect 7340 13880 7346 13932
rect 5534 13812 5540 13864
rect 5592 13852 5598 13864
rect 6730 13852 6736 13864
rect 5592 13824 6736 13852
rect 5592 13812 5598 13824
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 6914 13812 6920 13864
rect 6972 13852 6978 13864
rect 7009 13855 7067 13861
rect 7009 13852 7021 13855
rect 6972 13824 7021 13852
rect 6972 13812 6978 13824
rect 7009 13821 7021 13824
rect 7055 13821 7067 13855
rect 7009 13815 7067 13821
rect 7101 13855 7159 13861
rect 7101 13821 7113 13855
rect 7147 13821 7159 13855
rect 7101 13815 7159 13821
rect 3326 13784 3332 13796
rect 3287 13756 3332 13784
rect 3326 13744 3332 13756
rect 3384 13744 3390 13796
rect 7116 13784 7144 13815
rect 7190 13812 7196 13864
rect 7248 13852 7254 13864
rect 7248 13824 7293 13852
rect 7248 13812 7254 13824
rect 7392 13784 7420 13960
rect 7650 13880 7656 13932
rect 7708 13920 7714 13932
rect 8864 13920 8892 14028
rect 9677 14025 9689 14028
rect 9723 14056 9735 14059
rect 10226 14056 10232 14068
rect 9723 14028 9812 14056
rect 10187 14028 10232 14056
rect 9723 14025 9735 14028
rect 9677 14019 9735 14025
rect 9784 13988 9812 14028
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 10318 14016 10324 14068
rect 10376 14056 10382 14068
rect 20901 14059 20959 14065
rect 20901 14056 20913 14059
rect 10376 14028 20913 14056
rect 10376 14016 10382 14028
rect 20901 14025 20913 14028
rect 20947 14025 20959 14059
rect 20901 14019 20959 14025
rect 9950 13988 9956 14000
rect 9784 13960 9956 13988
rect 9950 13948 9956 13960
rect 10008 13948 10014 14000
rect 10134 13948 10140 14000
rect 10192 13948 10198 14000
rect 9674 13920 9680 13932
rect 7708 13892 8892 13920
rect 9508 13892 9680 13920
rect 7708 13880 7714 13892
rect 7466 13812 7472 13864
rect 7524 13852 7530 13864
rect 8021 13855 8079 13861
rect 8021 13852 8033 13855
rect 7524 13824 8033 13852
rect 7524 13812 7530 13824
rect 8021 13821 8033 13824
rect 8067 13821 8079 13855
rect 8021 13815 8079 13821
rect 8205 13855 8263 13861
rect 8205 13821 8217 13855
rect 8251 13852 8263 13855
rect 8570 13852 8576 13864
rect 8251 13824 8576 13852
rect 8251 13821 8263 13824
rect 8205 13815 8263 13821
rect 8570 13812 8576 13824
rect 8628 13812 8634 13864
rect 8680 13861 8708 13892
rect 9508 13861 9536 13892
rect 9674 13880 9680 13892
rect 9732 13920 9738 13932
rect 10152 13920 10180 13948
rect 9732 13892 10180 13920
rect 9732 13880 9738 13892
rect 14458 13880 14464 13932
rect 14516 13920 14522 13932
rect 17589 13923 17647 13929
rect 14516 13892 14688 13920
rect 14516 13880 14522 13892
rect 8665 13855 8723 13861
rect 8665 13821 8677 13855
rect 8711 13821 8723 13855
rect 8665 13815 8723 13821
rect 9493 13855 9551 13861
rect 9493 13821 9505 13855
rect 9539 13821 9551 13855
rect 9766 13852 9772 13864
rect 9727 13824 9772 13852
rect 9493 13815 9551 13821
rect 9766 13812 9772 13824
rect 9824 13812 9830 13864
rect 9861 13855 9919 13861
rect 9861 13821 9873 13855
rect 9907 13821 9919 13855
rect 9861 13815 9919 13821
rect 9953 13855 10011 13861
rect 9953 13821 9965 13855
rect 9999 13852 10011 13855
rect 10134 13852 10140 13864
rect 9999 13824 10140 13852
rect 9999 13821 10011 13824
rect 9953 13815 10011 13821
rect 7837 13787 7895 13793
rect 7837 13784 7849 13787
rect 7116 13756 7236 13784
rect 7392 13756 7849 13784
rect 7208 13716 7236 13756
rect 7837 13753 7849 13756
rect 7883 13753 7895 13787
rect 7837 13747 7895 13753
rect 9398 13744 9404 13796
rect 9456 13784 9462 13796
rect 9876 13784 9904 13815
rect 10134 13812 10140 13824
rect 10192 13812 10198 13864
rect 12158 13852 12164 13864
rect 12119 13824 12164 13852
rect 12158 13812 12164 13824
rect 12216 13812 12222 13864
rect 12250 13812 12256 13864
rect 12308 13852 12314 13864
rect 14274 13852 14280 13864
rect 12308 13824 12353 13852
rect 14235 13824 14280 13852
rect 12308 13812 12314 13824
rect 14274 13812 14280 13824
rect 14332 13812 14338 13864
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13852 14427 13855
rect 14550 13852 14556 13864
rect 14415 13824 14556 13852
rect 14415 13821 14427 13824
rect 14369 13815 14427 13821
rect 14550 13812 14556 13824
rect 14608 13812 14614 13864
rect 14660 13861 14688 13892
rect 17589 13889 17601 13923
rect 17635 13920 17647 13923
rect 18138 13920 18144 13932
rect 17635 13892 18144 13920
rect 17635 13889 17647 13892
rect 17589 13883 17647 13889
rect 18138 13880 18144 13892
rect 18196 13880 18202 13932
rect 18966 13920 18972 13932
rect 18927 13892 18972 13920
rect 18966 13880 18972 13892
rect 19024 13880 19030 13932
rect 20438 13920 20444 13932
rect 19076 13892 20444 13920
rect 14645 13855 14703 13861
rect 14645 13821 14657 13855
rect 14691 13821 14703 13855
rect 15194 13852 15200 13864
rect 14645 13815 14703 13821
rect 14752 13824 15200 13852
rect 9456 13756 9904 13784
rect 14461 13787 14519 13793
rect 9456 13744 9462 13756
rect 14461 13753 14473 13787
rect 14507 13784 14519 13787
rect 14752 13784 14780 13824
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 17494 13852 17500 13864
rect 17455 13824 17500 13852
rect 17494 13812 17500 13824
rect 17552 13812 17558 13864
rect 17678 13852 17684 13864
rect 17639 13824 17684 13852
rect 17678 13812 17684 13824
rect 17736 13812 17742 13864
rect 17770 13812 17776 13864
rect 17828 13852 17834 13864
rect 17828 13824 17873 13852
rect 17828 13812 17834 13824
rect 18046 13812 18052 13864
rect 18104 13852 18110 13864
rect 18690 13852 18696 13864
rect 18104 13824 18696 13852
rect 18104 13812 18110 13824
rect 18690 13812 18696 13824
rect 18748 13812 18754 13864
rect 18874 13852 18880 13864
rect 18835 13824 18880 13852
rect 18874 13812 18880 13824
rect 18932 13812 18938 13864
rect 19076 13861 19104 13892
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 19061 13855 19119 13861
rect 19061 13821 19073 13855
rect 19107 13821 19119 13855
rect 19061 13815 19119 13821
rect 19245 13855 19303 13861
rect 19245 13821 19257 13855
rect 19291 13821 19303 13855
rect 19245 13815 19303 13821
rect 14507 13756 14780 13784
rect 17696 13784 17724 13812
rect 19260 13784 19288 13815
rect 20622 13812 20628 13864
rect 20680 13852 20686 13864
rect 21085 13855 21143 13861
rect 21085 13852 21097 13855
rect 20680 13824 21097 13852
rect 20680 13812 20686 13824
rect 21085 13821 21097 13824
rect 21131 13821 21143 13855
rect 21085 13815 21143 13821
rect 20070 13784 20076 13796
rect 17696 13756 20076 13784
rect 14507 13753 14519 13756
rect 14461 13747 14519 13753
rect 20070 13744 20076 13756
rect 20128 13744 20134 13796
rect 7650 13716 7656 13728
rect 7208 13688 7656 13716
rect 7650 13676 7656 13688
rect 7708 13676 7714 13728
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 14090 13716 14096 13728
rect 12492 13688 12537 13716
rect 14051 13688 14096 13716
rect 12492 13676 12498 13688
rect 14090 13676 14096 13688
rect 14148 13676 14154 13728
rect 17310 13716 17316 13728
rect 17271 13688 17316 13716
rect 17310 13676 17316 13688
rect 17368 13676 17374 13728
rect 18509 13719 18567 13725
rect 18509 13685 18521 13719
rect 18555 13716 18567 13719
rect 18598 13716 18604 13728
rect 18555 13688 18604 13716
rect 18555 13685 18567 13688
rect 18509 13679 18567 13685
rect 18598 13676 18604 13688
rect 18656 13676 18662 13728
rect 1104 13626 21804 13648
rect 1104 13574 7882 13626
rect 7934 13574 7946 13626
rect 7998 13574 8010 13626
rect 8062 13574 8074 13626
rect 8126 13574 14782 13626
rect 14834 13574 14846 13626
rect 14898 13574 14910 13626
rect 14962 13574 14974 13626
rect 15026 13574 21804 13626
rect 1104 13552 21804 13574
rect 1578 13472 1584 13524
rect 1636 13512 1642 13524
rect 1857 13515 1915 13521
rect 1857 13512 1869 13515
rect 1636 13484 1869 13512
rect 1636 13472 1642 13484
rect 1857 13481 1869 13484
rect 1903 13481 1915 13515
rect 1857 13475 1915 13481
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 7374 13512 7380 13524
rect 7156 13484 7380 13512
rect 7156 13472 7162 13484
rect 7374 13472 7380 13484
rect 7432 13472 7438 13524
rect 8297 13515 8355 13521
rect 8297 13481 8309 13515
rect 8343 13512 8355 13515
rect 8386 13512 8392 13524
rect 8343 13484 8392 13512
rect 8343 13481 8355 13484
rect 8297 13475 8355 13481
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 18138 13512 18144 13524
rect 18099 13484 18144 13512
rect 18138 13472 18144 13484
rect 18196 13472 18202 13524
rect 6086 13444 6092 13456
rect 6047 13416 6092 13444
rect 6086 13404 6092 13416
rect 6144 13404 6150 13456
rect 6457 13447 6515 13453
rect 6457 13413 6469 13447
rect 6503 13444 6515 13447
rect 6914 13444 6920 13456
rect 6503 13416 6920 13444
rect 6503 13413 6515 13416
rect 6457 13407 6515 13413
rect 6914 13404 6920 13416
rect 6972 13444 6978 13456
rect 10042 13444 10048 13456
rect 6972 13416 10048 13444
rect 6972 13404 6978 13416
rect 1949 13379 2007 13385
rect 1949 13345 1961 13379
rect 1995 13376 2007 13379
rect 4890 13376 4896 13388
rect 1995 13348 4896 13376
rect 1995 13345 2007 13348
rect 1949 13339 2007 13345
rect 4890 13336 4896 13348
rect 4948 13336 4954 13388
rect 6273 13379 6331 13385
rect 6273 13345 6285 13379
rect 6319 13376 6331 13379
rect 6822 13376 6828 13388
rect 6319 13348 6828 13376
rect 6319 13345 6331 13348
rect 6273 13339 6331 13345
rect 6822 13336 6828 13348
rect 6880 13336 6886 13388
rect 7300 13385 7328 13416
rect 10042 13404 10048 13416
rect 10100 13444 10106 13456
rect 11241 13447 11299 13453
rect 11241 13444 11253 13447
rect 10100 13416 11253 13444
rect 10100 13404 10106 13416
rect 11241 13413 11253 13416
rect 11287 13413 11299 13447
rect 12066 13444 12072 13456
rect 12027 13416 12072 13444
rect 11241 13407 11299 13413
rect 12066 13404 12072 13416
rect 12124 13404 12130 13456
rect 12161 13447 12219 13453
rect 12161 13413 12173 13447
rect 12207 13413 12219 13447
rect 12161 13407 12219 13413
rect 12345 13447 12403 13453
rect 12345 13413 12357 13447
rect 12391 13444 12403 13447
rect 12434 13444 12440 13456
rect 12391 13416 12440 13444
rect 12391 13413 12403 13416
rect 12345 13407 12403 13413
rect 7285 13379 7343 13385
rect 7285 13345 7297 13379
rect 7331 13345 7343 13379
rect 8202 13376 8208 13388
rect 8163 13348 8208 13376
rect 7285 13339 7343 13345
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 8570 13336 8576 13388
rect 8628 13376 8634 13388
rect 9490 13376 9496 13388
rect 8628 13348 9496 13376
rect 8628 13336 8634 13348
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 9674 13376 9680 13388
rect 9635 13348 9680 13376
rect 9674 13336 9680 13348
rect 9732 13336 9738 13388
rect 10226 13336 10232 13388
rect 10284 13376 10290 13388
rect 11057 13379 11115 13385
rect 11057 13376 11069 13379
rect 10284 13348 11069 13376
rect 10284 13336 10290 13348
rect 11057 13345 11069 13348
rect 11103 13345 11115 13379
rect 11057 13339 11115 13345
rect 1765 13311 1823 13317
rect 1765 13277 1777 13311
rect 1811 13308 1823 13311
rect 2130 13308 2136 13320
rect 1811 13280 2136 13308
rect 1811 13277 1823 13280
rect 1765 13271 1823 13277
rect 2130 13268 2136 13280
rect 2188 13268 2194 13320
rect 6178 13268 6184 13320
rect 6236 13308 6242 13320
rect 12176 13308 12204 13407
rect 12434 13404 12440 13416
rect 12492 13404 12498 13456
rect 15194 13404 15200 13456
rect 15252 13444 15258 13456
rect 15657 13447 15715 13453
rect 15657 13444 15669 13447
rect 15252 13416 15669 13444
rect 15252 13404 15258 13416
rect 15657 13413 15669 13416
rect 15703 13413 15715 13447
rect 15657 13407 15715 13413
rect 17310 13404 17316 13456
rect 17368 13444 17374 13456
rect 17405 13447 17463 13453
rect 17405 13444 17417 13447
rect 17368 13416 17417 13444
rect 17368 13404 17374 13416
rect 17405 13413 17417 13416
rect 17451 13413 17463 13447
rect 17405 13407 17463 13413
rect 19886 13404 19892 13456
rect 19944 13444 19950 13456
rect 19944 13416 20576 13444
rect 19944 13404 19950 13416
rect 16390 13376 16396 13388
rect 16330 13348 16396 13376
rect 16390 13336 16396 13348
rect 16448 13336 16454 13388
rect 18046 13336 18052 13388
rect 18104 13376 18110 13388
rect 18325 13379 18383 13385
rect 18325 13376 18337 13379
rect 18104 13348 18337 13376
rect 18104 13336 18110 13348
rect 18325 13345 18337 13348
rect 18371 13345 18383 13379
rect 18325 13339 18383 13345
rect 18509 13379 18567 13385
rect 18509 13345 18521 13379
rect 18555 13345 18567 13379
rect 18509 13339 18567 13345
rect 6236 13280 12204 13308
rect 6236 13268 6242 13280
rect 13814 13268 13820 13320
rect 13872 13308 13878 13320
rect 17034 13308 17040 13320
rect 13872 13280 17040 13308
rect 13872 13268 13878 13280
rect 17034 13268 17040 13280
rect 17092 13308 17098 13320
rect 17678 13308 17684 13320
rect 17092 13280 17684 13308
rect 17092 13268 17098 13280
rect 17678 13268 17684 13280
rect 17736 13268 17742 13320
rect 18524 13308 18552 13339
rect 20070 13336 20076 13388
rect 20128 13385 20134 13388
rect 20128 13379 20177 13385
rect 20128 13345 20131 13379
rect 20165 13345 20177 13379
rect 20254 13376 20260 13388
rect 20215 13348 20260 13376
rect 20128 13339 20177 13345
rect 20128 13336 20134 13339
rect 20254 13336 20260 13348
rect 20312 13336 20318 13388
rect 20349 13379 20407 13385
rect 20349 13345 20361 13379
rect 20395 13376 20407 13379
rect 20438 13376 20444 13388
rect 20395 13348 20444 13376
rect 20395 13345 20407 13348
rect 20349 13339 20407 13345
rect 20438 13336 20444 13348
rect 20496 13336 20502 13388
rect 20548 13385 20576 13416
rect 20533 13379 20591 13385
rect 20533 13345 20545 13379
rect 20579 13345 20591 13379
rect 20533 13339 20591 13345
rect 18248 13280 18552 13308
rect 13078 13200 13084 13252
rect 13136 13240 13142 13252
rect 16298 13240 16304 13252
rect 13136 13212 16304 13240
rect 13136 13200 13142 13212
rect 16298 13200 16304 13212
rect 16356 13200 16362 13252
rect 2130 13132 2136 13184
rect 2188 13172 2194 13184
rect 2317 13175 2375 13181
rect 2317 13172 2329 13175
rect 2188 13144 2329 13172
rect 2188 13132 2194 13144
rect 2317 13141 2329 13144
rect 2363 13141 2375 13175
rect 2317 13135 2375 13141
rect 8662 13132 8668 13184
rect 8720 13172 8726 13184
rect 9306 13172 9312 13184
rect 8720 13144 9312 13172
rect 8720 13132 8726 13144
rect 9306 13132 9312 13144
rect 9364 13172 9370 13184
rect 9493 13175 9551 13181
rect 9493 13172 9505 13175
rect 9364 13144 9505 13172
rect 9364 13132 9370 13144
rect 9493 13141 9505 13144
rect 9539 13141 9551 13175
rect 9493 13135 9551 13141
rect 9861 13175 9919 13181
rect 9861 13141 9873 13175
rect 9907 13172 9919 13175
rect 11054 13172 11060 13184
rect 9907 13144 11060 13172
rect 9907 13141 9919 13144
rect 9861 13135 9919 13141
rect 11054 13132 11060 13144
rect 11112 13132 11118 13184
rect 11425 13175 11483 13181
rect 11425 13141 11437 13175
rect 11471 13172 11483 13175
rect 11790 13172 11796 13184
rect 11471 13144 11796 13172
rect 11471 13141 11483 13144
rect 11425 13135 11483 13141
rect 11790 13132 11796 13144
rect 11848 13132 11854 13184
rect 12621 13175 12679 13181
rect 12621 13141 12633 13175
rect 12667 13172 12679 13175
rect 14182 13172 14188 13184
rect 12667 13144 14188 13172
rect 12667 13141 12679 13144
rect 12621 13135 12679 13141
rect 14182 13132 14188 13144
rect 14240 13132 14246 13184
rect 17402 13132 17408 13184
rect 17460 13172 17466 13184
rect 18248 13172 18276 13280
rect 17460 13144 18276 13172
rect 18509 13175 18567 13181
rect 17460 13132 17466 13144
rect 18509 13141 18521 13175
rect 18555 13172 18567 13175
rect 18874 13172 18880 13184
rect 18555 13144 18880 13172
rect 18555 13141 18567 13144
rect 18509 13135 18567 13141
rect 18874 13132 18880 13144
rect 18932 13132 18938 13184
rect 19610 13132 19616 13184
rect 19668 13172 19674 13184
rect 19981 13175 20039 13181
rect 19981 13172 19993 13175
rect 19668 13144 19993 13172
rect 19668 13132 19674 13144
rect 19981 13141 19993 13144
rect 20027 13141 20039 13175
rect 19981 13135 20039 13141
rect 1104 13082 21804 13104
rect 1104 13030 4432 13082
rect 4484 13030 4496 13082
rect 4548 13030 4560 13082
rect 4612 13030 4624 13082
rect 4676 13030 11332 13082
rect 11384 13030 11396 13082
rect 11448 13030 11460 13082
rect 11512 13030 11524 13082
rect 11576 13030 18232 13082
rect 18284 13030 18296 13082
rect 18348 13030 18360 13082
rect 18412 13030 18424 13082
rect 18476 13030 21804 13082
rect 1104 13008 21804 13030
rect 1486 12968 1492 12980
rect 1447 12940 1492 12968
rect 1486 12928 1492 12940
rect 1544 12928 1550 12980
rect 2685 12971 2743 12977
rect 2685 12937 2697 12971
rect 2731 12968 2743 12971
rect 3326 12968 3332 12980
rect 2731 12940 3332 12968
rect 2731 12937 2743 12940
rect 2685 12931 2743 12937
rect 3326 12928 3332 12940
rect 3384 12968 3390 12980
rect 3513 12971 3571 12977
rect 3513 12968 3525 12971
rect 3384 12940 3525 12968
rect 3384 12928 3390 12940
rect 3513 12937 3525 12940
rect 3559 12937 3571 12971
rect 4890 12968 4896 12980
rect 4851 12940 4896 12968
rect 3513 12931 3571 12937
rect 4890 12928 4896 12940
rect 4948 12928 4954 12980
rect 5261 12971 5319 12977
rect 5261 12937 5273 12971
rect 5307 12937 5319 12971
rect 5261 12931 5319 12937
rect 5276 12900 5304 12931
rect 9766 12928 9772 12980
rect 9824 12968 9830 12980
rect 9953 12971 10011 12977
rect 9953 12968 9965 12971
rect 9824 12940 9965 12968
rect 9824 12928 9830 12940
rect 9953 12937 9965 12940
rect 9999 12937 10011 12971
rect 9953 12931 10011 12937
rect 10042 12928 10048 12980
rect 10100 12968 10106 12980
rect 10318 12968 10324 12980
rect 10100 12940 10324 12968
rect 10100 12928 10106 12940
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 10965 12971 11023 12977
rect 10965 12937 10977 12971
rect 11011 12968 11023 12971
rect 11698 12968 11704 12980
rect 11011 12940 11704 12968
rect 11011 12937 11023 12940
rect 10965 12931 11023 12937
rect 11698 12928 11704 12940
rect 11756 12968 11762 12980
rect 12250 12968 12256 12980
rect 11756 12940 12256 12968
rect 11756 12928 11762 12940
rect 12250 12928 12256 12940
rect 12308 12928 12314 12980
rect 14550 12928 14556 12980
rect 14608 12968 14614 12980
rect 15565 12971 15623 12977
rect 15565 12968 15577 12971
rect 14608 12940 15577 12968
rect 14608 12928 14614 12940
rect 15565 12937 15577 12940
rect 15611 12937 15623 12971
rect 16390 12968 16396 12980
rect 16351 12940 16396 12968
rect 15565 12931 15623 12937
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 17405 12971 17463 12977
rect 17405 12937 17417 12971
rect 17451 12968 17463 12971
rect 17494 12968 17500 12980
rect 17451 12940 17500 12968
rect 17451 12937 17463 12940
rect 17405 12931 17463 12937
rect 17494 12928 17500 12940
rect 17552 12928 17558 12980
rect 20254 12928 20260 12980
rect 20312 12968 20318 12980
rect 21085 12971 21143 12977
rect 21085 12968 21097 12971
rect 20312 12940 21097 12968
rect 20312 12928 20318 12940
rect 21085 12937 21097 12940
rect 21131 12937 21143 12971
rect 21085 12931 21143 12937
rect 6822 12900 6828 12912
rect 5276 12872 6828 12900
rect 6822 12860 6828 12872
rect 6880 12900 6886 12912
rect 9398 12900 9404 12912
rect 6880 12872 9404 12900
rect 6880 12860 6886 12872
rect 9398 12860 9404 12872
rect 9456 12860 9462 12912
rect 3145 12835 3203 12841
rect 3145 12832 3157 12835
rect 2148 12804 3157 12832
rect 2148 12776 2176 12804
rect 3145 12801 3157 12804
rect 3191 12801 3203 12835
rect 9784 12832 9812 12928
rect 17678 12860 17684 12912
rect 17736 12900 17742 12912
rect 17736 12872 19380 12900
rect 17736 12860 17742 12872
rect 3145 12795 3203 12801
rect 8956 12804 10916 12832
rect 8956 12776 8984 12804
rect 2130 12764 2136 12776
rect 2091 12736 2136 12764
rect 2130 12724 2136 12736
rect 2188 12724 2194 12776
rect 2685 12767 2743 12773
rect 2685 12733 2697 12767
rect 2731 12764 2743 12767
rect 2774 12764 2780 12776
rect 2731 12736 2780 12764
rect 2731 12733 2743 12736
rect 2685 12727 2743 12733
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 3326 12724 3332 12776
rect 3384 12764 3390 12776
rect 3513 12767 3571 12773
rect 3513 12764 3525 12767
rect 3384 12736 3525 12764
rect 3384 12724 3390 12736
rect 3513 12733 3525 12736
rect 3559 12733 3571 12767
rect 5166 12764 5172 12776
rect 5127 12736 5172 12764
rect 3513 12727 3571 12733
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 5261 12767 5319 12773
rect 5261 12733 5273 12767
rect 5307 12733 5319 12767
rect 5261 12727 5319 12733
rect 1581 12699 1639 12705
rect 1581 12665 1593 12699
rect 1627 12696 1639 12699
rect 3234 12696 3240 12708
rect 1627 12668 3240 12696
rect 1627 12665 1639 12668
rect 1581 12659 1639 12665
rect 3234 12656 3240 12668
rect 3292 12656 3298 12708
rect 4982 12656 4988 12708
rect 5040 12696 5046 12708
rect 5276 12696 5304 12727
rect 7190 12724 7196 12776
rect 7248 12764 7254 12776
rect 7374 12764 7380 12776
rect 7248 12736 7380 12764
rect 7248 12724 7254 12736
rect 7374 12724 7380 12736
rect 7432 12764 7438 12776
rect 7745 12767 7803 12773
rect 7745 12764 7757 12767
rect 7432 12736 7757 12764
rect 7432 12724 7438 12736
rect 7745 12733 7757 12736
rect 7791 12733 7803 12767
rect 7745 12727 7803 12733
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 8665 12767 8723 12773
rect 8665 12764 8677 12767
rect 8444 12736 8677 12764
rect 8444 12724 8450 12736
rect 8665 12733 8677 12736
rect 8711 12733 8723 12767
rect 8938 12764 8944 12776
rect 8851 12736 8944 12764
rect 8665 12727 8723 12733
rect 8938 12724 8944 12736
rect 8996 12724 9002 12776
rect 9674 12764 9680 12776
rect 9635 12736 9680 12764
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 9861 12767 9919 12773
rect 9861 12733 9873 12767
rect 9907 12764 9919 12767
rect 9950 12764 9956 12776
rect 9907 12736 9956 12764
rect 9907 12733 9919 12736
rect 9861 12727 9919 12733
rect 9950 12724 9956 12736
rect 10008 12724 10014 12776
rect 10134 12724 10140 12776
rect 10192 12764 10198 12776
rect 10594 12764 10600 12776
rect 10192 12736 10600 12764
rect 10192 12724 10198 12736
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 10888 12773 10916 12804
rect 12066 12792 12072 12844
rect 12124 12832 12130 12844
rect 12342 12832 12348 12844
rect 12124 12804 12348 12832
rect 12124 12792 12130 12804
rect 12342 12792 12348 12804
rect 12400 12832 12406 12844
rect 13173 12835 13231 12841
rect 13173 12832 13185 12835
rect 12400 12804 13185 12832
rect 12400 12792 12406 12804
rect 13173 12801 13185 12804
rect 13219 12801 13231 12835
rect 13814 12832 13820 12844
rect 13775 12804 13820 12832
rect 13173 12795 13231 12801
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 14090 12832 14096 12844
rect 14051 12804 14096 12832
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 17313 12835 17371 12841
rect 17313 12801 17325 12835
rect 17359 12832 17371 12835
rect 17402 12832 17408 12844
rect 17359 12804 17408 12832
rect 17359 12801 17371 12804
rect 17313 12795 17371 12801
rect 17402 12792 17408 12804
rect 17460 12792 17466 12844
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12832 17555 12835
rect 18874 12832 18880 12844
rect 17543 12804 18880 12832
rect 17543 12801 17555 12804
rect 17497 12795 17555 12801
rect 18874 12792 18880 12804
rect 18932 12792 18938 12844
rect 19352 12841 19380 12872
rect 19337 12835 19395 12841
rect 19337 12801 19349 12835
rect 19383 12801 19395 12835
rect 19610 12832 19616 12844
rect 19571 12804 19616 12832
rect 19337 12795 19395 12801
rect 19610 12792 19616 12804
rect 19668 12792 19674 12844
rect 10873 12767 10931 12773
rect 10873 12733 10885 12767
rect 10919 12733 10931 12767
rect 11054 12764 11060 12776
rect 11015 12736 11060 12764
rect 10873 12727 10931 12733
rect 11054 12724 11060 12736
rect 11112 12724 11118 12776
rect 13078 12764 13084 12776
rect 13039 12736 13084 12764
rect 13078 12724 13084 12736
rect 13136 12724 13142 12776
rect 16206 12764 16212 12776
rect 16167 12736 16212 12764
rect 16206 12724 16212 12736
rect 16264 12724 16270 12776
rect 17589 12767 17647 12773
rect 17589 12733 17601 12767
rect 17635 12764 17647 12767
rect 18046 12764 18052 12776
rect 17635 12736 18052 12764
rect 17635 12733 17647 12736
rect 17589 12727 17647 12733
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 18509 12767 18567 12773
rect 18509 12733 18521 12767
rect 18555 12764 18567 12767
rect 18598 12764 18604 12776
rect 18555 12736 18604 12764
rect 18555 12733 18567 12736
rect 18509 12727 18567 12733
rect 18598 12724 18604 12736
rect 18656 12724 18662 12776
rect 5040 12668 5304 12696
rect 5040 12656 5046 12668
rect 5276 12628 5304 12668
rect 6914 12656 6920 12708
rect 6972 12696 6978 12708
rect 7561 12699 7619 12705
rect 7561 12696 7573 12699
rect 6972 12668 7573 12696
rect 6972 12656 6978 12668
rect 7561 12665 7573 12668
rect 7607 12696 7619 12699
rect 7650 12696 7656 12708
rect 7607 12668 7656 12696
rect 7607 12665 7619 12668
rect 7561 12659 7619 12665
rect 7650 12656 7656 12668
rect 7708 12656 7714 12708
rect 10413 12699 10471 12705
rect 10413 12665 10425 12699
rect 10459 12696 10471 12699
rect 10459 12668 14504 12696
rect 10459 12665 10471 12668
rect 10413 12659 10471 12665
rect 7837 12631 7895 12637
rect 7837 12628 7849 12631
rect 5276 12600 7849 12628
rect 7837 12597 7849 12600
rect 7883 12628 7895 12631
rect 8202 12628 8208 12640
rect 7883 12600 8208 12628
rect 7883 12597 7895 12600
rect 7837 12591 7895 12597
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 8849 12631 8907 12637
rect 8849 12597 8861 12631
rect 8895 12628 8907 12631
rect 9214 12628 9220 12640
rect 8895 12600 9220 12628
rect 8895 12597 8907 12600
rect 8849 12591 8907 12597
rect 9214 12588 9220 12600
rect 9272 12588 9278 12640
rect 12618 12628 12624 12640
rect 12579 12600 12624 12628
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 12986 12628 12992 12640
rect 12947 12600 12992 12628
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 14476 12628 14504 12668
rect 15102 12656 15108 12708
rect 15160 12656 15166 12708
rect 17770 12656 17776 12708
rect 17828 12696 17834 12708
rect 18693 12699 18751 12705
rect 18693 12696 18705 12699
rect 17828 12668 18705 12696
rect 17828 12656 17834 12668
rect 18693 12665 18705 12668
rect 18739 12665 18751 12699
rect 18693 12659 18751 12665
rect 20622 12656 20628 12708
rect 20680 12656 20686 12708
rect 17954 12628 17960 12640
rect 14476 12600 17960 12628
rect 17954 12588 17960 12600
rect 18012 12588 18018 12640
rect 18874 12628 18880 12640
rect 18835 12600 18880 12628
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 1104 12538 21804 12560
rect 1104 12486 7882 12538
rect 7934 12486 7946 12538
rect 7998 12486 8010 12538
rect 8062 12486 8074 12538
rect 8126 12486 14782 12538
rect 14834 12486 14846 12538
rect 14898 12486 14910 12538
rect 14962 12486 14974 12538
rect 15026 12486 21804 12538
rect 1104 12464 21804 12486
rect 5534 12424 5540 12436
rect 5495 12396 5540 12424
rect 5534 12384 5540 12396
rect 5592 12384 5598 12436
rect 11054 12384 11060 12436
rect 11112 12424 11118 12436
rect 11885 12427 11943 12433
rect 11885 12424 11897 12427
rect 11112 12396 11897 12424
rect 11112 12384 11118 12396
rect 11885 12393 11897 12396
rect 11931 12393 11943 12427
rect 11885 12387 11943 12393
rect 12158 12384 12164 12436
rect 12216 12424 12222 12436
rect 12253 12427 12311 12433
rect 12253 12424 12265 12427
rect 12216 12396 12265 12424
rect 12216 12384 12222 12396
rect 12253 12393 12265 12396
rect 12299 12393 12311 12427
rect 12253 12387 12311 12393
rect 12986 12384 12992 12436
rect 13044 12424 13050 12436
rect 13081 12427 13139 12433
rect 13081 12424 13093 12427
rect 13044 12396 13093 12424
rect 13044 12384 13050 12396
rect 13081 12393 13093 12396
rect 13127 12393 13139 12427
rect 13081 12387 13139 12393
rect 14921 12427 14979 12433
rect 14921 12393 14933 12427
rect 14967 12424 14979 12427
rect 15102 12424 15108 12436
rect 14967 12396 15108 12424
rect 14967 12393 14979 12396
rect 14921 12387 14979 12393
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 20622 12424 20628 12436
rect 20583 12396 20628 12424
rect 20622 12384 20628 12396
rect 20680 12384 20686 12436
rect 3326 12356 3332 12368
rect 3287 12328 3332 12356
rect 3326 12316 3332 12328
rect 3384 12316 3390 12368
rect 11790 12356 11796 12368
rect 11751 12328 11796 12356
rect 11790 12316 11796 12328
rect 11848 12356 11854 12368
rect 12713 12359 12771 12365
rect 12713 12356 12725 12359
rect 11848 12328 12725 12356
rect 11848 12316 11854 12328
rect 12713 12325 12725 12328
rect 12759 12325 12771 12359
rect 12713 12319 12771 12325
rect 2958 12248 2964 12300
rect 3016 12288 3022 12300
rect 3145 12291 3203 12297
rect 3145 12288 3157 12291
rect 3016 12260 3157 12288
rect 3016 12248 3022 12260
rect 3145 12257 3157 12260
rect 3191 12257 3203 12291
rect 3145 12251 3203 12257
rect 5166 12248 5172 12300
rect 5224 12288 5230 12300
rect 5629 12291 5687 12297
rect 5629 12288 5641 12291
rect 5224 12260 5641 12288
rect 5224 12248 5230 12260
rect 5629 12257 5641 12260
rect 5675 12257 5687 12291
rect 5629 12251 5687 12257
rect 5718 12248 5724 12300
rect 5776 12288 5782 12300
rect 6365 12291 6423 12297
rect 6365 12288 6377 12291
rect 5776 12260 6377 12288
rect 5776 12248 5782 12260
rect 6365 12257 6377 12260
rect 6411 12288 6423 12291
rect 6914 12288 6920 12300
rect 6411 12260 6920 12288
rect 6411 12257 6423 12260
rect 6365 12251 6423 12257
rect 6914 12248 6920 12260
rect 6972 12248 6978 12300
rect 7558 12288 7564 12300
rect 7519 12260 7564 12288
rect 7558 12248 7564 12260
rect 7616 12248 7622 12300
rect 12897 12291 12955 12297
rect 12897 12288 12909 12291
rect 12406 12260 12909 12288
rect 5537 12223 5595 12229
rect 5537 12189 5549 12223
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 5552 12152 5580 12183
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 6457 12223 6515 12229
rect 6457 12220 6469 12223
rect 5960 12192 6469 12220
rect 5960 12180 5966 12192
rect 6457 12189 6469 12192
rect 6503 12189 6515 12223
rect 6457 12183 6515 12189
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 6822 12220 6828 12232
rect 6687 12192 6828 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 6181 12155 6239 12161
rect 6181 12152 6193 12155
rect 5552 12124 6193 12152
rect 6181 12121 6193 12124
rect 6227 12121 6239 12155
rect 6181 12115 6239 12121
rect 6564 12152 6592 12183
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 7837 12223 7895 12229
rect 7837 12189 7849 12223
rect 7883 12220 7895 12223
rect 8202 12220 8208 12232
rect 7883 12192 8208 12220
rect 7883 12189 7895 12192
rect 7837 12183 7895 12189
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 10410 12180 10416 12232
rect 10468 12220 10474 12232
rect 11609 12223 11667 12229
rect 11609 12220 11621 12223
rect 10468 12192 11621 12220
rect 10468 12180 10474 12192
rect 11609 12189 11621 12192
rect 11655 12220 11667 12223
rect 12406 12220 12434 12260
rect 12897 12257 12909 12260
rect 12943 12257 12955 12291
rect 12897 12251 12955 12257
rect 14737 12291 14795 12297
rect 14737 12257 14749 12291
rect 14783 12288 14795 12291
rect 16206 12288 16212 12300
rect 14783 12260 16212 12288
rect 14783 12257 14795 12260
rect 14737 12251 14795 12257
rect 16206 12248 16212 12260
rect 16264 12288 16270 12300
rect 20070 12288 20076 12300
rect 16264 12260 20076 12288
rect 16264 12248 16270 12260
rect 20070 12248 20076 12260
rect 20128 12288 20134 12300
rect 20809 12291 20867 12297
rect 20809 12288 20821 12291
rect 20128 12260 20821 12288
rect 20128 12248 20134 12260
rect 20809 12257 20821 12260
rect 20855 12288 20867 12291
rect 20898 12288 20904 12300
rect 20855 12260 20904 12288
rect 20855 12257 20867 12260
rect 20809 12251 20867 12257
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 11655 12192 12434 12220
rect 11655 12189 11667 12192
rect 11609 12183 11667 12189
rect 6730 12152 6736 12164
rect 6564 12124 6736 12152
rect 5074 12084 5080 12096
rect 5035 12056 5080 12084
rect 5074 12044 5080 12056
rect 5132 12044 5138 12096
rect 5626 12044 5632 12096
rect 5684 12084 5690 12096
rect 6564 12084 6592 12124
rect 6730 12112 6736 12124
rect 6788 12112 6794 12164
rect 7466 12112 7472 12164
rect 7524 12152 7530 12164
rect 7745 12155 7803 12161
rect 7745 12152 7757 12155
rect 7524 12124 7757 12152
rect 7524 12112 7530 12124
rect 7745 12121 7757 12124
rect 7791 12121 7803 12155
rect 7745 12115 7803 12121
rect 7650 12084 7656 12096
rect 5684 12056 6592 12084
rect 7611 12056 7656 12084
rect 5684 12044 5690 12056
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 1104 11994 21804 12016
rect 1104 11942 4432 11994
rect 4484 11942 4496 11994
rect 4548 11942 4560 11994
rect 4612 11942 4624 11994
rect 4676 11942 11332 11994
rect 11384 11942 11396 11994
rect 11448 11942 11460 11994
rect 11512 11942 11524 11994
rect 11576 11942 18232 11994
rect 18284 11942 18296 11994
rect 18348 11942 18360 11994
rect 18412 11942 18424 11994
rect 18476 11942 21804 11994
rect 1104 11920 21804 11942
rect 2958 11880 2964 11892
rect 2919 11852 2964 11880
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 7374 11880 7380 11892
rect 5552 11852 7380 11880
rect 5552 11753 5580 11852
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11713 5595 11747
rect 5718 11744 5724 11756
rect 5679 11716 5724 11744
rect 5537 11707 5595 11713
rect 5718 11704 5724 11716
rect 5776 11704 5782 11756
rect 5994 11704 6000 11756
rect 6052 11744 6058 11756
rect 6822 11744 6828 11756
rect 6052 11716 6828 11744
rect 6052 11704 6058 11716
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 2961 11679 3019 11685
rect 2961 11676 2973 11679
rect 2832 11648 2973 11676
rect 2832 11636 2838 11648
rect 2961 11645 2973 11648
rect 3007 11645 3019 11679
rect 3510 11676 3516 11688
rect 3471 11648 3516 11676
rect 2961 11639 3019 11645
rect 2976 11608 3004 11639
rect 3510 11636 3516 11648
rect 3568 11636 3574 11688
rect 5626 11636 5632 11688
rect 5684 11676 5690 11688
rect 7208 11685 7236 11852
rect 7374 11840 7380 11852
rect 7432 11840 7438 11892
rect 8202 11840 8208 11892
rect 8260 11880 8266 11892
rect 8389 11883 8447 11889
rect 8389 11880 8401 11883
rect 8260 11852 8401 11880
rect 8260 11840 8266 11852
rect 8389 11849 8401 11852
rect 8435 11849 8447 11883
rect 8389 11843 8447 11849
rect 9214 11840 9220 11892
rect 9272 11880 9278 11892
rect 9272 11852 10824 11880
rect 9272 11840 9278 11852
rect 9401 11815 9459 11821
rect 9401 11812 9413 11815
rect 8036 11784 9413 11812
rect 7650 11704 7656 11756
rect 7708 11744 7714 11756
rect 7929 11747 7987 11753
rect 7929 11744 7941 11747
rect 7708 11716 7941 11744
rect 7708 11704 7714 11716
rect 7929 11713 7941 11716
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 8036 11685 8064 11784
rect 9401 11781 9413 11784
rect 9447 11781 9459 11815
rect 9401 11775 9459 11781
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11744 8263 11747
rect 8938 11744 8944 11756
rect 8251 11716 8944 11744
rect 8251 11713 8263 11716
rect 8205 11707 8263 11713
rect 8938 11704 8944 11716
rect 8996 11744 9002 11756
rect 8996 11716 9628 11744
rect 8996 11704 9002 11716
rect 5813 11679 5871 11685
rect 5684 11648 5729 11676
rect 5684 11636 5690 11648
rect 5813 11645 5825 11679
rect 5859 11676 5871 11679
rect 7009 11679 7067 11685
rect 7009 11676 7021 11679
rect 5859 11648 7021 11676
rect 5859 11645 5871 11648
rect 5813 11639 5871 11645
rect 7009 11645 7021 11648
rect 7055 11645 7067 11679
rect 7009 11639 7067 11645
rect 7193 11679 7251 11685
rect 7193 11645 7205 11679
rect 7239 11676 7251 11679
rect 8021 11679 8079 11685
rect 8021 11676 8033 11679
rect 7239 11648 8033 11676
rect 7239 11645 7251 11648
rect 7193 11639 7251 11645
rect 8021 11645 8033 11648
rect 8067 11645 8079 11679
rect 8021 11639 8079 11645
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11676 8171 11679
rect 9306 11676 9312 11688
rect 8159 11648 9312 11676
rect 8159 11645 8171 11648
rect 8113 11639 8171 11645
rect 4062 11608 4068 11620
rect 2976 11580 4068 11608
rect 4062 11568 4068 11580
rect 4120 11568 4126 11620
rect 5258 11568 5264 11620
rect 5316 11608 5322 11620
rect 5828 11608 5856 11639
rect 5316 11580 5856 11608
rect 7024 11608 7052 11639
rect 7282 11608 7288 11620
rect 7024 11580 7288 11608
rect 5316 11568 5322 11580
rect 7282 11568 7288 11580
rect 7340 11568 7346 11620
rect 7742 11568 7748 11620
rect 7800 11608 7806 11620
rect 8128 11608 8156 11639
rect 9306 11636 9312 11648
rect 9364 11636 9370 11688
rect 9600 11685 9628 11716
rect 10318 11704 10324 11756
rect 10376 11744 10382 11756
rect 10505 11747 10563 11753
rect 10505 11744 10517 11747
rect 10376 11716 10517 11744
rect 10376 11704 10382 11716
rect 10505 11713 10517 11716
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 10796 11685 10824 11852
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11645 9643 11679
rect 10597 11679 10655 11685
rect 10597 11676 10609 11679
rect 9585 11639 9643 11645
rect 9784 11648 10609 11676
rect 9674 11608 9680 11620
rect 7800 11580 8156 11608
rect 9600 11580 9680 11608
rect 7800 11568 7806 11580
rect 4982 11500 4988 11552
rect 5040 11540 5046 11552
rect 5353 11543 5411 11549
rect 5353 11540 5365 11543
rect 5040 11512 5365 11540
rect 5040 11500 5046 11512
rect 5353 11509 5365 11512
rect 5399 11509 5411 11543
rect 7300 11540 7328 11568
rect 9600 11540 9628 11580
rect 9674 11568 9680 11580
rect 9732 11568 9738 11620
rect 9784 11552 9812 11648
rect 10597 11645 10609 11648
rect 10643 11645 10655 11679
rect 10597 11639 10655 11645
rect 10781 11679 10839 11685
rect 10781 11645 10793 11679
rect 10827 11645 10839 11679
rect 10781 11639 10839 11645
rect 9766 11540 9772 11552
rect 7300 11512 9628 11540
rect 9727 11512 9772 11540
rect 5353 11503 5411 11509
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 10965 11543 11023 11549
rect 10965 11509 10977 11543
rect 11011 11540 11023 11543
rect 18414 11540 18420 11552
rect 11011 11512 18420 11540
rect 11011 11509 11023 11512
rect 10965 11503 11023 11509
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 1104 11450 21804 11472
rect 1104 11398 7882 11450
rect 7934 11398 7946 11450
rect 7998 11398 8010 11450
rect 8062 11398 8074 11450
rect 8126 11398 14782 11450
rect 14834 11398 14846 11450
rect 14898 11398 14910 11450
rect 14962 11398 14974 11450
rect 15026 11398 21804 11450
rect 1104 11376 21804 11398
rect 1854 11296 1860 11348
rect 1912 11336 1918 11348
rect 2041 11339 2099 11345
rect 2041 11336 2053 11339
rect 1912 11308 2053 11336
rect 1912 11296 1918 11308
rect 2041 11305 2053 11308
rect 2087 11305 2099 11339
rect 2958 11336 2964 11348
rect 2919 11308 2964 11336
rect 2041 11299 2099 11305
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 4356 11308 8953 11336
rect 4246 11268 4252 11280
rect 2746 11240 4252 11268
rect 1949 11203 2007 11209
rect 1949 11169 1961 11203
rect 1995 11200 2007 11203
rect 2746 11200 2774 11240
rect 4246 11228 4252 11240
rect 4304 11228 4310 11280
rect 4356 11200 4384 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 8941 11299 8999 11305
rect 9766 11296 9772 11348
rect 9824 11336 9830 11348
rect 10250 11339 10308 11345
rect 10250 11336 10262 11339
rect 9824 11308 10262 11336
rect 9824 11296 9830 11308
rect 10250 11305 10262 11308
rect 10296 11305 10308 11339
rect 10250 11299 10308 11305
rect 12710 11296 12716 11348
rect 12768 11336 12774 11348
rect 12897 11339 12955 11345
rect 12897 11336 12909 11339
rect 12768 11308 12909 11336
rect 12768 11296 12774 11308
rect 12897 11305 12909 11308
rect 12943 11305 12955 11339
rect 18509 11339 18567 11345
rect 12897 11299 12955 11305
rect 15028 11308 18368 11336
rect 5626 11228 5632 11280
rect 5684 11268 5690 11280
rect 7009 11271 7067 11277
rect 5684 11240 6316 11268
rect 5684 11228 5690 11240
rect 1995 11172 2774 11200
rect 3988 11172 4384 11200
rect 4433 11203 4491 11209
rect 1995 11169 2007 11172
rect 1949 11163 2007 11169
rect 2222 11132 2228 11144
rect 2183 11104 2228 11132
rect 2222 11092 2228 11104
rect 2280 11092 2286 11144
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 3329 11135 3387 11141
rect 3329 11101 3341 11135
rect 3375 11132 3387 11135
rect 3510 11132 3516 11144
rect 3375 11104 3516 11132
rect 3375 11101 3387 11104
rect 3329 11095 3387 11101
rect 2976 11064 3004 11095
rect 3510 11092 3516 11104
rect 3568 11132 3574 11144
rect 3988 11132 4016 11172
rect 4433 11169 4445 11203
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 3568 11104 4016 11132
rect 3568 11092 3574 11104
rect 4062 11092 4068 11144
rect 4120 11132 4126 11144
rect 4448 11132 4476 11163
rect 5534 11160 5540 11212
rect 5592 11200 5598 11212
rect 5902 11200 5908 11212
rect 5592 11172 5908 11200
rect 5592 11160 5598 11172
rect 5902 11160 5908 11172
rect 5960 11200 5966 11212
rect 6288 11209 6316 11240
rect 7009 11237 7021 11271
rect 7055 11268 7067 11271
rect 7055 11240 7696 11268
rect 7055 11237 7067 11240
rect 7009 11231 7067 11237
rect 7668 11212 7696 11240
rect 9674 11228 9680 11280
rect 9732 11268 9738 11280
rect 10042 11268 10048 11280
rect 9732 11240 10048 11268
rect 9732 11228 9738 11240
rect 10042 11228 10048 11240
rect 10100 11268 10106 11280
rect 10410 11268 10416 11280
rect 10100 11240 10416 11268
rect 10100 11228 10106 11240
rect 10410 11228 10416 11240
rect 10468 11228 10474 11280
rect 11609 11271 11667 11277
rect 11609 11237 11621 11271
rect 11655 11268 11667 11271
rect 11698 11268 11704 11280
rect 11655 11240 11704 11268
rect 11655 11237 11667 11240
rect 11609 11231 11667 11237
rect 11698 11228 11704 11240
rect 11756 11228 11762 11280
rect 11793 11271 11851 11277
rect 11793 11237 11805 11271
rect 11839 11268 11851 11271
rect 15028 11268 15056 11308
rect 18138 11268 18144 11280
rect 11839 11240 15056 11268
rect 15120 11240 18144 11268
rect 11839 11237 11851 11240
rect 11793 11231 11851 11237
rect 6170 11203 6228 11209
rect 6170 11200 6182 11203
rect 5960 11172 6182 11200
rect 5960 11160 5966 11172
rect 6170 11169 6182 11172
rect 6216 11169 6228 11203
rect 6170 11163 6228 11169
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11169 6331 11203
rect 6273 11163 6331 11169
rect 6822 11160 6828 11212
rect 6880 11200 6886 11212
rect 6917 11203 6975 11209
rect 6917 11200 6929 11203
rect 6880 11172 6929 11200
rect 6880 11160 6886 11172
rect 6917 11169 6929 11172
rect 6963 11169 6975 11203
rect 6917 11163 6975 11169
rect 7098 11160 7104 11212
rect 7156 11200 7162 11212
rect 7561 11203 7619 11209
rect 7561 11200 7573 11203
rect 7156 11172 7573 11200
rect 7156 11160 7162 11172
rect 7561 11169 7573 11172
rect 7607 11169 7619 11203
rect 7561 11163 7619 11169
rect 7650 11160 7656 11212
rect 7708 11200 7714 11212
rect 7745 11203 7803 11209
rect 7745 11200 7757 11203
rect 7708 11172 7757 11200
rect 7708 11160 7714 11172
rect 7745 11169 7757 11172
rect 7791 11169 7803 11203
rect 7745 11163 7803 11169
rect 8113 11203 8171 11209
rect 8113 11169 8125 11203
rect 8159 11200 8171 11203
rect 8202 11200 8208 11212
rect 8159 11172 8208 11200
rect 8159 11169 8171 11172
rect 8113 11163 8171 11169
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 12989 11203 13047 11209
rect 12989 11200 13001 11203
rect 8312 11172 13001 11200
rect 4120 11104 4476 11132
rect 4120 11092 4126 11104
rect 5994 11092 6000 11144
rect 6052 11132 6058 11144
rect 6089 11135 6147 11141
rect 6089 11132 6101 11135
rect 6052 11104 6101 11132
rect 6052 11092 6058 11104
rect 6089 11101 6101 11104
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 6365 11135 6423 11141
rect 6365 11101 6377 11135
rect 6411 11132 6423 11135
rect 7374 11132 7380 11144
rect 6411 11104 7380 11132
rect 6411 11101 6423 11104
rect 6365 11095 6423 11101
rect 7374 11092 7380 11104
rect 7432 11132 7438 11144
rect 8312 11132 8340 11172
rect 12989 11169 13001 11172
rect 13035 11169 13047 11203
rect 15010 11200 15016 11212
rect 14971 11172 15016 11200
rect 12989 11163 13047 11169
rect 15010 11160 15016 11172
rect 15068 11160 15074 11212
rect 7432 11104 8340 11132
rect 8941 11135 8999 11141
rect 7432 11092 7438 11104
rect 8941 11101 8953 11135
rect 8987 11132 8999 11135
rect 11885 11135 11943 11141
rect 8987 11104 11376 11132
rect 8987 11101 8999 11104
rect 8941 11095 8999 11101
rect 4249 11067 4307 11073
rect 4249 11064 4261 11067
rect 2976 11036 4261 11064
rect 4249 11033 4261 11036
rect 4295 11033 4307 11067
rect 4249 11027 4307 11033
rect 7282 11024 7288 11076
rect 7340 11064 7346 11076
rect 7745 11067 7803 11073
rect 7745 11064 7757 11067
rect 7340 11036 7757 11064
rect 7340 11024 7346 11036
rect 7745 11033 7757 11036
rect 7791 11033 7803 11067
rect 10410 11064 10416 11076
rect 10371 11036 10416 11064
rect 7745 11027 7803 11033
rect 10410 11024 10416 11036
rect 10468 11064 10474 11076
rect 10594 11064 10600 11076
rect 10468 11036 10600 11064
rect 10468 11024 10474 11036
rect 10594 11024 10600 11036
rect 10652 11024 10658 11076
rect 11348 11073 11376 11104
rect 11885 11101 11897 11135
rect 11931 11132 11943 11135
rect 12342 11132 12348 11144
rect 11931 11104 12348 11132
rect 11931 11101 11943 11104
rect 11885 11095 11943 11101
rect 12342 11092 12348 11104
rect 12400 11132 12406 11144
rect 12713 11135 12771 11141
rect 12713 11132 12725 11135
rect 12400 11104 12725 11132
rect 12400 11092 12406 11104
rect 12713 11101 12725 11104
rect 12759 11132 12771 11135
rect 15120 11132 15148 11240
rect 18138 11228 18144 11240
rect 18196 11228 18202 11280
rect 18340 11268 18368 11308
rect 18509 11305 18521 11339
rect 18555 11336 18567 11339
rect 20990 11336 20996 11348
rect 18555 11308 20996 11336
rect 18555 11305 18567 11308
rect 18509 11299 18567 11305
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 20898 11268 20904 11280
rect 18340 11240 20904 11268
rect 20898 11228 20904 11240
rect 20956 11228 20962 11280
rect 16942 11200 16948 11212
rect 16903 11172 16948 11200
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 17405 11203 17463 11209
rect 17405 11169 17417 11203
rect 17451 11169 17463 11203
rect 18414 11200 18420 11212
rect 18375 11172 18420 11200
rect 17405 11163 17463 11169
rect 16482 11132 16488 11144
rect 12759 11104 15148 11132
rect 15212 11104 16488 11132
rect 12759 11101 12771 11104
rect 12713 11095 12771 11101
rect 15212 11076 15240 11104
rect 16482 11092 16488 11104
rect 16540 11132 16546 11144
rect 17420 11132 17448 11163
rect 18414 11160 18420 11172
rect 18472 11160 18478 11212
rect 20070 11200 20076 11212
rect 20031 11172 20076 11200
rect 20070 11160 20076 11172
rect 20128 11160 20134 11212
rect 16540 11104 17448 11132
rect 16540 11092 16546 11104
rect 18322 11092 18328 11144
rect 18380 11132 18386 11144
rect 18598 11132 18604 11144
rect 18380 11104 18604 11132
rect 18380 11092 18386 11104
rect 18598 11092 18604 11104
rect 18656 11092 18662 11144
rect 11333 11067 11391 11073
rect 11333 11033 11345 11067
rect 11379 11033 11391 11067
rect 11333 11027 11391 11033
rect 13357 11067 13415 11073
rect 13357 11033 13369 11067
rect 13403 11064 13415 11067
rect 14826 11064 14832 11076
rect 13403 11036 14832 11064
rect 13403 11033 13415 11036
rect 13357 11027 13415 11033
rect 14826 11024 14832 11036
rect 14884 11024 14890 11076
rect 15194 11064 15200 11076
rect 15155 11036 15200 11064
rect 15194 11024 15200 11036
rect 15252 11024 15258 11076
rect 17589 11067 17647 11073
rect 17589 11033 17601 11067
rect 17635 11064 17647 11067
rect 18046 11064 18052 11076
rect 17635 11036 17908 11064
rect 18007 11036 18052 11064
rect 17635 11033 17647 11036
rect 17589 11027 17647 11033
rect 1578 10996 1584 11008
rect 1539 10968 1584 10996
rect 1578 10956 1584 10968
rect 1636 10956 1642 11008
rect 5902 10996 5908 11008
rect 5863 10968 5908 10996
rect 5902 10956 5908 10968
rect 5960 10956 5966 11008
rect 9858 10956 9864 11008
rect 9916 10996 9922 11008
rect 10226 10996 10232 11008
rect 9916 10968 10232 10996
rect 9916 10956 9922 10968
rect 10226 10956 10232 10968
rect 10284 10956 10290 11008
rect 16850 10996 16856 11008
rect 16811 10968 16856 10996
rect 16850 10956 16856 10968
rect 16908 10956 16914 11008
rect 17880 10996 17908 11036
rect 18046 11024 18052 11036
rect 18104 11024 18110 11076
rect 20162 11024 20168 11076
rect 20220 11064 20226 11076
rect 20257 11067 20315 11073
rect 20257 11064 20269 11067
rect 20220 11036 20269 11064
rect 20220 11024 20226 11036
rect 20257 11033 20269 11036
rect 20303 11033 20315 11067
rect 20257 11027 20315 11033
rect 18690 10996 18696 11008
rect 17880 10968 18696 10996
rect 18690 10956 18696 10968
rect 18748 10956 18754 11008
rect 1104 10906 21804 10928
rect 1104 10854 4432 10906
rect 4484 10854 4496 10906
rect 4548 10854 4560 10906
rect 4612 10854 4624 10906
rect 4676 10854 11332 10906
rect 11384 10854 11396 10906
rect 11448 10854 11460 10906
rect 11512 10854 11524 10906
rect 11576 10854 18232 10906
rect 18284 10854 18296 10906
rect 18348 10854 18360 10906
rect 18412 10854 18424 10906
rect 18476 10854 21804 10906
rect 1104 10832 21804 10854
rect 4246 10752 4252 10804
rect 4304 10792 4310 10804
rect 4617 10795 4675 10801
rect 4617 10792 4629 10795
rect 4304 10764 4629 10792
rect 4304 10752 4310 10764
rect 4617 10761 4629 10764
rect 4663 10761 4675 10795
rect 4617 10755 4675 10761
rect 4890 10752 4896 10804
rect 4948 10792 4954 10804
rect 4985 10795 5043 10801
rect 4985 10792 4997 10795
rect 4948 10764 4997 10792
rect 4948 10752 4954 10764
rect 4985 10761 4997 10764
rect 5031 10761 5043 10795
rect 7558 10792 7564 10804
rect 7519 10764 7564 10792
rect 4985 10755 5043 10761
rect 7558 10752 7564 10764
rect 7616 10752 7622 10804
rect 13449 10795 13507 10801
rect 13449 10761 13461 10795
rect 13495 10792 13507 10795
rect 13814 10792 13820 10804
rect 13495 10764 13820 10792
rect 13495 10761 13507 10764
rect 13449 10755 13507 10761
rect 13814 10752 13820 10764
rect 13872 10792 13878 10804
rect 15010 10792 15016 10804
rect 13872 10764 15016 10792
rect 13872 10752 13878 10764
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 20438 10752 20444 10804
rect 20496 10792 20502 10804
rect 20901 10795 20959 10801
rect 20901 10792 20913 10795
rect 20496 10764 20913 10792
rect 20496 10752 20502 10764
rect 20901 10761 20913 10764
rect 20947 10761 20959 10795
rect 20901 10755 20959 10761
rect 7650 10684 7656 10736
rect 7708 10684 7714 10736
rect 16209 10727 16267 10733
rect 16209 10693 16221 10727
rect 16255 10724 16267 10727
rect 16850 10724 16856 10736
rect 16255 10696 16856 10724
rect 16255 10693 16267 10696
rect 16209 10687 16267 10693
rect 16850 10684 16856 10696
rect 16908 10684 16914 10736
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10656 5135 10659
rect 5626 10656 5632 10668
rect 5123 10628 5632 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 5626 10616 5632 10628
rect 5684 10616 5690 10668
rect 7377 10659 7435 10665
rect 7377 10625 7389 10659
rect 7423 10656 7435 10659
rect 7668 10656 7696 10684
rect 9674 10656 9680 10668
rect 7423 10628 7696 10656
rect 9048 10628 9680 10656
rect 7423 10625 7435 10628
rect 7377 10619 7435 10625
rect 2682 10588 2688 10600
rect 2643 10560 2688 10588
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 4801 10591 4859 10597
rect 4801 10557 4813 10591
rect 4847 10588 4859 10591
rect 5258 10588 5264 10600
rect 4847 10560 5264 10588
rect 4847 10557 4859 10560
rect 4801 10551 4859 10557
rect 5258 10548 5264 10560
rect 5316 10548 5322 10600
rect 7653 10591 7711 10597
rect 7653 10557 7665 10591
rect 7699 10588 7711 10591
rect 7742 10588 7748 10600
rect 7699 10560 7748 10588
rect 7699 10557 7711 10560
rect 7653 10551 7711 10557
rect 7742 10548 7748 10560
rect 7800 10548 7806 10600
rect 9048 10597 9076 10628
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 12618 10616 12624 10668
rect 12676 10656 12682 10668
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 12676 10628 13093 10656
rect 12676 10616 12682 10628
rect 13081 10625 13093 10628
rect 13127 10625 13139 10659
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 13081 10619 13139 10625
rect 14844 10628 15853 10656
rect 14844 10600 14872 10628
rect 15841 10625 15853 10628
rect 15887 10625 15899 10659
rect 15841 10619 15899 10625
rect 18325 10659 18383 10665
rect 18325 10625 18337 10659
rect 18371 10656 18383 10659
rect 18598 10656 18604 10668
rect 18371 10628 18604 10656
rect 18371 10625 18383 10628
rect 18325 10619 18383 10625
rect 18598 10616 18604 10628
rect 18656 10616 18662 10668
rect 18874 10616 18880 10668
rect 18932 10656 18938 10668
rect 19429 10659 19487 10665
rect 19429 10656 19441 10659
rect 18932 10628 19441 10656
rect 18932 10616 18938 10628
rect 19429 10625 19441 10628
rect 19475 10625 19487 10659
rect 19429 10619 19487 10625
rect 9033 10591 9091 10597
rect 9033 10557 9045 10591
rect 9079 10557 9091 10591
rect 9033 10551 9091 10557
rect 9490 10548 9496 10600
rect 9548 10588 9554 10600
rect 9585 10591 9643 10597
rect 9585 10588 9597 10591
rect 9548 10560 9597 10588
rect 9548 10548 9554 10560
rect 9585 10557 9597 10560
rect 9631 10557 9643 10591
rect 13446 10588 13452 10600
rect 13407 10560 13452 10588
rect 9585 10551 9643 10557
rect 13446 10548 13452 10560
rect 13504 10548 13510 10600
rect 14826 10588 14832 10600
rect 14787 10560 14832 10588
rect 14826 10548 14832 10560
rect 14884 10548 14890 10600
rect 15194 10548 15200 10600
rect 15252 10588 15258 10600
rect 15381 10591 15439 10597
rect 15381 10588 15393 10591
rect 15252 10560 15393 10588
rect 15252 10548 15258 10560
rect 15381 10557 15393 10560
rect 15427 10557 15439 10591
rect 15381 10551 15439 10557
rect 17678 10548 17684 10600
rect 17736 10548 17742 10600
rect 17954 10548 17960 10600
rect 18012 10588 18018 10600
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 18012 10560 18061 10588
rect 18012 10548 18018 10560
rect 18049 10557 18061 10560
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 19153 10591 19211 10597
rect 19153 10557 19165 10591
rect 19199 10557 19211 10591
rect 19153 10551 19211 10557
rect 1581 10523 1639 10529
rect 1581 10489 1593 10523
rect 1627 10520 1639 10523
rect 2038 10520 2044 10532
rect 1627 10492 2044 10520
rect 1627 10489 1639 10492
rect 1581 10483 1639 10489
rect 2038 10480 2044 10492
rect 2096 10480 2102 10532
rect 2866 10520 2872 10532
rect 2827 10492 2872 10520
rect 2866 10480 2872 10492
rect 2924 10480 2930 10532
rect 8478 10520 8484 10532
rect 8439 10492 8484 10520
rect 8478 10480 8484 10492
rect 8536 10480 8542 10532
rect 15289 10523 15347 10529
rect 15289 10489 15301 10523
rect 15335 10489 15347 10523
rect 15289 10483 15347 10489
rect 1486 10452 1492 10464
rect 1447 10424 1492 10452
rect 1486 10412 1492 10424
rect 1544 10412 1550 10464
rect 7377 10455 7435 10461
rect 7377 10421 7389 10455
rect 7423 10452 7435 10455
rect 7650 10452 7656 10464
rect 7423 10424 7656 10452
rect 7423 10421 7435 10424
rect 7377 10415 7435 10421
rect 7650 10412 7656 10424
rect 7708 10412 7714 10464
rect 8570 10412 8576 10464
rect 8628 10452 8634 10464
rect 9582 10452 9588 10464
rect 8628 10424 9588 10452
rect 8628 10412 8634 10424
rect 9582 10412 9588 10424
rect 9640 10452 9646 10464
rect 9677 10455 9735 10461
rect 9677 10452 9689 10455
rect 9640 10424 9689 10452
rect 9640 10412 9646 10424
rect 9677 10421 9689 10424
rect 9723 10421 9735 10455
rect 15304 10452 15332 10483
rect 17402 10480 17408 10532
rect 17460 10520 17466 10532
rect 17696 10520 17724 10548
rect 19168 10520 19196 10551
rect 17460 10492 19196 10520
rect 17460 10480 17466 10492
rect 20162 10480 20168 10532
rect 20220 10480 20226 10532
rect 16209 10455 16267 10461
rect 16209 10452 16221 10455
rect 15304 10424 16221 10452
rect 9677 10415 9735 10421
rect 16209 10421 16221 10424
rect 16255 10452 16267 10455
rect 17310 10452 17316 10464
rect 16255 10424 17316 10452
rect 16255 10421 16267 10424
rect 16209 10415 16267 10421
rect 17310 10412 17316 10424
rect 17368 10412 17374 10464
rect 17681 10455 17739 10461
rect 17681 10421 17693 10455
rect 17727 10452 17739 10455
rect 17770 10452 17776 10464
rect 17727 10424 17776 10452
rect 17727 10421 17739 10424
rect 17681 10415 17739 10421
rect 17770 10412 17776 10424
rect 17828 10412 17834 10464
rect 18141 10455 18199 10461
rect 18141 10421 18153 10455
rect 18187 10452 18199 10455
rect 18782 10452 18788 10464
rect 18187 10424 18788 10452
rect 18187 10421 18199 10424
rect 18141 10415 18199 10421
rect 18782 10412 18788 10424
rect 18840 10412 18846 10464
rect 1104 10362 21804 10384
rect 1104 10310 7882 10362
rect 7934 10310 7946 10362
rect 7998 10310 8010 10362
rect 8062 10310 8074 10362
rect 8126 10310 14782 10362
rect 14834 10310 14846 10362
rect 14898 10310 14910 10362
rect 14962 10310 14974 10362
rect 15026 10310 21804 10362
rect 1104 10288 21804 10310
rect 2222 10248 2228 10260
rect 2183 10220 2228 10248
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 5261 10251 5319 10257
rect 5261 10217 5273 10251
rect 5307 10248 5319 10251
rect 5350 10248 5356 10260
rect 5307 10220 5356 10248
rect 5307 10217 5319 10220
rect 5261 10211 5319 10217
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 6733 10251 6791 10257
rect 6733 10217 6745 10251
rect 6779 10248 6791 10251
rect 7006 10248 7012 10260
rect 6779 10220 7012 10248
rect 6779 10217 6791 10220
rect 6733 10211 6791 10217
rect 7006 10208 7012 10220
rect 7064 10208 7070 10260
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 7561 10251 7619 10257
rect 7561 10248 7573 10251
rect 7432 10220 7573 10248
rect 7432 10208 7438 10220
rect 7561 10217 7573 10220
rect 7607 10217 7619 10251
rect 7561 10211 7619 10217
rect 11885 10251 11943 10257
rect 11885 10217 11897 10251
rect 11931 10248 11943 10251
rect 12434 10248 12440 10260
rect 11931 10220 12440 10248
rect 11931 10217 11943 10220
rect 11885 10211 11943 10217
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 18233 10251 18291 10257
rect 18233 10217 18245 10251
rect 18279 10217 18291 10251
rect 20898 10248 20904 10260
rect 20859 10220 20904 10248
rect 18233 10211 18291 10217
rect 5445 10183 5503 10189
rect 5445 10149 5457 10183
rect 5491 10180 5503 10183
rect 5902 10180 5908 10192
rect 5491 10152 5908 10180
rect 5491 10149 5503 10152
rect 5445 10143 5503 10149
rect 5902 10140 5908 10152
rect 5960 10140 5966 10192
rect 6641 10183 6699 10189
rect 6641 10149 6653 10183
rect 6687 10180 6699 10183
rect 9214 10180 9220 10192
rect 6687 10152 9220 10180
rect 6687 10149 6699 10152
rect 6641 10143 6699 10149
rect 1578 10072 1584 10124
rect 1636 10112 1642 10124
rect 1857 10115 1915 10121
rect 1857 10112 1869 10115
rect 1636 10084 1869 10112
rect 1636 10072 1642 10084
rect 1857 10081 1869 10084
rect 1903 10081 1915 10115
rect 1857 10075 1915 10081
rect 7653 10115 7711 10121
rect 7653 10081 7665 10115
rect 7699 10112 7711 10115
rect 8202 10112 8208 10124
rect 7699 10084 8208 10112
rect 7699 10081 7711 10084
rect 7653 10075 7711 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 8312 10121 8340 10152
rect 9214 10140 9220 10152
rect 9272 10180 9278 10192
rect 13357 10183 13415 10189
rect 9272 10152 9996 10180
rect 9272 10140 9278 10152
rect 8297 10115 8355 10121
rect 8297 10081 8309 10115
rect 8343 10081 8355 10115
rect 8570 10112 8576 10124
rect 8531 10084 8576 10112
rect 8297 10075 8355 10081
rect 8570 10072 8576 10084
rect 8628 10072 8634 10124
rect 9398 10072 9404 10124
rect 9456 10112 9462 10124
rect 9968 10121 9996 10152
rect 13357 10149 13369 10183
rect 13403 10180 13415 10183
rect 13814 10180 13820 10192
rect 13403 10152 13820 10180
rect 13403 10149 13415 10152
rect 13357 10143 13415 10149
rect 13814 10140 13820 10152
rect 13872 10140 13878 10192
rect 16942 10140 16948 10192
rect 17000 10180 17006 10192
rect 17313 10183 17371 10189
rect 17313 10180 17325 10183
rect 17000 10152 17325 10180
rect 17000 10140 17006 10152
rect 17313 10149 17325 10152
rect 17359 10180 17371 10183
rect 18248 10180 18276 10211
rect 20898 10208 20904 10220
rect 20956 10208 20962 10260
rect 17359 10152 18276 10180
rect 17359 10149 17371 10152
rect 17313 10143 17371 10149
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 9456 10084 9689 10112
rect 9456 10072 9462 10084
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 9953 10115 10011 10121
rect 9953 10081 9965 10115
rect 9999 10081 10011 10115
rect 9953 10075 10011 10081
rect 12618 10072 12624 10124
rect 12676 10112 12682 10124
rect 12897 10115 12955 10121
rect 12897 10112 12909 10115
rect 12676 10084 12909 10112
rect 12676 10072 12682 10084
rect 12897 10081 12909 10084
rect 12943 10081 12955 10115
rect 12897 10075 12955 10081
rect 12986 10072 12992 10124
rect 13044 10112 13050 10124
rect 13449 10115 13507 10121
rect 13449 10112 13461 10115
rect 13044 10084 13461 10112
rect 13044 10072 13050 10084
rect 13449 10081 13461 10084
rect 13495 10081 13507 10115
rect 13449 10075 13507 10081
rect 16482 10072 16488 10124
rect 16540 10112 16546 10124
rect 17221 10115 17279 10121
rect 17221 10112 17233 10115
rect 16540 10084 17233 10112
rect 16540 10072 16546 10084
rect 17221 10081 17233 10084
rect 17267 10081 17279 10115
rect 17770 10112 17776 10124
rect 17731 10084 17776 10112
rect 17221 10075 17279 10081
rect 17770 10072 17776 10084
rect 17828 10112 17834 10124
rect 18601 10115 18659 10121
rect 18601 10112 18613 10115
rect 17828 10084 18613 10112
rect 17828 10072 17834 10084
rect 18601 10081 18613 10084
rect 18647 10081 18659 10115
rect 21082 10112 21088 10124
rect 21043 10084 21088 10112
rect 18601 10075 18659 10081
rect 21082 10072 21088 10084
rect 21140 10072 21146 10124
rect 5166 10044 5172 10056
rect 5127 10016 5172 10044
rect 5166 10004 5172 10016
rect 5224 10044 5230 10056
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 5224 10016 6837 10044
rect 5224 10004 5230 10016
rect 6825 10013 6837 10016
rect 6871 10013 6883 10047
rect 6825 10007 6883 10013
rect 8481 10047 8539 10053
rect 8481 10013 8493 10047
rect 8527 10044 8539 10047
rect 9766 10044 9772 10056
rect 8527 10016 9772 10044
rect 8527 10013 8539 10016
rect 8481 10007 8539 10013
rect 9766 10004 9772 10016
rect 9824 10004 9830 10056
rect 11146 10004 11152 10056
rect 11204 10044 11210 10056
rect 11517 10047 11575 10053
rect 11517 10044 11529 10047
rect 11204 10016 11529 10044
rect 11204 10004 11210 10016
rect 11517 10013 11529 10016
rect 11563 10013 11575 10047
rect 11517 10007 11575 10013
rect 18233 10047 18291 10053
rect 18233 10013 18245 10047
rect 18279 10044 18291 10047
rect 18690 10044 18696 10056
rect 18279 10016 18696 10044
rect 18279 10013 18291 10016
rect 18233 10007 18291 10013
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 2225 9979 2283 9985
rect 2225 9945 2237 9979
rect 2271 9976 2283 9979
rect 2774 9976 2780 9988
rect 2271 9948 2780 9976
rect 2271 9945 2283 9948
rect 2225 9939 2283 9945
rect 2774 9936 2780 9948
rect 2832 9936 2838 9988
rect 5721 9979 5779 9985
rect 5721 9945 5733 9979
rect 5767 9976 5779 9979
rect 10226 9976 10232 9988
rect 5767 9948 10232 9976
rect 5767 9945 5779 9948
rect 5721 9939 5779 9945
rect 10226 9936 10232 9948
rect 10284 9936 10290 9988
rect 11882 9976 11888 9988
rect 11843 9948 11888 9976
rect 11882 9936 11888 9948
rect 11940 9936 11946 9988
rect 6178 9868 6184 9920
rect 6236 9908 6242 9920
rect 6273 9911 6331 9917
rect 6273 9908 6285 9911
rect 6236 9880 6285 9908
rect 6236 9868 6242 9880
rect 6273 9877 6285 9880
rect 6319 9877 6331 9911
rect 6273 9871 6331 9877
rect 8113 9911 8171 9917
rect 8113 9877 8125 9911
rect 8159 9908 8171 9911
rect 8754 9908 8760 9920
rect 8159 9880 8760 9908
rect 8159 9877 8171 9880
rect 8113 9871 8171 9877
rect 8754 9868 8760 9880
rect 8812 9868 8818 9920
rect 10137 9911 10195 9917
rect 10137 9877 10149 9911
rect 10183 9908 10195 9911
rect 13354 9908 13360 9920
rect 10183 9880 13360 9908
rect 10183 9877 10195 9880
rect 10137 9871 10195 9877
rect 13354 9868 13360 9880
rect 13412 9868 13418 9920
rect 1104 9818 21804 9840
rect 1104 9766 4432 9818
rect 4484 9766 4496 9818
rect 4548 9766 4560 9818
rect 4612 9766 4624 9818
rect 4676 9766 11332 9818
rect 11384 9766 11396 9818
rect 11448 9766 11460 9818
rect 11512 9766 11524 9818
rect 11576 9766 18232 9818
rect 18284 9766 18296 9818
rect 18348 9766 18360 9818
rect 18412 9766 18424 9818
rect 18476 9766 21804 9818
rect 1104 9744 21804 9766
rect 2222 9664 2228 9716
rect 2280 9704 2286 9716
rect 2317 9707 2375 9713
rect 2317 9704 2329 9707
rect 2280 9676 2329 9704
rect 2280 9664 2286 9676
rect 2317 9673 2329 9676
rect 2363 9673 2375 9707
rect 2317 9667 2375 9673
rect 13173 9707 13231 9713
rect 13173 9673 13185 9707
rect 13219 9704 13231 9707
rect 13446 9704 13452 9716
rect 13219 9676 13452 9704
rect 13219 9673 13231 9676
rect 13173 9667 13231 9673
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 2774 9596 2780 9648
rect 2832 9636 2838 9648
rect 5261 9639 5319 9645
rect 2832 9608 2877 9636
rect 2832 9596 2838 9608
rect 5261 9605 5273 9639
rect 5307 9636 5319 9639
rect 11146 9636 11152 9648
rect 5307 9608 11152 9636
rect 5307 9605 5319 9608
rect 5261 9599 5319 9605
rect 11146 9596 11152 9608
rect 11204 9596 11210 9648
rect 7190 9528 7196 9580
rect 7248 9568 7254 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 7248 9540 7389 9568
rect 7248 9528 7254 9540
rect 7377 9537 7389 9540
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 9585 9571 9643 9577
rect 9585 9537 9597 9571
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 9677 9571 9735 9577
rect 9677 9537 9689 9571
rect 9723 9568 9735 9571
rect 10502 9568 10508 9580
rect 9723 9540 10508 9568
rect 9723 9537 9735 9540
rect 9677 9531 9735 9537
rect 1578 9460 1584 9512
rect 1636 9500 1642 9512
rect 1765 9503 1823 9509
rect 1765 9500 1777 9503
rect 1636 9472 1777 9500
rect 1636 9460 1642 9472
rect 1765 9469 1777 9472
rect 1811 9469 1823 9503
rect 1765 9463 1823 9469
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9500 2375 9503
rect 2866 9500 2872 9512
rect 2363 9472 2872 9500
rect 2363 9469 2375 9472
rect 2317 9463 2375 9469
rect 2866 9460 2872 9472
rect 2924 9500 2930 9512
rect 2961 9503 3019 9509
rect 2961 9500 2973 9503
rect 2924 9472 2973 9500
rect 2924 9460 2930 9472
rect 2961 9469 2973 9472
rect 3007 9469 3019 9503
rect 4982 9500 4988 9512
rect 4943 9472 4988 9500
rect 2961 9463 3019 9469
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 7558 9500 7564 9512
rect 7519 9472 7564 9500
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 8297 9503 8355 9509
rect 8297 9469 8309 9503
rect 8343 9500 8355 9503
rect 8478 9500 8484 9512
rect 8343 9472 8484 9500
rect 8343 9469 8355 9472
rect 8297 9463 8355 9469
rect 2406 9392 2412 9444
rect 2464 9432 2470 9444
rect 4709 9435 4767 9441
rect 4709 9432 4721 9435
rect 2464 9404 4721 9432
rect 2464 9392 2470 9404
rect 4709 9401 4721 9404
rect 4755 9432 4767 9435
rect 5166 9432 5172 9444
rect 4755 9404 5172 9432
rect 4755 9401 4767 9404
rect 4709 9395 4767 9401
rect 5166 9392 5172 9404
rect 5224 9432 5230 9444
rect 5442 9432 5448 9444
rect 5224 9404 5448 9432
rect 5224 9392 5230 9404
rect 5442 9392 5448 9404
rect 5500 9432 5506 9444
rect 8312 9432 8340 9463
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 9600 9500 9628 9531
rect 10502 9528 10508 9540
rect 10560 9528 10566 9580
rect 11164 9500 11192 9596
rect 12434 9528 12440 9580
rect 12492 9568 12498 9580
rect 12492 9540 13124 9568
rect 12492 9528 12498 9540
rect 12069 9503 12127 9509
rect 12069 9500 12081 9503
rect 9600 9472 9720 9500
rect 11164 9472 12081 9500
rect 9692 9444 9720 9472
rect 12069 9469 12081 9472
rect 12115 9469 12127 9503
rect 12069 9463 12127 9469
rect 12621 9503 12679 9509
rect 12621 9469 12633 9503
rect 12667 9500 12679 9503
rect 12986 9500 12992 9512
rect 12667 9472 12992 9500
rect 12667 9469 12679 9472
rect 12621 9463 12679 9469
rect 12986 9460 12992 9472
rect 13044 9460 13050 9512
rect 13096 9509 13124 9540
rect 13081 9503 13139 9509
rect 13081 9469 13093 9503
rect 13127 9469 13139 9503
rect 14274 9500 14280 9512
rect 14235 9472 14280 9500
rect 13081 9463 13139 9469
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 9674 9432 9680 9444
rect 5500 9404 8340 9432
rect 9587 9404 9680 9432
rect 5500 9392 5506 9404
rect 9674 9392 9680 9404
rect 9732 9432 9738 9444
rect 12342 9432 12348 9444
rect 9732 9404 12348 9432
rect 9732 9392 9738 9404
rect 12342 9392 12348 9404
rect 12400 9392 12406 9444
rect 4798 9364 4804 9376
rect 4759 9336 4804 9364
rect 4798 9324 4804 9336
rect 4856 9324 4862 9376
rect 9769 9367 9827 9373
rect 9769 9333 9781 9367
rect 9815 9364 9827 9367
rect 9950 9364 9956 9376
rect 9815 9336 9956 9364
rect 9815 9333 9827 9336
rect 9769 9327 9827 9333
rect 9950 9324 9956 9336
rect 10008 9324 10014 9376
rect 10134 9364 10140 9376
rect 10095 9336 10140 9364
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 14461 9367 14519 9373
rect 14461 9333 14473 9367
rect 14507 9364 14519 9367
rect 15194 9364 15200 9376
rect 14507 9336 15200 9364
rect 14507 9333 14519 9336
rect 14461 9327 14519 9333
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 1104 9274 21804 9296
rect 1104 9222 7882 9274
rect 7934 9222 7946 9274
rect 7998 9222 8010 9274
rect 8062 9222 8074 9274
rect 8126 9222 14782 9274
rect 14834 9222 14846 9274
rect 14898 9222 14910 9274
rect 14962 9222 14974 9274
rect 15026 9222 21804 9274
rect 1104 9200 21804 9222
rect 2222 9120 2228 9172
rect 2280 9160 2286 9172
rect 2685 9163 2743 9169
rect 2685 9160 2697 9163
rect 2280 9132 2697 9160
rect 2280 9120 2286 9132
rect 2685 9129 2697 9132
rect 2731 9129 2743 9163
rect 9950 9160 9956 9172
rect 2685 9123 2743 9129
rect 4908 9132 7052 9160
rect 9911 9132 9956 9160
rect 1394 9052 1400 9104
rect 1452 9092 1458 9104
rect 4908 9092 4936 9132
rect 1452 9064 4936 9092
rect 1452 9052 1458 9064
rect 5534 9052 5540 9104
rect 5592 9052 5598 9104
rect 5810 9092 5816 9104
rect 5771 9064 5816 9092
rect 5810 9052 5816 9064
rect 5868 9052 5874 9104
rect 5994 9092 6000 9104
rect 5955 9064 6000 9092
rect 5994 9052 6000 9064
rect 6052 9052 6058 9104
rect 4709 9027 4767 9033
rect 4709 8993 4721 9027
rect 4755 8993 4767 9027
rect 4709 8987 4767 8993
rect 4893 9027 4951 9033
rect 4893 8993 4905 9027
rect 4939 8993 4951 9027
rect 4893 8987 4951 8993
rect 2498 8848 2504 8900
rect 2556 8888 2562 8900
rect 4525 8891 4583 8897
rect 4525 8888 4537 8891
rect 2556 8860 4537 8888
rect 2556 8848 2562 8860
rect 4525 8857 4537 8860
rect 4571 8857 4583 8891
rect 4724 8888 4752 8987
rect 4908 8956 4936 8987
rect 4982 8984 4988 9036
rect 5040 9024 5046 9036
rect 5040 8996 5085 9024
rect 5040 8984 5046 8996
rect 5552 8956 5580 9052
rect 6825 9027 6883 9033
rect 6825 8993 6837 9027
rect 6871 9024 6883 9027
rect 6914 9024 6920 9036
rect 6871 8996 6920 9024
rect 6871 8993 6883 8996
rect 6825 8987 6883 8993
rect 6914 8984 6920 8996
rect 6972 8984 6978 9036
rect 7024 9033 7052 9132
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 11882 9120 11888 9172
rect 11940 9160 11946 9172
rect 12161 9163 12219 9169
rect 12161 9160 12173 9163
rect 11940 9132 12173 9160
rect 11940 9120 11946 9132
rect 12161 9129 12173 9132
rect 12207 9129 12219 9163
rect 15194 9160 15200 9172
rect 15155 9132 15200 9160
rect 12161 9123 12219 9129
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 15286 9120 15292 9172
rect 15344 9160 15350 9172
rect 18598 9160 18604 9172
rect 15344 9132 15389 9160
rect 18559 9132 18604 9160
rect 15344 9120 15350 9132
rect 18598 9120 18604 9132
rect 18656 9120 18662 9172
rect 17310 9092 17316 9104
rect 17271 9064 17316 9092
rect 17310 9052 17316 9064
rect 17368 9052 17374 9104
rect 7009 9027 7067 9033
rect 7009 8993 7021 9027
rect 7055 8993 7067 9027
rect 7009 8987 7067 8993
rect 8113 9027 8171 9033
rect 8113 8993 8125 9027
rect 8159 9024 8171 9027
rect 8386 9024 8392 9036
rect 8159 8996 8392 9024
rect 8159 8993 8171 8996
rect 8113 8987 8171 8993
rect 8386 8984 8392 8996
rect 8444 8984 8450 9036
rect 9582 9024 9588 9036
rect 9543 8996 9588 9024
rect 9582 8984 9588 8996
rect 9640 8984 9646 9036
rect 9769 9027 9827 9033
rect 9769 8993 9781 9027
rect 9815 9024 9827 9027
rect 10042 9024 10048 9036
rect 9815 8996 10048 9024
rect 9815 8993 9827 8996
rect 9769 8987 9827 8993
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 10686 8984 10692 9036
rect 10744 9024 10750 9036
rect 11517 9027 11575 9033
rect 11517 9024 11529 9027
rect 10744 8996 11529 9024
rect 10744 8984 10750 8996
rect 11517 8993 11529 8996
rect 11563 8993 11575 9027
rect 11517 8987 11575 8993
rect 11701 9027 11759 9033
rect 11701 8993 11713 9027
rect 11747 9024 11759 9027
rect 12345 9027 12403 9033
rect 12345 9024 12357 9027
rect 11747 8996 12357 9024
rect 11747 8993 11759 8996
rect 11701 8987 11759 8993
rect 12345 8993 12357 8996
rect 12391 9024 12403 9027
rect 12986 9024 12992 9036
rect 12391 8996 12992 9024
rect 12391 8993 12403 8996
rect 12345 8987 12403 8993
rect 12986 8984 12992 8996
rect 13044 8984 13050 9036
rect 14458 8984 14464 9036
rect 14516 9024 14522 9036
rect 16209 9027 16267 9033
rect 16209 9024 16221 9027
rect 14516 8996 16221 9024
rect 14516 8984 14522 8996
rect 16209 8993 16221 8996
rect 16255 8993 16267 9027
rect 16209 8987 16267 8993
rect 16761 9027 16819 9033
rect 16761 8993 16773 9027
rect 16807 9024 16819 9027
rect 17497 9027 17555 9033
rect 17497 9024 17509 9027
rect 16807 8996 17509 9024
rect 16807 8993 16819 8996
rect 16761 8987 16819 8993
rect 17497 8993 17509 8996
rect 17543 8993 17555 9027
rect 17497 8987 17555 8993
rect 4908 8928 5580 8956
rect 5718 8916 5724 8968
rect 5776 8956 5782 8968
rect 7377 8959 7435 8965
rect 5776 8928 5821 8956
rect 5776 8916 5782 8928
rect 7377 8925 7389 8959
rect 7423 8956 7435 8959
rect 7558 8956 7564 8968
rect 7423 8928 7564 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 9493 8959 9551 8965
rect 9493 8925 9505 8959
rect 9539 8956 9551 8959
rect 9539 8928 9812 8956
rect 9539 8925 9551 8928
rect 9493 8919 9551 8925
rect 9784 8900 9812 8928
rect 12618 8916 12624 8968
rect 12676 8956 12682 8968
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 12676 8928 15393 8956
rect 12676 8916 12682 8928
rect 15381 8925 15393 8928
rect 15427 8925 15439 8959
rect 16574 8956 16580 8968
rect 16535 8928 16580 8956
rect 15381 8919 15439 8925
rect 16574 8916 16580 8928
rect 16632 8916 16638 8968
rect 17512 8956 17540 8987
rect 18046 8984 18052 9036
rect 18104 9024 18110 9036
rect 18233 9027 18291 9033
rect 18233 9024 18245 9027
rect 18104 8996 18245 9024
rect 18104 8984 18110 8996
rect 18233 8993 18245 8996
rect 18279 8993 18291 9027
rect 18233 8987 18291 8993
rect 18690 8956 18696 8968
rect 17512 8928 18696 8956
rect 18690 8916 18696 8928
rect 18748 8916 18754 8968
rect 7650 8888 7656 8900
rect 4724 8860 7656 8888
rect 4525 8851 4583 8857
rect 7650 8848 7656 8860
rect 7708 8848 7714 8900
rect 9766 8848 9772 8900
rect 9824 8848 9830 8900
rect 18601 8891 18659 8897
rect 18601 8857 18613 8891
rect 18647 8888 18659 8891
rect 19150 8888 19156 8900
rect 18647 8860 19156 8888
rect 18647 8857 18659 8860
rect 18601 8851 18659 8857
rect 19150 8848 19156 8860
rect 19208 8848 19214 8900
rect 2777 8823 2835 8829
rect 2777 8789 2789 8823
rect 2823 8820 2835 8823
rect 3878 8820 3884 8832
rect 2823 8792 3884 8820
rect 2823 8789 2835 8792
rect 2777 8783 2835 8789
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 6270 8820 6276 8832
rect 6231 8792 6276 8820
rect 6270 8780 6276 8792
rect 6328 8780 6334 8832
rect 7742 8780 7748 8832
rect 7800 8820 7806 8832
rect 7929 8823 7987 8829
rect 7929 8820 7941 8823
rect 7800 8792 7941 8820
rect 7800 8780 7806 8792
rect 7929 8789 7941 8792
rect 7975 8789 7987 8823
rect 7929 8783 7987 8789
rect 14642 8780 14648 8832
rect 14700 8820 14706 8832
rect 14829 8823 14887 8829
rect 14829 8820 14841 8823
rect 14700 8792 14841 8820
rect 14700 8780 14706 8792
rect 14829 8789 14841 8792
rect 14875 8789 14887 8823
rect 14829 8783 14887 8789
rect 1104 8730 21804 8752
rect 1104 8678 4432 8730
rect 4484 8678 4496 8730
rect 4548 8678 4560 8730
rect 4612 8678 4624 8730
rect 4676 8678 11332 8730
rect 11384 8678 11396 8730
rect 11448 8678 11460 8730
rect 11512 8678 11524 8730
rect 11576 8678 18232 8730
rect 18284 8678 18296 8730
rect 18348 8678 18360 8730
rect 18412 8678 18424 8730
rect 18476 8678 21804 8730
rect 1104 8656 21804 8678
rect 2130 8616 2136 8628
rect 2043 8588 2136 8616
rect 2130 8576 2136 8588
rect 2188 8616 2194 8628
rect 2188 8588 3372 8616
rect 2188 8576 2194 8588
rect 1581 8551 1639 8557
rect 1581 8517 1593 8551
rect 1627 8548 1639 8551
rect 1627 8520 2636 8548
rect 1627 8517 1639 8520
rect 1581 8511 1639 8517
rect 2608 8489 2636 8520
rect 3344 8489 3372 8588
rect 4982 8576 4988 8628
rect 5040 8616 5046 8628
rect 9401 8619 9459 8625
rect 9401 8616 9413 8619
rect 5040 8588 9413 8616
rect 5040 8576 5046 8588
rect 9401 8585 9413 8588
rect 9447 8585 9459 8619
rect 9582 8616 9588 8628
rect 9543 8588 9588 8616
rect 9401 8579 9459 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 16574 8576 16580 8628
rect 16632 8616 16638 8628
rect 17681 8619 17739 8625
rect 17681 8616 17693 8619
rect 16632 8588 17693 8616
rect 16632 8576 16638 8588
rect 17681 8585 17693 8588
rect 17727 8585 17739 8619
rect 17681 8579 17739 8585
rect 18598 8576 18604 8628
rect 18656 8616 18662 8628
rect 18693 8619 18751 8625
rect 18693 8616 18705 8619
rect 18656 8588 18705 8616
rect 18656 8576 18662 8588
rect 18693 8585 18705 8588
rect 18739 8585 18751 8619
rect 19150 8616 19156 8628
rect 19111 8588 19156 8616
rect 18693 8579 18751 8585
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 6270 8508 6276 8560
rect 6328 8548 6334 8560
rect 14458 8548 14464 8560
rect 6328 8520 14464 8548
rect 6328 8508 6334 8520
rect 14458 8508 14464 8520
rect 14516 8508 14522 8560
rect 14553 8551 14611 8557
rect 14553 8517 14565 8551
rect 14599 8548 14611 8551
rect 15013 8551 15071 8557
rect 15013 8548 15025 8551
rect 14599 8520 15025 8548
rect 14599 8517 14611 8520
rect 14553 8511 14611 8517
rect 15013 8517 15025 8520
rect 15059 8517 15071 8551
rect 15013 8511 15071 8517
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8449 2651 8483
rect 2593 8443 2651 8449
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 3329 8483 3387 8489
rect 3329 8449 3341 8483
rect 3375 8449 3387 8483
rect 3878 8480 3884 8492
rect 3839 8452 3884 8480
rect 3329 8443 3387 8449
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 2498 8412 2504 8424
rect 2459 8384 2504 8412
rect 2498 8372 2504 8384
rect 2556 8372 2562 8424
rect 2406 8304 2412 8356
rect 2464 8344 2470 8356
rect 2700 8344 2728 8443
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8480 7159 8483
rect 9401 8483 9459 8489
rect 7147 8452 8340 8480
rect 7147 8449 7159 8452
rect 7101 8443 7159 8449
rect 7558 8412 7564 8424
rect 7519 8384 7564 8412
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 8312 8421 8340 8452
rect 9401 8449 9413 8483
rect 9447 8480 9459 8483
rect 9585 8483 9643 8489
rect 9585 8480 9597 8483
rect 9447 8452 9597 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 9585 8449 9597 8452
rect 9631 8480 9643 8483
rect 9766 8480 9772 8492
rect 9631 8452 9772 8480
rect 9631 8449 9643 8452
rect 9585 8443 9643 8449
rect 9766 8440 9772 8452
rect 9824 8480 9830 8492
rect 14182 8480 14188 8492
rect 9824 8452 12112 8480
rect 14143 8452 14188 8480
rect 9824 8440 9830 8452
rect 8297 8415 8355 8421
rect 8297 8381 8309 8415
rect 8343 8381 8355 8415
rect 8297 8375 8355 8381
rect 9493 8415 9551 8421
rect 9493 8381 9505 8415
rect 9539 8412 9551 8415
rect 10042 8412 10048 8424
rect 9539 8384 10048 8412
rect 9539 8381 9551 8384
rect 9493 8375 9551 8381
rect 10042 8372 10048 8384
rect 10100 8372 10106 8424
rect 12084 8421 12112 8452
rect 14182 8440 14188 8452
rect 14240 8440 14246 8492
rect 14476 8480 14504 8508
rect 17313 8483 17371 8489
rect 17313 8480 17325 8483
rect 14476 8452 17325 8480
rect 17313 8449 17325 8452
rect 17359 8449 17371 8483
rect 17313 8443 17371 8449
rect 12069 8415 12127 8421
rect 12069 8381 12081 8415
rect 12115 8381 12127 8415
rect 14274 8412 14280 8424
rect 12069 8375 12127 8381
rect 12268 8384 14280 8412
rect 3786 8344 3792 8356
rect 2464 8316 2728 8344
rect 3747 8316 3792 8344
rect 2464 8304 2470 8316
rect 3786 8304 3792 8316
rect 3844 8304 3850 8356
rect 8205 8347 8263 8353
rect 8205 8313 8217 8347
rect 8251 8344 8263 8347
rect 8386 8344 8392 8356
rect 8251 8316 8392 8344
rect 8251 8313 8263 8316
rect 8205 8307 8263 8313
rect 8386 8304 8392 8316
rect 8444 8344 8450 8356
rect 9214 8344 9220 8356
rect 8444 8316 9220 8344
rect 8444 8304 8450 8316
rect 9214 8304 9220 8316
rect 9272 8304 9278 8356
rect 10060 8344 10088 8372
rect 12268 8353 12296 8384
rect 14274 8372 14280 8384
rect 14332 8372 14338 8424
rect 15197 8415 15255 8421
rect 15197 8381 15209 8415
rect 15243 8412 15255 8415
rect 15286 8412 15292 8424
rect 15243 8384 15292 8412
rect 15243 8381 15255 8384
rect 15197 8375 15255 8381
rect 15286 8372 15292 8384
rect 15344 8372 15350 8424
rect 17681 8415 17739 8421
rect 17681 8381 17693 8415
rect 17727 8412 17739 8415
rect 18046 8412 18052 8424
rect 17727 8384 18052 8412
rect 17727 8381 17739 8384
rect 17681 8375 17739 8381
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 18138 8372 18144 8424
rect 18196 8412 18202 8424
rect 18690 8412 18696 8424
rect 18196 8384 18241 8412
rect 18651 8384 18696 8412
rect 18196 8372 18202 8384
rect 18690 8372 18696 8384
rect 18748 8412 18754 8424
rect 19337 8415 19395 8421
rect 19337 8412 19349 8415
rect 18748 8384 19349 8412
rect 18748 8372 18754 8384
rect 19337 8381 19349 8384
rect 19383 8381 19395 8415
rect 21082 8412 21088 8424
rect 21043 8384 21088 8412
rect 19337 8375 19395 8381
rect 21082 8372 21088 8384
rect 21140 8372 21146 8424
rect 12253 8347 12311 8353
rect 12253 8344 12265 8347
rect 10060 8316 12265 8344
rect 12253 8313 12265 8316
rect 12299 8313 12311 8347
rect 12253 8307 12311 8313
rect 12342 8304 12348 8356
rect 12400 8344 12406 8356
rect 12618 8344 12624 8356
rect 12400 8316 12624 8344
rect 12400 8304 12406 8316
rect 12618 8304 12624 8316
rect 12676 8304 12682 8356
rect 9858 8276 9864 8288
rect 9819 8248 9864 8276
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 12434 8236 12440 8288
rect 12492 8276 12498 8288
rect 14550 8276 14556 8288
rect 12492 8248 12537 8276
rect 14511 8248 14556 8276
rect 12492 8236 12498 8248
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 20898 8276 20904 8288
rect 20859 8248 20904 8276
rect 20898 8236 20904 8248
rect 20956 8236 20962 8288
rect 1104 8186 21804 8208
rect 1104 8134 7882 8186
rect 7934 8134 7946 8186
rect 7998 8134 8010 8186
rect 8062 8134 8074 8186
rect 8126 8134 14782 8186
rect 14834 8134 14846 8186
rect 14898 8134 14910 8186
rect 14962 8134 14974 8186
rect 15026 8134 21804 8186
rect 1104 8112 21804 8134
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12805 8075 12863 8081
rect 12805 8072 12817 8075
rect 12492 8044 12817 8072
rect 12492 8032 12498 8044
rect 12805 8041 12817 8044
rect 12851 8041 12863 8075
rect 12805 8035 12863 8041
rect 18417 8075 18475 8081
rect 18417 8041 18429 8075
rect 18463 8072 18475 8075
rect 18598 8072 18604 8084
rect 18463 8044 18604 8072
rect 18463 8041 18475 8044
rect 18417 8035 18475 8041
rect 18598 8032 18604 8044
rect 18656 8032 18662 8084
rect 8021 8007 8079 8013
rect 8021 7973 8033 8007
rect 8067 8004 8079 8007
rect 8294 8004 8300 8016
rect 8067 7976 8300 8004
rect 8067 7973 8079 7976
rect 8021 7967 8079 7973
rect 8294 7964 8300 7976
rect 8352 7964 8358 8016
rect 14550 7964 14556 8016
rect 14608 8004 14614 8016
rect 15197 8007 15255 8013
rect 15197 8004 15209 8007
rect 14608 7976 15209 8004
rect 14608 7964 14614 7976
rect 15197 7973 15209 7976
rect 15243 7973 15255 8007
rect 15197 7967 15255 7973
rect 16393 8007 16451 8013
rect 16393 7973 16405 8007
rect 16439 8004 16451 8007
rect 16574 8004 16580 8016
rect 16439 7976 16580 8004
rect 16439 7973 16451 7976
rect 16393 7967 16451 7973
rect 16574 7964 16580 7976
rect 16632 7964 16638 8016
rect 18046 7964 18052 8016
rect 18104 8004 18110 8016
rect 18233 8007 18291 8013
rect 18233 8004 18245 8007
rect 18104 7976 18245 8004
rect 18104 7964 18110 7976
rect 18233 7973 18245 7976
rect 18279 7973 18291 8007
rect 18233 7967 18291 7973
rect 2130 7936 2136 7948
rect 2091 7908 2136 7936
rect 2130 7896 2136 7908
rect 2188 7896 2194 7948
rect 2682 7936 2688 7948
rect 2643 7908 2688 7936
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 7742 7936 7748 7948
rect 7703 7908 7748 7936
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 9861 7939 9919 7945
rect 9861 7905 9873 7939
rect 9907 7936 9919 7939
rect 10318 7936 10324 7948
rect 9907 7908 10324 7936
rect 9907 7905 9919 7908
rect 9861 7899 9919 7905
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 14182 7896 14188 7948
rect 14240 7936 14246 7948
rect 14737 7939 14795 7945
rect 14737 7936 14749 7939
rect 14240 7908 14749 7936
rect 14240 7896 14246 7908
rect 14737 7905 14749 7908
rect 14783 7905 14795 7939
rect 15286 7936 15292 7948
rect 15247 7908 15292 7936
rect 14737 7899 14795 7905
rect 15286 7896 15292 7908
rect 15344 7936 15350 7948
rect 16209 7939 16267 7945
rect 16209 7936 16221 7939
rect 15344 7908 16221 7936
rect 15344 7896 15350 7908
rect 16209 7905 16221 7908
rect 16255 7905 16267 7939
rect 16209 7899 16267 7905
rect 12618 7868 12624 7880
rect 12579 7840 12624 7868
rect 12618 7828 12624 7840
rect 12676 7828 12682 7880
rect 12713 7871 12771 7877
rect 12713 7837 12725 7871
rect 12759 7868 12771 7871
rect 20898 7868 20904 7880
rect 12759 7840 20904 7868
rect 12759 7837 12771 7840
rect 12713 7831 12771 7837
rect 20898 7828 20904 7840
rect 20956 7828 20962 7880
rect 2685 7735 2743 7741
rect 2685 7701 2697 7735
rect 2731 7732 2743 7735
rect 3786 7732 3792 7744
rect 2731 7704 3792 7732
rect 2731 7701 2743 7704
rect 2685 7695 2743 7701
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 9490 7692 9496 7744
rect 9548 7732 9554 7744
rect 9769 7735 9827 7741
rect 9769 7732 9781 7735
rect 9548 7704 9781 7732
rect 9548 7692 9554 7704
rect 9769 7701 9781 7704
rect 9815 7701 9827 7735
rect 9769 7695 9827 7701
rect 13173 7735 13231 7741
rect 13173 7701 13185 7735
rect 13219 7732 13231 7735
rect 13262 7732 13268 7744
rect 13219 7704 13268 7732
rect 13219 7701 13231 7704
rect 13173 7695 13231 7701
rect 13262 7692 13268 7704
rect 13320 7692 13326 7744
rect 1104 7642 21804 7664
rect 1104 7590 4432 7642
rect 4484 7590 4496 7642
rect 4548 7590 4560 7642
rect 4612 7590 4624 7642
rect 4676 7590 11332 7642
rect 11384 7590 11396 7642
rect 11448 7590 11460 7642
rect 11512 7590 11524 7642
rect 11576 7590 18232 7642
rect 18284 7590 18296 7642
rect 18348 7590 18360 7642
rect 18412 7590 18424 7642
rect 18476 7590 21804 7642
rect 1104 7568 21804 7590
rect 3789 7531 3847 7537
rect 3789 7497 3801 7531
rect 3835 7528 3847 7531
rect 4062 7528 4068 7540
rect 3835 7500 4068 7528
rect 3835 7497 3847 7500
rect 3789 7491 3847 7497
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 12805 7531 12863 7537
rect 12805 7497 12817 7531
rect 12851 7528 12863 7531
rect 13446 7528 13452 7540
rect 12851 7500 13452 7528
rect 12851 7497 12863 7500
rect 12805 7491 12863 7497
rect 13446 7488 13452 7500
rect 13504 7528 13510 7540
rect 13633 7531 13691 7537
rect 13633 7528 13645 7531
rect 13504 7500 13645 7528
rect 13504 7488 13510 7500
rect 13633 7497 13645 7500
rect 13679 7497 13691 7531
rect 13633 7491 13691 7497
rect 4246 7352 4252 7404
rect 4304 7392 4310 7404
rect 4709 7395 4767 7401
rect 4709 7392 4721 7395
rect 4304 7364 4721 7392
rect 4304 7352 4310 7364
rect 4709 7361 4721 7364
rect 4755 7392 4767 7395
rect 5074 7392 5080 7404
rect 4755 7364 5080 7392
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 5074 7352 5080 7364
rect 5132 7352 5138 7404
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7392 8171 7395
rect 13262 7392 13268 7404
rect 8159 7364 9996 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 7742 7324 7748 7336
rect 7655 7296 7748 7324
rect 7742 7284 7748 7296
rect 7800 7324 7806 7336
rect 8573 7327 8631 7333
rect 8573 7324 8585 7327
rect 7800 7296 8585 7324
rect 7800 7284 7806 7296
rect 8573 7293 8585 7296
rect 8619 7293 8631 7327
rect 9490 7324 9496 7336
rect 9451 7296 9496 7324
rect 8573 7287 8631 7293
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 9968 7333 9996 7364
rect 12406 7364 13268 7392
rect 9953 7327 10011 7333
rect 9953 7293 9965 7327
rect 9999 7293 10011 7327
rect 10686 7324 10692 7336
rect 10647 7296 10692 7324
rect 9953 7287 10011 7293
rect 10686 7284 10692 7296
rect 10744 7284 10750 7336
rect 12253 7327 12311 7333
rect 12253 7293 12265 7327
rect 12299 7324 12311 7327
rect 12406 7324 12434 7364
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 15286 7392 15292 7404
rect 13556 7364 15292 7392
rect 12299 7296 12434 7324
rect 12805 7327 12863 7333
rect 12299 7293 12311 7296
rect 12253 7287 12311 7293
rect 12805 7293 12817 7327
rect 12851 7324 12863 7327
rect 13556 7324 13584 7364
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 12851 7296 13584 7324
rect 13633 7327 13691 7333
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 13633 7293 13645 7327
rect 13679 7324 13691 7327
rect 14093 7327 14151 7333
rect 14093 7324 14105 7327
rect 13679 7296 14105 7324
rect 13679 7293 13691 7296
rect 13633 7287 13691 7293
rect 14093 7293 14105 7296
rect 14139 7293 14151 7327
rect 14093 7287 14151 7293
rect 14277 7327 14335 7333
rect 14277 7293 14289 7327
rect 14323 7324 14335 7327
rect 14550 7324 14556 7336
rect 14323 7296 14556 7324
rect 14323 7293 14335 7296
rect 14277 7287 14335 7293
rect 14550 7284 14556 7296
rect 14608 7284 14614 7336
rect 3878 7256 3884 7268
rect 3839 7228 3884 7256
rect 3878 7216 3884 7228
rect 3936 7256 3942 7268
rect 5169 7259 5227 7265
rect 5169 7256 5181 7259
rect 3936 7228 5181 7256
rect 3936 7216 3942 7228
rect 5169 7225 5181 7228
rect 5215 7225 5227 7259
rect 5169 7219 5227 7225
rect 5261 7259 5319 7265
rect 5261 7225 5273 7259
rect 5307 7256 5319 7259
rect 5721 7259 5779 7265
rect 5721 7256 5733 7259
rect 5307 7228 5733 7256
rect 5307 7225 5319 7228
rect 5261 7219 5319 7225
rect 5721 7225 5733 7228
rect 5767 7225 5779 7259
rect 5721 7219 5779 7225
rect 7558 7216 7564 7268
rect 7616 7256 7622 7268
rect 7929 7259 7987 7265
rect 7929 7256 7941 7259
rect 7616 7228 7941 7256
rect 7616 7216 7622 7228
rect 7929 7225 7941 7228
rect 7975 7225 7987 7259
rect 9214 7256 9220 7268
rect 9127 7228 9220 7256
rect 7929 7219 7987 7225
rect 9214 7216 9220 7228
rect 9272 7256 9278 7268
rect 10704 7256 10732 7284
rect 9272 7228 10732 7256
rect 10873 7259 10931 7265
rect 9272 7216 9278 7228
rect 10873 7225 10885 7259
rect 10919 7256 10931 7259
rect 10962 7256 10968 7268
rect 10919 7228 10968 7256
rect 10919 7225 10931 7228
rect 10873 7219 10931 7225
rect 10962 7216 10968 7228
rect 11020 7216 11026 7268
rect 5902 7188 5908 7200
rect 5863 7160 5908 7188
rect 5902 7148 5908 7160
rect 5960 7148 5966 7200
rect 1104 7098 21804 7120
rect 1104 7046 7882 7098
rect 7934 7046 7946 7098
rect 7998 7046 8010 7098
rect 8062 7046 8074 7098
rect 8126 7046 14782 7098
rect 14834 7046 14846 7098
rect 14898 7046 14910 7098
rect 14962 7046 14974 7098
rect 15026 7046 21804 7098
rect 1104 7024 21804 7046
rect 7742 6944 7748 6996
rect 7800 6984 7806 6996
rect 7837 6987 7895 6993
rect 7837 6984 7849 6987
rect 7800 6956 7849 6984
rect 7800 6944 7806 6956
rect 7837 6953 7849 6956
rect 7883 6953 7895 6987
rect 10870 6984 10876 6996
rect 10831 6956 10876 6984
rect 7837 6947 7895 6953
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 17770 6984 17776 6996
rect 17731 6956 17776 6984
rect 17770 6944 17776 6956
rect 17828 6944 17834 6996
rect 3878 6876 3884 6928
rect 3936 6916 3942 6928
rect 4893 6919 4951 6925
rect 4893 6916 4905 6919
rect 3936 6888 4905 6916
rect 3936 6876 3942 6888
rect 4893 6885 4905 6888
rect 4939 6885 4951 6919
rect 4893 6879 4951 6885
rect 5721 6919 5779 6925
rect 5721 6885 5733 6919
rect 5767 6916 5779 6919
rect 5902 6916 5908 6928
rect 5767 6888 5908 6916
rect 5767 6885 5779 6888
rect 5721 6879 5779 6885
rect 5902 6876 5908 6888
rect 5960 6876 5966 6928
rect 7650 6876 7656 6928
rect 7708 6916 7714 6928
rect 8205 6919 8263 6925
rect 8205 6916 8217 6919
rect 7708 6888 8217 6916
rect 7708 6876 7714 6888
rect 8205 6885 8217 6888
rect 8251 6885 8263 6919
rect 10318 6916 10324 6928
rect 10279 6888 10324 6916
rect 8205 6879 8263 6885
rect 10318 6876 10324 6888
rect 10376 6876 10382 6928
rect 4246 6848 4252 6860
rect 4207 6820 4252 6848
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 5169 6851 5227 6857
rect 5169 6817 5181 6851
rect 5215 6848 5227 6851
rect 5626 6848 5632 6860
rect 5215 6820 5632 6848
rect 5215 6817 5227 6820
rect 5169 6811 5227 6817
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 6178 6848 6184 6860
rect 6139 6820 6184 6848
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 8297 6851 8355 6857
rect 8297 6817 8309 6851
rect 8343 6848 8355 6851
rect 9861 6851 9919 6857
rect 8343 6820 9674 6848
rect 8343 6817 8355 6820
rect 8297 6811 8355 6817
rect 8481 6783 8539 6789
rect 8481 6749 8493 6783
rect 8527 6749 8539 6783
rect 9646 6780 9674 6820
rect 9861 6817 9873 6851
rect 9907 6848 9919 6851
rect 10134 6848 10140 6860
rect 9907 6820 10140 6848
rect 9907 6817 9919 6820
rect 9861 6811 9919 6817
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 10413 6851 10471 6857
rect 10413 6817 10425 6851
rect 10459 6848 10471 6851
rect 10962 6848 10968 6860
rect 10459 6820 10968 6848
rect 10459 6817 10471 6820
rect 10413 6811 10471 6817
rect 10962 6808 10968 6820
rect 11020 6848 11026 6860
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 11020 6820 11069 6848
rect 11020 6808 11026 6820
rect 11057 6817 11069 6820
rect 11103 6817 11115 6851
rect 15930 6848 15936 6860
rect 15891 6820 15936 6848
rect 11057 6811 11115 6817
rect 15930 6808 15936 6820
rect 15988 6808 15994 6860
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6848 16083 6851
rect 17402 6848 17408 6860
rect 16071 6820 17408 6848
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 17773 6851 17831 6857
rect 17773 6817 17785 6851
rect 17819 6817 17831 6851
rect 17773 6811 17831 6817
rect 16206 6780 16212 6792
rect 9646 6752 11008 6780
rect 16167 6752 16212 6780
rect 8481 6743 8539 6749
rect 8496 6712 8524 6743
rect 9674 6712 9680 6724
rect 8496 6684 9680 6712
rect 9674 6672 9680 6684
rect 9732 6672 9738 6724
rect 10980 6712 11008 6752
rect 16206 6740 16212 6752
rect 16264 6740 16270 6792
rect 17494 6740 17500 6792
rect 17552 6780 17558 6792
rect 17589 6783 17647 6789
rect 17589 6780 17601 6783
rect 17552 6752 17601 6780
rect 17552 6740 17558 6752
rect 17589 6749 17601 6752
rect 17635 6749 17647 6783
rect 17788 6780 17816 6811
rect 17862 6808 17868 6860
rect 17920 6848 17926 6860
rect 17957 6851 18015 6857
rect 17957 6848 17969 6851
rect 17920 6820 17969 6848
rect 17920 6808 17926 6820
rect 17957 6817 17969 6820
rect 18003 6817 18015 6851
rect 17957 6811 18015 6817
rect 18690 6780 18696 6792
rect 17788 6752 18696 6780
rect 17589 6743 17647 6749
rect 18690 6740 18696 6752
rect 18748 6740 18754 6792
rect 20898 6712 20904 6724
rect 10980 6684 20904 6712
rect 20898 6672 20904 6684
rect 20956 6672 20962 6724
rect 2038 6604 2044 6656
rect 2096 6644 2102 6656
rect 15565 6647 15623 6653
rect 15565 6644 15577 6647
rect 2096 6616 15577 6644
rect 2096 6604 2102 6616
rect 15565 6613 15577 6616
rect 15611 6613 15623 6647
rect 15565 6607 15623 6613
rect 1104 6554 21804 6576
rect 1104 6502 4432 6554
rect 4484 6502 4496 6554
rect 4548 6502 4560 6554
rect 4612 6502 4624 6554
rect 4676 6502 11332 6554
rect 11384 6502 11396 6554
rect 11448 6502 11460 6554
rect 11512 6502 11524 6554
rect 11576 6502 18232 6554
rect 18284 6502 18296 6554
rect 18348 6502 18360 6554
rect 18412 6502 18424 6554
rect 18476 6502 21804 6554
rect 1104 6480 21804 6502
rect 5905 6375 5963 6381
rect 5905 6341 5917 6375
rect 5951 6372 5963 6375
rect 6825 6375 6883 6381
rect 6825 6372 6837 6375
rect 5951 6344 6837 6372
rect 5951 6341 5963 6344
rect 5905 6335 5963 6341
rect 6825 6341 6837 6344
rect 6871 6341 6883 6375
rect 6825 6335 6883 6341
rect 10229 6375 10287 6381
rect 10229 6341 10241 6375
rect 10275 6372 10287 6375
rect 10870 6372 10876 6384
rect 10275 6344 10876 6372
rect 10275 6341 10287 6344
rect 10229 6335 10287 6341
rect 10870 6332 10876 6344
rect 10928 6332 10934 6384
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6304 5595 6307
rect 6178 6304 6184 6316
rect 5583 6276 6184 6304
rect 5583 6273 5595 6276
rect 5537 6267 5595 6273
rect 6178 6264 6184 6276
rect 6236 6264 6242 6316
rect 9861 6307 9919 6313
rect 9861 6273 9873 6307
rect 9907 6304 9919 6307
rect 10134 6304 10140 6316
rect 9907 6276 10140 6304
rect 9907 6273 9919 6276
rect 9861 6267 9919 6273
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 14642 6304 14648 6316
rect 14603 6276 14648 6304
rect 14642 6264 14648 6276
rect 14700 6264 14706 6316
rect 16206 6264 16212 6316
rect 16264 6304 16270 6316
rect 17313 6307 17371 6313
rect 17313 6304 17325 6307
rect 16264 6276 17325 6304
rect 16264 6264 16270 6276
rect 17313 6273 17325 6276
rect 17359 6273 17371 6307
rect 17313 6267 17371 6273
rect 3478 6239 3536 6245
rect 3478 6205 3490 6239
rect 3524 6236 3536 6239
rect 3878 6236 3884 6248
rect 3524 6208 3884 6236
rect 3524 6205 3536 6208
rect 3478 6199 3536 6205
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 5626 6196 5632 6248
rect 5684 6236 5690 6248
rect 6822 6236 6828 6248
rect 5684 6208 6828 6236
rect 5684 6196 5690 6208
rect 6822 6196 6828 6208
rect 6880 6236 6886 6248
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 6880 6208 7021 6236
rect 6880 6196 6886 6208
rect 7009 6205 7021 6208
rect 7055 6205 7067 6239
rect 7009 6199 7067 6205
rect 15013 6239 15071 6245
rect 15013 6205 15025 6239
rect 15059 6236 15071 6239
rect 15102 6236 15108 6248
rect 15059 6208 15108 6236
rect 15059 6205 15071 6208
rect 15013 6199 15071 6205
rect 15102 6196 15108 6208
rect 15160 6196 15166 6248
rect 17494 6236 17500 6248
rect 17455 6208 17500 6236
rect 17494 6196 17500 6208
rect 17552 6196 17558 6248
rect 17678 6236 17684 6248
rect 17639 6208 17684 6236
rect 17678 6196 17684 6208
rect 17736 6196 17742 6248
rect 17862 6236 17868 6248
rect 17823 6208 17868 6236
rect 17862 6196 17868 6208
rect 17920 6236 17926 6248
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 17920 6208 18429 6236
rect 17920 6196 17926 6208
rect 18417 6205 18429 6208
rect 18463 6205 18475 6239
rect 18690 6236 18696 6248
rect 18651 6208 18696 6236
rect 18417 6199 18475 6205
rect 18690 6196 18696 6208
rect 18748 6196 18754 6248
rect 18874 6236 18880 6248
rect 18835 6208 18880 6236
rect 18874 6196 18880 6208
rect 18932 6196 18938 6248
rect 2774 6060 2780 6112
rect 2832 6100 2838 6112
rect 3375 6103 3433 6109
rect 3375 6100 3387 6103
rect 2832 6072 3387 6100
rect 2832 6060 2838 6072
rect 3375 6069 3387 6072
rect 3421 6069 3433 6103
rect 5902 6100 5908 6112
rect 5863 6072 5908 6100
rect 3375 6063 3433 6069
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 10229 6103 10287 6109
rect 10229 6069 10241 6103
rect 10275 6100 10287 6103
rect 10318 6100 10324 6112
rect 10275 6072 10324 6100
rect 10275 6069 10287 6072
rect 10229 6063 10287 6069
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 15013 6103 15071 6109
rect 15013 6069 15025 6103
rect 15059 6100 15071 6103
rect 15194 6100 15200 6112
rect 15059 6072 15200 6100
rect 15059 6069 15071 6072
rect 15013 6063 15071 6069
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 18598 6060 18604 6112
rect 18656 6100 18662 6112
rect 18693 6103 18751 6109
rect 18693 6100 18705 6103
rect 18656 6072 18705 6100
rect 18656 6060 18662 6072
rect 18693 6069 18705 6072
rect 18739 6069 18751 6103
rect 18693 6063 18751 6069
rect 1104 6010 21804 6032
rect 1104 5958 7882 6010
rect 7934 5958 7946 6010
rect 7998 5958 8010 6010
rect 8062 5958 8074 6010
rect 8126 5958 14782 6010
rect 14834 5958 14846 6010
rect 14898 5958 14910 6010
rect 14962 5958 14974 6010
rect 15026 5958 21804 6010
rect 1104 5936 21804 5958
rect 6822 5856 6828 5908
rect 6880 5896 6886 5908
rect 6917 5899 6975 5905
rect 6917 5896 6929 5899
rect 6880 5868 6929 5896
rect 6880 5856 6886 5868
rect 6917 5865 6929 5868
rect 6963 5865 6975 5899
rect 6917 5859 6975 5865
rect 15930 5856 15936 5908
rect 15988 5896 15994 5908
rect 16117 5899 16175 5905
rect 16117 5896 16129 5899
rect 15988 5868 16129 5896
rect 15988 5856 15994 5868
rect 16117 5865 16129 5868
rect 16163 5865 16175 5899
rect 16117 5859 16175 5865
rect 18601 5899 18659 5905
rect 18601 5865 18613 5899
rect 18647 5896 18659 5899
rect 18690 5896 18696 5908
rect 18647 5868 18696 5896
rect 18647 5865 18659 5868
rect 18601 5859 18659 5865
rect 18690 5856 18696 5868
rect 18748 5856 18754 5908
rect 20898 5896 20904 5908
rect 20859 5868 20904 5896
rect 20898 5856 20904 5868
rect 20956 5856 20962 5908
rect 1581 5831 1639 5837
rect 1581 5797 1593 5831
rect 1627 5828 1639 5831
rect 4982 5828 4988 5840
rect 1627 5800 4988 5828
rect 1627 5797 1639 5800
rect 1581 5791 1639 5797
rect 4982 5788 4988 5800
rect 5040 5788 5046 5840
rect 13446 5828 13452 5840
rect 13407 5800 13452 5828
rect 13446 5788 13452 5800
rect 13504 5788 13510 5840
rect 14826 5788 14832 5840
rect 14884 5828 14890 5840
rect 15194 5828 15200 5840
rect 14884 5800 15200 5828
rect 14884 5788 14890 5800
rect 15194 5788 15200 5800
rect 15252 5788 15258 5840
rect 17678 5788 17684 5840
rect 17736 5828 17742 5840
rect 17736 5800 18736 5828
rect 17736 5788 17742 5800
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 7009 5763 7067 5769
rect 2832 5732 2877 5760
rect 2832 5720 2838 5732
rect 7009 5729 7021 5763
rect 7055 5760 7067 5763
rect 8294 5760 8300 5772
rect 7055 5732 8300 5760
rect 7055 5729 7067 5732
rect 7009 5723 7067 5729
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 12710 5760 12716 5772
rect 12671 5732 12716 5760
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 14642 5720 14648 5772
rect 14700 5760 14706 5772
rect 14737 5763 14795 5769
rect 14737 5760 14749 5763
rect 14700 5732 14749 5760
rect 14700 5720 14706 5732
rect 14737 5729 14749 5732
rect 14783 5729 14795 5763
rect 15286 5760 15292 5772
rect 15247 5732 15292 5760
rect 14737 5723 14795 5729
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5760 16543 5763
rect 17310 5760 17316 5772
rect 16531 5732 17316 5760
rect 16531 5729 16543 5732
rect 16485 5723 16543 5729
rect 17310 5720 17316 5732
rect 17368 5720 17374 5772
rect 17788 5769 17816 5800
rect 17773 5763 17831 5769
rect 17773 5729 17785 5763
rect 17819 5729 17831 5763
rect 17773 5723 17831 5729
rect 17862 5720 17868 5772
rect 17920 5760 17926 5772
rect 18708 5769 18736 5800
rect 17957 5763 18015 5769
rect 17957 5760 17969 5763
rect 17920 5732 17969 5760
rect 17920 5720 17926 5732
rect 17957 5729 17969 5732
rect 18003 5729 18015 5763
rect 17957 5723 18015 5729
rect 18693 5763 18751 5769
rect 18693 5729 18705 5763
rect 18739 5760 18751 5763
rect 20806 5760 20812 5772
rect 18739 5732 20812 5760
rect 18739 5729 18751 5732
rect 18693 5723 18751 5729
rect 20806 5720 20812 5732
rect 20864 5720 20870 5772
rect 21082 5760 21088 5772
rect 21043 5732 21088 5760
rect 21082 5720 21088 5732
rect 21140 5720 21146 5772
rect 15194 5652 15200 5704
rect 15252 5692 15258 5704
rect 16577 5695 16635 5701
rect 16577 5692 16589 5695
rect 15252 5664 16589 5692
rect 15252 5652 15258 5664
rect 16577 5661 16589 5664
rect 16623 5661 16635 5695
rect 16577 5655 16635 5661
rect 16761 5695 16819 5701
rect 16761 5661 16773 5695
rect 16807 5692 16819 5695
rect 17405 5695 17463 5701
rect 17405 5692 17417 5695
rect 16807 5664 17417 5692
rect 16807 5661 16819 5664
rect 16761 5655 16819 5661
rect 17405 5661 17417 5664
rect 17451 5661 17463 5695
rect 17405 5655 17463 5661
rect 17589 5695 17647 5701
rect 17589 5661 17601 5695
rect 17635 5692 17647 5695
rect 18874 5692 18880 5704
rect 17635 5664 18880 5692
rect 17635 5661 17647 5664
rect 17589 5655 17647 5661
rect 18874 5652 18880 5664
rect 18932 5652 18938 5704
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 13265 5627 13323 5633
rect 13265 5624 13277 5627
rect 9732 5596 13277 5624
rect 9732 5584 9738 5596
rect 13265 5593 13277 5596
rect 13311 5593 13323 5627
rect 13265 5587 13323 5593
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 2682 5556 2688 5568
rect 2643 5528 2688 5556
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 12618 5556 12624 5568
rect 12579 5528 12624 5556
rect 12618 5516 12624 5528
rect 12676 5516 12682 5568
rect 1104 5466 21804 5488
rect 1104 5414 4432 5466
rect 4484 5414 4496 5466
rect 4548 5414 4560 5466
rect 4612 5414 4624 5466
rect 4676 5414 11332 5466
rect 11384 5414 11396 5466
rect 11448 5414 11460 5466
rect 11512 5414 11524 5466
rect 11576 5414 18232 5466
rect 18284 5414 18296 5466
rect 18348 5414 18360 5466
rect 18412 5414 18424 5466
rect 18476 5414 21804 5466
rect 1104 5392 21804 5414
rect 8113 5355 8171 5361
rect 8113 5321 8125 5355
rect 8159 5352 8171 5355
rect 8294 5352 8300 5364
rect 8159 5324 8300 5352
rect 8159 5321 8171 5324
rect 8113 5315 8171 5321
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 12710 5312 12716 5364
rect 12768 5352 12774 5364
rect 12989 5355 13047 5361
rect 12989 5352 13001 5355
rect 12768 5324 13001 5352
rect 12768 5312 12774 5324
rect 12989 5321 13001 5324
rect 13035 5352 13047 5355
rect 13817 5355 13875 5361
rect 13817 5352 13829 5355
rect 13035 5324 13829 5352
rect 13035 5321 13047 5324
rect 12989 5315 13047 5321
rect 13817 5321 13829 5324
rect 13863 5321 13875 5355
rect 15102 5352 15108 5364
rect 15063 5324 15108 5352
rect 13817 5315 13875 5321
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 17310 5352 17316 5364
rect 17271 5324 17316 5352
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 18601 5355 18659 5361
rect 18601 5321 18613 5355
rect 18647 5352 18659 5355
rect 18874 5352 18880 5364
rect 18647 5324 18880 5352
rect 18647 5321 18659 5324
rect 18601 5315 18659 5321
rect 18874 5312 18880 5324
rect 18932 5312 18938 5364
rect 15194 5284 15200 5296
rect 7024 5256 15200 5284
rect 3234 5216 3240 5228
rect 3195 5188 3240 5216
rect 3234 5176 3240 5188
rect 3292 5216 3298 5228
rect 3292 5188 5028 5216
rect 3292 5176 3298 5188
rect 2038 5108 2044 5160
rect 2096 5148 2102 5160
rect 2682 5148 2688 5160
rect 2096 5120 2688 5148
rect 2096 5108 2102 5120
rect 2682 5108 2688 5120
rect 2740 5148 2746 5160
rect 5000 5157 5028 5188
rect 7024 5160 7052 5256
rect 15194 5244 15200 5256
rect 15252 5244 15258 5296
rect 13449 5219 13507 5225
rect 13449 5216 13461 5219
rect 12452 5188 13461 5216
rect 2961 5151 3019 5157
rect 2961 5148 2973 5151
rect 2740 5120 2973 5148
rect 2740 5108 2746 5120
rect 2961 5117 2973 5120
rect 3007 5117 3019 5151
rect 2961 5111 3019 5117
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5148 5043 5151
rect 7006 5148 7012 5160
rect 5031 5120 7012 5148
rect 5031 5117 5043 5120
rect 4985 5111 5043 5117
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 7558 5148 7564 5160
rect 7519 5120 7564 5148
rect 7558 5108 7564 5120
rect 7616 5108 7622 5160
rect 8113 5151 8171 5157
rect 8113 5117 8125 5151
rect 8159 5148 8171 5151
rect 9674 5148 9680 5160
rect 8159 5120 9680 5148
rect 8159 5117 8171 5120
rect 8113 5111 8171 5117
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 10226 5148 10232 5160
rect 10187 5120 10232 5148
rect 10226 5108 10232 5120
rect 10284 5108 10290 5160
rect 11054 5108 11060 5160
rect 11112 5148 11118 5160
rect 12452 5157 12480 5188
rect 13449 5185 13461 5188
rect 13495 5185 13507 5219
rect 13449 5179 13507 5185
rect 17770 5176 17776 5228
rect 17828 5216 17834 5228
rect 17865 5219 17923 5225
rect 17865 5216 17877 5219
rect 17828 5188 17877 5216
rect 17828 5176 17834 5188
rect 17865 5185 17877 5188
rect 17911 5185 17923 5219
rect 17865 5179 17923 5185
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 11112 5120 12449 5148
rect 11112 5108 11118 5120
rect 12437 5117 12449 5120
rect 12483 5117 12495 5151
rect 12437 5111 12495 5117
rect 12989 5151 13047 5157
rect 12989 5117 13001 5151
rect 13035 5117 13047 5151
rect 12989 5111 13047 5117
rect 13817 5151 13875 5157
rect 13817 5117 13829 5151
rect 13863 5148 13875 5151
rect 14461 5151 14519 5157
rect 14461 5148 14473 5151
rect 13863 5120 14473 5148
rect 13863 5117 13875 5120
rect 13817 5111 13875 5117
rect 14461 5117 14473 5120
rect 14507 5117 14519 5151
rect 14461 5111 14519 5117
rect 14645 5151 14703 5157
rect 14645 5117 14657 5151
rect 14691 5148 14703 5151
rect 14826 5148 14832 5160
rect 14691 5120 14832 5148
rect 14691 5117 14703 5120
rect 14645 5111 14703 5117
rect 6270 5080 6276 5092
rect 4462 5052 6276 5080
rect 6270 5040 6276 5052
rect 6328 5040 6334 5092
rect 10962 5080 10968 5092
rect 10923 5052 10968 5080
rect 10962 5040 10968 5052
rect 11020 5040 11026 5092
rect 11149 5083 11207 5089
rect 11149 5049 11161 5083
rect 11195 5080 11207 5083
rect 12618 5080 12624 5092
rect 11195 5052 12624 5080
rect 11195 5049 11207 5052
rect 11149 5043 11207 5049
rect 12618 5040 12624 5052
rect 12676 5040 12682 5092
rect 13004 5080 13032 5111
rect 14826 5108 14832 5120
rect 14884 5108 14890 5160
rect 15286 5148 15292 5160
rect 15199 5120 15292 5148
rect 15286 5108 15292 5120
rect 15344 5108 15350 5160
rect 17494 5108 17500 5160
rect 17552 5148 17558 5160
rect 18509 5151 18567 5157
rect 18509 5148 18521 5151
rect 17552 5120 18521 5148
rect 17552 5108 17558 5120
rect 18509 5117 18521 5120
rect 18555 5117 18567 5151
rect 18509 5111 18567 5117
rect 15304 5080 15332 5108
rect 13004 5052 15332 5080
rect 17678 5012 17684 5024
rect 17639 4984 17684 5012
rect 17678 4972 17684 4984
rect 17736 4972 17742 5024
rect 17770 4972 17776 5024
rect 17828 5012 17834 5024
rect 17828 4984 17873 5012
rect 17828 4972 17834 4984
rect 1104 4922 21804 4944
rect 1104 4870 7882 4922
rect 7934 4870 7946 4922
rect 7998 4870 8010 4922
rect 8062 4870 8074 4922
rect 8126 4870 14782 4922
rect 14834 4870 14846 4922
rect 14898 4870 14910 4922
rect 14962 4870 14974 4922
rect 15026 4870 21804 4922
rect 1104 4848 21804 4870
rect 7558 4768 7564 4820
rect 7616 4808 7622 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7616 4780 7849 4808
rect 7616 4768 7622 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 7837 4771 7895 4777
rect 17678 4768 17684 4820
rect 17736 4808 17742 4820
rect 17957 4811 18015 4817
rect 17957 4808 17969 4811
rect 17736 4780 17969 4808
rect 17736 4768 17742 4780
rect 17957 4777 17969 4780
rect 18003 4777 18015 4811
rect 17957 4771 18015 4777
rect 18417 4811 18475 4817
rect 18417 4777 18429 4811
rect 18463 4808 18475 4811
rect 19610 4808 19616 4820
rect 18463 4780 19616 4808
rect 18463 4777 18475 4780
rect 18417 4771 18475 4777
rect 19610 4768 19616 4780
rect 19668 4808 19674 4820
rect 20714 4808 20720 4820
rect 19668 4780 20720 4808
rect 19668 4768 19674 4780
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 6270 4700 6276 4752
rect 6328 4740 6334 4752
rect 6730 4740 6736 4752
rect 6328 4712 6736 4740
rect 6328 4700 6334 4712
rect 6730 4700 6736 4712
rect 6788 4700 6794 4752
rect 7466 4700 7472 4752
rect 7524 4740 7530 4752
rect 8205 4743 8263 4749
rect 8205 4740 8217 4743
rect 7524 4712 8217 4740
rect 7524 4700 7530 4712
rect 8205 4709 8217 4712
rect 8251 4709 8263 4743
rect 8205 4703 8263 4709
rect 10962 4700 10968 4752
rect 11020 4740 11026 4752
rect 11149 4743 11207 4749
rect 11149 4740 11161 4743
rect 11020 4712 11161 4740
rect 11020 4700 11026 4712
rect 11149 4709 11161 4712
rect 11195 4709 11207 4743
rect 11149 4703 11207 4709
rect 4982 4672 4988 4684
rect 4895 4644 4988 4672
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 7006 4632 7012 4684
rect 7064 4672 7070 4684
rect 7064 4644 7109 4672
rect 7064 4632 7070 4644
rect 10226 4632 10232 4684
rect 10284 4672 10290 4684
rect 10505 4675 10563 4681
rect 10505 4672 10517 4675
rect 10284 4644 10517 4672
rect 10284 4632 10290 4644
rect 10505 4641 10517 4644
rect 10551 4641 10563 4675
rect 10505 4635 10563 4641
rect 11425 4675 11483 4681
rect 11425 4641 11437 4675
rect 11471 4672 11483 4675
rect 12158 4672 12164 4684
rect 11471 4644 12164 4672
rect 11471 4641 11483 4644
rect 11425 4635 11483 4641
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 18325 4675 18383 4681
rect 18325 4641 18337 4675
rect 18371 4672 18383 4675
rect 19426 4672 19432 4684
rect 18371 4644 19432 4672
rect 18371 4641 18383 4644
rect 18325 4635 18383 4641
rect 19426 4632 19432 4644
rect 19484 4632 19490 4684
rect 5000 4604 5028 4632
rect 6733 4607 6791 4613
rect 6733 4604 6745 4607
rect 5000 4576 6745 4604
rect 6733 4573 6745 4576
rect 6779 4604 6791 4607
rect 6779 4576 6960 4604
rect 6779 4573 6791 4576
rect 6733 4567 6791 4573
rect 6932 4536 6960 4576
rect 8202 4564 8208 4616
rect 8260 4604 8266 4616
rect 8297 4607 8355 4613
rect 8297 4604 8309 4607
rect 8260 4576 8309 4604
rect 8260 4564 8266 4576
rect 8297 4573 8309 4576
rect 8343 4573 8355 4607
rect 8478 4604 8484 4616
rect 8439 4576 8484 4604
rect 8297 4567 8355 4573
rect 8478 4564 8484 4576
rect 8536 4604 8542 4616
rect 9766 4604 9772 4616
rect 8536 4576 9772 4604
rect 8536 4564 8542 4576
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 18598 4604 18604 4616
rect 18559 4576 18604 4604
rect 18598 4564 18604 4576
rect 18656 4564 18662 4616
rect 6932 4508 12434 4536
rect 12406 4468 12434 4508
rect 17310 4468 17316 4480
rect 12406 4440 17316 4468
rect 17310 4428 17316 4440
rect 17368 4468 17374 4480
rect 17770 4468 17776 4480
rect 17368 4440 17776 4468
rect 17368 4428 17374 4440
rect 17770 4428 17776 4440
rect 17828 4428 17834 4480
rect 1104 4378 21804 4400
rect 1104 4326 4432 4378
rect 4484 4326 4496 4378
rect 4548 4326 4560 4378
rect 4612 4326 4624 4378
rect 4676 4326 11332 4378
rect 11384 4326 11396 4378
rect 11448 4326 11460 4378
rect 11512 4326 11524 4378
rect 11576 4326 18232 4378
rect 18284 4326 18296 4378
rect 18348 4326 18360 4378
rect 18412 4326 18424 4378
rect 18476 4326 21804 4378
rect 1104 4304 21804 4326
rect 8294 4264 8300 4276
rect 8255 4236 8300 4264
rect 8294 4224 8300 4236
rect 8352 4224 8358 4276
rect 12158 4264 12164 4276
rect 12119 4236 12164 4264
rect 12158 4224 12164 4236
rect 12216 4224 12222 4276
rect 18404 4267 18462 4273
rect 18404 4233 18416 4267
rect 18450 4264 18462 4267
rect 19426 4264 19432 4276
rect 18450 4236 19432 4264
rect 18450 4233 18462 4236
rect 18404 4227 18462 4233
rect 19426 4224 19432 4236
rect 19484 4264 19490 4276
rect 20162 4264 20168 4276
rect 19484 4236 20168 4264
rect 19484 4224 19490 4236
rect 20162 4224 20168 4236
rect 20220 4224 20226 4276
rect 15286 4156 15292 4208
rect 15344 4196 15350 4208
rect 15381 4199 15439 4205
rect 15381 4196 15393 4199
rect 15344 4168 15393 4196
rect 15344 4156 15350 4168
rect 15381 4165 15393 4168
rect 15427 4165 15439 4199
rect 15381 4159 15439 4165
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 7929 4131 7987 4137
rect 7929 4128 7941 4131
rect 7616 4100 7941 4128
rect 7616 4088 7622 4100
rect 7929 4097 7941 4100
rect 7975 4097 7987 4131
rect 7929 4091 7987 4097
rect 9585 4131 9643 4137
rect 9585 4097 9597 4131
rect 9631 4128 9643 4131
rect 9766 4128 9772 4140
rect 9631 4100 9772 4128
rect 9631 4097 9643 4100
rect 9585 4091 9643 4097
rect 9766 4088 9772 4100
rect 9824 4128 9830 4140
rect 10502 4128 10508 4140
rect 9824 4100 10508 4128
rect 9824 4088 9830 4100
rect 10502 4088 10508 4100
rect 10560 4088 10566 4140
rect 18141 4131 18199 4137
rect 18141 4097 18153 4131
rect 18187 4128 18199 4131
rect 19610 4128 19616 4140
rect 18187 4100 19616 4128
rect 18187 4097 18199 4100
rect 18141 4091 18199 4097
rect 19610 4088 19616 4100
rect 19668 4088 19674 4140
rect 8297 4063 8355 4069
rect 8297 4029 8309 4063
rect 8343 4060 8355 4063
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 8343 4032 8769 4060
rect 8343 4029 8355 4032
rect 8297 4023 8355 4029
rect 8757 4029 8769 4032
rect 8803 4029 8815 4063
rect 9858 4060 9864 4072
rect 9819 4032 9864 4060
rect 8757 4023 8815 4029
rect 9858 4020 9864 4032
rect 9916 4020 9922 4072
rect 1670 3952 1676 4004
rect 1728 3992 1734 4004
rect 11698 3992 11704 4004
rect 1728 3964 11704 3992
rect 1728 3952 1734 3964
rect 11698 3952 11704 3964
rect 11756 3952 11762 4004
rect 15562 3992 15568 4004
rect 15523 3964 15568 3992
rect 15562 3952 15568 3964
rect 15620 3952 15626 4004
rect 18046 3952 18052 4004
rect 18104 3992 18110 4004
rect 18104 3964 18906 3992
rect 18104 3952 18110 3964
rect 8938 3924 8944 3936
rect 8899 3896 8944 3924
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 9766 3924 9772 3936
rect 9727 3896 9772 3924
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 10229 3927 10287 3933
rect 10229 3893 10241 3927
rect 10275 3924 10287 3927
rect 11054 3924 11060 3936
rect 10275 3896 11060 3924
rect 10275 3893 10287 3896
rect 10229 3887 10287 3893
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 12069 3927 12127 3933
rect 12069 3924 12081 3927
rect 11204 3896 12081 3924
rect 11204 3884 11210 3896
rect 12069 3893 12081 3896
rect 12115 3893 12127 3927
rect 12069 3887 12127 3893
rect 14642 3884 14648 3936
rect 14700 3924 14706 3936
rect 14737 3927 14795 3933
rect 14737 3924 14749 3927
rect 14700 3896 14749 3924
rect 14700 3884 14706 3896
rect 14737 3893 14749 3896
rect 14783 3893 14795 3927
rect 14737 3887 14795 3893
rect 14829 3927 14887 3933
rect 14829 3893 14841 3927
rect 14875 3924 14887 3927
rect 15378 3924 15384 3936
rect 14875 3896 15384 3924
rect 14875 3893 14887 3896
rect 14829 3887 14887 3893
rect 15378 3884 15384 3896
rect 15436 3884 15442 3936
rect 20162 3924 20168 3936
rect 20123 3896 20168 3924
rect 20162 3884 20168 3896
rect 20220 3884 20226 3936
rect 1104 3834 21804 3856
rect 1104 3782 7882 3834
rect 7934 3782 7946 3834
rect 7998 3782 8010 3834
rect 8062 3782 8074 3834
rect 8126 3782 14782 3834
rect 14834 3782 14846 3834
rect 14898 3782 14910 3834
rect 14962 3782 14974 3834
rect 15026 3782 21804 3834
rect 1104 3760 21804 3782
rect 8573 3723 8631 3729
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 8938 3720 8944 3732
rect 8619 3692 8944 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 8938 3680 8944 3692
rect 8996 3720 9002 3732
rect 10042 3720 10048 3732
rect 8996 3692 10048 3720
rect 8996 3680 9002 3692
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 10410 3680 10416 3732
rect 10468 3720 10474 3732
rect 11241 3723 11299 3729
rect 11241 3720 11253 3723
rect 10468 3692 11253 3720
rect 10468 3680 10474 3692
rect 11241 3689 11253 3692
rect 11287 3689 11299 3723
rect 11241 3683 11299 3689
rect 11333 3723 11391 3729
rect 11333 3689 11345 3723
rect 11379 3720 11391 3723
rect 12713 3723 12771 3729
rect 12713 3720 12725 3723
rect 11379 3692 12725 3720
rect 11379 3689 11391 3692
rect 11333 3683 11391 3689
rect 12713 3689 12725 3692
rect 12759 3689 12771 3723
rect 15562 3720 15568 3732
rect 12713 3683 12771 3689
rect 15028 3692 15568 3720
rect 3786 3612 3792 3664
rect 3844 3652 3850 3664
rect 4341 3655 4399 3661
rect 4341 3652 4353 3655
rect 3844 3624 4353 3652
rect 3844 3612 3850 3624
rect 4341 3621 4353 3624
rect 4387 3621 4399 3655
rect 4341 3615 4399 3621
rect 10502 3612 10508 3664
rect 10560 3652 10566 3664
rect 13170 3652 13176 3664
rect 10560 3624 13176 3652
rect 10560 3612 10566 3624
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 6914 3584 6920 3596
rect 6875 3556 6920 3584
rect 6914 3544 6920 3556
rect 6972 3544 6978 3596
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3516 8263 3519
rect 9030 3516 9036 3528
rect 8251 3488 9036 3516
rect 8251 3485 8263 3488
rect 8205 3479 8263 3485
rect 9030 3476 9036 3488
rect 9088 3476 9094 3528
rect 11440 3525 11468 3624
rect 13170 3612 13176 3624
rect 13228 3612 13234 3664
rect 15028 3661 15056 3692
rect 15562 3680 15568 3692
rect 15620 3720 15626 3732
rect 15933 3723 15991 3729
rect 15933 3720 15945 3723
rect 15620 3692 15945 3720
rect 15620 3680 15626 3692
rect 15933 3689 15945 3692
rect 15979 3689 15991 3723
rect 15933 3683 15991 3689
rect 15013 3655 15071 3661
rect 15013 3621 15025 3655
rect 15059 3621 15071 3655
rect 15013 3615 15071 3621
rect 15378 3612 15384 3664
rect 15436 3652 15442 3664
rect 15436 3624 15976 3652
rect 15436 3612 15442 3624
rect 12253 3587 12311 3593
rect 12253 3553 12265 3587
rect 12299 3584 12311 3587
rect 12618 3584 12624 3596
rect 12299 3556 12624 3584
rect 12299 3553 12311 3556
rect 12253 3547 12311 3553
rect 12618 3544 12624 3556
rect 12676 3544 12682 3596
rect 12897 3587 12955 3593
rect 12897 3553 12909 3587
rect 12943 3553 12955 3587
rect 12897 3547 12955 3553
rect 11425 3519 11483 3525
rect 11425 3485 11437 3519
rect 11471 3485 11483 3519
rect 11425 3479 11483 3485
rect 11974 3476 11980 3528
rect 12032 3516 12038 3528
rect 12912 3516 12940 3547
rect 13906 3544 13912 3596
rect 13964 3584 13970 3596
rect 15948 3593 15976 3624
rect 14921 3587 14979 3593
rect 14921 3584 14933 3587
rect 13964 3556 14933 3584
rect 13964 3544 13970 3556
rect 14921 3553 14933 3556
rect 14967 3553 14979 3587
rect 14921 3547 14979 3553
rect 15473 3587 15531 3593
rect 15473 3553 15485 3587
rect 15519 3553 15531 3587
rect 15473 3547 15531 3553
rect 15933 3587 15991 3593
rect 15933 3553 15945 3587
rect 15979 3553 15991 3587
rect 21082 3584 21088 3596
rect 21043 3556 21088 3584
rect 15933 3547 15991 3553
rect 15488 3516 15516 3547
rect 21082 3544 21088 3556
rect 21140 3544 21146 3596
rect 15562 3516 15568 3528
rect 12032 3488 12940 3516
rect 15475 3488 15568 3516
rect 12032 3476 12038 3488
rect 15562 3476 15568 3488
rect 15620 3516 15626 3528
rect 16301 3519 16359 3525
rect 16301 3516 16313 3519
rect 15620 3488 16313 3516
rect 15620 3476 15626 3488
rect 16301 3485 16313 3488
rect 16347 3485 16359 3519
rect 16301 3479 16359 3485
rect 8573 3451 8631 3457
rect 8573 3417 8585 3451
rect 8619 3448 8631 3451
rect 9493 3451 9551 3457
rect 9493 3448 9505 3451
rect 8619 3420 9505 3448
rect 8619 3417 8631 3420
rect 8573 3411 8631 3417
rect 9493 3417 9505 3420
rect 9539 3417 9551 3451
rect 20806 3448 20812 3460
rect 9493 3411 9551 3417
rect 10336 3420 20812 3448
rect 1578 3380 1584 3392
rect 1539 3352 1584 3380
rect 1578 3340 1584 3352
rect 1636 3340 1642 3392
rect 4433 3383 4491 3389
rect 4433 3349 4445 3383
rect 4479 3380 4491 3383
rect 6638 3380 6644 3392
rect 4479 3352 6644 3380
rect 4479 3349 4491 3352
rect 4433 3343 4491 3349
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 6730 3340 6736 3392
rect 6788 3380 6794 3392
rect 6788 3352 6833 3380
rect 6788 3340 6794 3352
rect 8202 3340 8208 3392
rect 8260 3380 8266 3392
rect 10336 3380 10364 3420
rect 20806 3408 20812 3420
rect 20864 3408 20870 3460
rect 10870 3380 10876 3392
rect 8260 3352 10364 3380
rect 10831 3352 10876 3380
rect 8260 3340 8266 3352
rect 10870 3340 10876 3352
rect 10928 3340 10934 3392
rect 12066 3380 12072 3392
rect 12027 3352 12072 3380
rect 12066 3340 12072 3352
rect 12124 3340 12130 3392
rect 16022 3340 16028 3392
rect 16080 3380 16086 3392
rect 20901 3383 20959 3389
rect 20901 3380 20913 3383
rect 16080 3352 20913 3380
rect 16080 3340 16086 3352
rect 20901 3349 20913 3352
rect 20947 3349 20959 3383
rect 20901 3343 20959 3349
rect 1104 3290 21804 3312
rect 1104 3238 4432 3290
rect 4484 3238 4496 3290
rect 4548 3238 4560 3290
rect 4612 3238 4624 3290
rect 4676 3238 11332 3290
rect 11384 3238 11396 3290
rect 11448 3238 11460 3290
rect 11512 3238 11524 3290
rect 11576 3238 18232 3290
rect 18284 3238 18296 3290
rect 18348 3238 18360 3290
rect 18412 3238 18424 3290
rect 18476 3238 21804 3290
rect 1104 3216 21804 3238
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 9030 3176 9036 3188
rect 6696 3148 8708 3176
rect 8991 3148 9036 3176
rect 6696 3136 6702 3148
rect 1578 3068 1584 3120
rect 1636 3108 1642 3120
rect 8680 3108 8708 3148
rect 9030 3136 9036 3148
rect 9088 3136 9094 3188
rect 10042 3176 10048 3188
rect 10003 3148 10048 3176
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 11146 3176 11152 3188
rect 11107 3148 11152 3176
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 12161 3179 12219 3185
rect 12161 3145 12173 3179
rect 12207 3176 12219 3179
rect 12526 3176 12532 3188
rect 12207 3148 12532 3176
rect 12207 3145 12219 3148
rect 12161 3139 12219 3145
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 14642 3176 14648 3188
rect 14603 3148 14648 3176
rect 14642 3136 14648 3148
rect 14700 3136 14706 3188
rect 15562 3176 15568 3188
rect 15523 3148 15568 3176
rect 15562 3136 15568 3148
rect 15620 3136 15626 3188
rect 20806 3136 20812 3188
rect 20864 3176 20870 3188
rect 20901 3179 20959 3185
rect 20901 3176 20913 3179
rect 20864 3148 20913 3176
rect 20864 3136 20870 3148
rect 20901 3145 20913 3148
rect 20947 3145 20959 3179
rect 20901 3139 20959 3145
rect 13906 3108 13912 3120
rect 1636 3080 2774 3108
rect 8680 3080 13912 3108
rect 1636 3068 1642 3080
rect 474 2932 480 2984
rect 532 2972 538 2984
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 532 2944 1409 2972
rect 532 2932 538 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 2746 2972 2774 3080
rect 13906 3068 13912 3080
rect 13964 3068 13970 3120
rect 14016 3080 16160 3108
rect 8478 3040 8484 3052
rect 8439 3012 8484 3040
rect 8478 3000 8484 3012
rect 8536 3000 8542 3052
rect 12618 3040 12624 3052
rect 11164 3012 12624 3040
rect 8573 2975 8631 2981
rect 8573 2972 8585 2975
rect 2746 2944 8585 2972
rect 1397 2935 1455 2941
rect 8573 2941 8585 2944
rect 8619 2941 8631 2975
rect 8573 2935 8631 2941
rect 8665 2975 8723 2981
rect 8665 2941 8677 2975
rect 8711 2972 8723 2975
rect 8754 2972 8760 2984
rect 8711 2944 8760 2972
rect 8711 2941 8723 2944
rect 8665 2935 8723 2941
rect 8754 2932 8760 2944
rect 8812 2932 8818 2984
rect 9030 2932 9036 2984
rect 9088 2972 9094 2984
rect 9493 2975 9551 2981
rect 9493 2972 9505 2975
rect 9088 2944 9505 2972
rect 9088 2932 9094 2944
rect 9493 2941 9505 2944
rect 9539 2941 9551 2975
rect 9493 2935 9551 2941
rect 9674 2932 9680 2984
rect 9732 2972 9738 2984
rect 10045 2975 10103 2981
rect 10045 2972 10057 2975
rect 9732 2944 10057 2972
rect 9732 2932 9738 2944
rect 10045 2941 10057 2944
rect 10091 2941 10103 2975
rect 10045 2935 10103 2941
rect 10597 2975 10655 2981
rect 10597 2941 10609 2975
rect 10643 2972 10655 2975
rect 10870 2972 10876 2984
rect 10643 2944 10876 2972
rect 10643 2941 10655 2944
rect 10597 2935 10655 2941
rect 10870 2932 10876 2944
rect 10928 2932 10934 2984
rect 11164 2981 11192 3012
rect 12618 3000 12624 3012
rect 12676 3000 12682 3052
rect 13170 3040 13176 3052
rect 13131 3012 13176 3040
rect 13170 3000 13176 3012
rect 13228 3040 13234 3052
rect 14016 3040 14044 3080
rect 16132 3052 16160 3080
rect 16022 3040 16028 3052
rect 13228 3012 14044 3040
rect 14108 3012 15884 3040
rect 15983 3012 16028 3040
rect 13228 3000 13234 3012
rect 11149 2975 11207 2981
rect 11149 2941 11161 2975
rect 11195 2941 11207 2975
rect 11149 2935 11207 2941
rect 11698 2932 11704 2984
rect 11756 2972 11762 2984
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 11756 2944 12081 2972
rect 11756 2932 11762 2944
rect 12069 2941 12081 2944
rect 12115 2941 12127 2975
rect 14108 2972 14136 3012
rect 14274 2972 14280 2984
rect 12069 2935 12127 2941
rect 12406 2944 14136 2972
rect 14235 2944 14280 2972
rect 6730 2864 6736 2916
rect 6788 2904 6794 2916
rect 12406 2904 12434 2944
rect 14274 2932 14280 2944
rect 14332 2932 14338 2984
rect 14642 2972 14648 2984
rect 14603 2944 14648 2972
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 15856 2972 15884 3012
rect 16022 3000 16028 3012
rect 16080 3000 16086 3052
rect 16114 3000 16120 3052
rect 16172 3040 16178 3052
rect 17310 3040 17316 3052
rect 16172 3012 16265 3040
rect 17271 3012 17316 3040
rect 16172 3000 16178 3012
rect 17310 3000 17316 3012
rect 17368 3000 17374 3052
rect 17589 3043 17647 3049
rect 17589 3009 17601 3043
rect 17635 3040 17647 3043
rect 17635 3012 19380 3040
rect 17635 3009 17647 3012
rect 17589 3003 17647 3009
rect 19352 2981 19380 3012
rect 19337 2975 19395 2981
rect 15856 2944 16436 2972
rect 15933 2907 15991 2913
rect 15933 2904 15945 2907
rect 6788 2876 12434 2904
rect 12820 2876 15945 2904
rect 6788 2864 6794 2876
rect 1581 2839 1639 2845
rect 1581 2805 1593 2839
rect 1627 2836 1639 2839
rect 1670 2836 1676 2848
rect 1627 2808 1676 2836
rect 1627 2805 1639 2808
rect 1581 2799 1639 2805
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 7282 2796 7288 2848
rect 7340 2836 7346 2848
rect 12820 2836 12848 2876
rect 15933 2873 15945 2876
rect 15979 2873 15991 2907
rect 15933 2867 15991 2873
rect 7340 2808 12848 2836
rect 7340 2796 7346 2808
rect 12894 2796 12900 2848
rect 12952 2836 12958 2848
rect 13357 2839 13415 2845
rect 13357 2836 13369 2839
rect 12952 2808 13369 2836
rect 12952 2796 12958 2808
rect 13357 2805 13369 2808
rect 13403 2805 13415 2839
rect 13357 2799 13415 2805
rect 13446 2796 13452 2848
rect 13504 2836 13510 2848
rect 13814 2836 13820 2848
rect 13504 2808 13549 2836
rect 13775 2808 13820 2836
rect 13504 2796 13510 2808
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 16408 2836 16436 2944
rect 19337 2941 19349 2975
rect 19383 2972 19395 2975
rect 19610 2972 19616 2984
rect 19383 2944 19616 2972
rect 19383 2941 19395 2944
rect 19337 2935 19395 2941
rect 19610 2932 19616 2944
rect 19668 2932 19674 2984
rect 21085 2975 21143 2981
rect 21085 2941 21097 2975
rect 21131 2972 21143 2975
rect 22094 2972 22100 2984
rect 21131 2944 22100 2972
rect 21131 2941 21143 2944
rect 21085 2935 21143 2941
rect 22094 2932 22100 2944
rect 22152 2932 22158 2984
rect 18046 2864 18052 2916
rect 18104 2864 18110 2916
rect 18064 2836 18092 2864
rect 16408 2808 18092 2836
rect 1104 2746 21804 2768
rect 1104 2694 7882 2746
rect 7934 2694 7946 2746
rect 7998 2694 8010 2746
rect 8062 2694 8074 2746
rect 8126 2694 14782 2746
rect 14834 2694 14846 2746
rect 14898 2694 14910 2746
rect 14962 2694 14974 2746
rect 15026 2694 21804 2746
rect 1104 2672 21804 2694
rect 4433 2635 4491 2641
rect 4433 2601 4445 2635
rect 4479 2632 4491 2635
rect 4798 2632 4804 2644
rect 4479 2604 4804 2632
rect 4479 2601 4491 2604
rect 4433 2595 4491 2601
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 5721 2635 5779 2641
rect 5721 2601 5733 2635
rect 5767 2632 5779 2635
rect 5810 2632 5816 2644
rect 5767 2604 5816 2632
rect 5767 2601 5779 2604
rect 5721 2595 5779 2601
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 6914 2592 6920 2644
rect 6972 2632 6978 2644
rect 7009 2635 7067 2641
rect 7009 2632 7021 2635
rect 6972 2604 7021 2632
rect 6972 2592 6978 2604
rect 7009 2601 7021 2604
rect 7055 2601 7067 2635
rect 9766 2632 9772 2644
rect 9727 2604 9772 2632
rect 7009 2595 7067 2601
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 11146 2592 11152 2644
rect 11204 2632 11210 2644
rect 11333 2635 11391 2641
rect 11333 2632 11345 2635
rect 11204 2604 11345 2632
rect 11204 2592 11210 2604
rect 11333 2601 11345 2604
rect 11379 2601 11391 2635
rect 12894 2632 12900 2644
rect 12855 2604 12900 2632
rect 11333 2595 11391 2601
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 14642 2592 14648 2644
rect 14700 2632 14706 2644
rect 14921 2635 14979 2641
rect 14921 2632 14933 2635
rect 14700 2604 14933 2632
rect 14700 2592 14706 2604
rect 14921 2601 14933 2604
rect 14967 2601 14979 2635
rect 14921 2595 14979 2601
rect 18782 2592 18788 2644
rect 18840 2632 18846 2644
rect 18877 2635 18935 2641
rect 18877 2632 18889 2635
rect 18840 2604 18889 2632
rect 18840 2592 18846 2604
rect 18877 2601 18889 2604
rect 18923 2601 18935 2635
rect 18877 2595 18935 2601
rect 2038 2564 2044 2576
rect 1999 2536 2044 2564
rect 2038 2524 2044 2536
rect 2096 2524 2102 2576
rect 13814 2564 13820 2576
rect 13372 2536 13820 2564
rect 3694 2456 3700 2508
rect 3752 2496 3758 2508
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 3752 2468 4261 2496
rect 3752 2456 3758 2468
rect 4249 2465 4261 2468
rect 4295 2465 4307 2499
rect 5534 2496 5540 2508
rect 5495 2468 5540 2496
rect 4249 2459 4307 2465
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 7101 2499 7159 2505
rect 7101 2496 7113 2499
rect 6972 2468 7113 2496
rect 6972 2456 6978 2468
rect 7101 2465 7113 2468
rect 7147 2465 7159 2499
rect 7101 2459 7159 2465
rect 8754 2456 8760 2508
rect 8812 2496 8818 2508
rect 9585 2499 9643 2505
rect 9585 2496 9597 2499
rect 8812 2468 9597 2496
rect 8812 2456 8818 2468
rect 9585 2465 9597 2468
rect 9631 2465 9643 2499
rect 9585 2459 9643 2465
rect 10321 2499 10379 2505
rect 10321 2465 10333 2499
rect 10367 2496 10379 2499
rect 10594 2496 10600 2508
rect 10367 2468 10600 2496
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 10594 2456 10600 2468
rect 10652 2456 10658 2508
rect 10870 2456 10876 2508
rect 10928 2496 10934 2508
rect 10965 2499 11023 2505
rect 10965 2496 10977 2499
rect 10928 2468 10977 2496
rect 10928 2456 10934 2468
rect 10965 2465 10977 2468
rect 11011 2465 11023 2499
rect 10965 2459 11023 2465
rect 11333 2499 11391 2505
rect 11333 2465 11345 2499
rect 11379 2496 11391 2499
rect 12066 2496 12072 2508
rect 11379 2468 12072 2496
rect 11379 2465 11391 2468
rect 11333 2459 11391 2465
rect 12066 2456 12072 2468
rect 12124 2456 12130 2508
rect 13372 2505 13400 2536
rect 13814 2524 13820 2536
rect 13872 2564 13878 2576
rect 14274 2564 14280 2576
rect 13872 2536 14280 2564
rect 13872 2524 13878 2536
rect 14274 2524 14280 2536
rect 14332 2524 14338 2576
rect 17862 2564 17868 2576
rect 17823 2536 17868 2564
rect 17862 2524 17868 2536
rect 17920 2524 17926 2576
rect 20162 2524 20168 2576
rect 20220 2564 20226 2576
rect 20901 2567 20959 2573
rect 20901 2564 20913 2567
rect 20220 2536 20913 2564
rect 20220 2524 20226 2536
rect 20901 2533 20913 2536
rect 20947 2533 20959 2567
rect 20901 2527 20959 2533
rect 12713 2499 12771 2505
rect 12713 2465 12725 2499
rect 12759 2465 12771 2499
rect 12713 2459 12771 2465
rect 13357 2499 13415 2505
rect 13357 2465 13369 2499
rect 13403 2465 13415 2499
rect 13906 2496 13912 2508
rect 13867 2468 13912 2496
rect 13357 2459 13415 2465
rect 12728 2428 12756 2459
rect 13906 2456 13912 2468
rect 13964 2496 13970 2508
rect 15105 2499 15163 2505
rect 15105 2496 15117 2499
rect 13964 2468 15117 2496
rect 13964 2456 13970 2468
rect 15105 2465 15117 2468
rect 15151 2465 15163 2499
rect 15654 2496 15660 2508
rect 15615 2468 15660 2496
rect 15105 2459 15163 2465
rect 15654 2456 15660 2468
rect 15712 2456 15718 2508
rect 17034 2456 17040 2508
rect 17092 2496 17098 2508
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 17092 2468 17693 2496
rect 17092 2456 17098 2468
rect 17681 2465 17693 2468
rect 17727 2465 17739 2499
rect 17681 2459 17739 2465
rect 18874 2456 18880 2508
rect 18932 2496 18938 2508
rect 19061 2499 19119 2505
rect 19061 2496 19073 2499
rect 18932 2468 19073 2496
rect 18932 2456 18938 2468
rect 19061 2465 19073 2468
rect 19107 2465 19119 2499
rect 19061 2459 19119 2465
rect 13814 2428 13820 2440
rect 12728 2400 13820 2428
rect 13814 2388 13820 2400
rect 13872 2388 13878 2440
rect 16114 2428 16120 2440
rect 16075 2400 16120 2428
rect 16114 2388 16120 2400
rect 16172 2388 16178 2440
rect 1854 2360 1860 2372
rect 1815 2332 1860 2360
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 10505 2363 10563 2369
rect 10505 2329 10517 2363
rect 10551 2360 10563 2363
rect 20714 2360 20720 2372
rect 10551 2332 16574 2360
rect 20675 2332 20720 2360
rect 10551 2329 10563 2332
rect 10505 2323 10563 2329
rect 13909 2295 13967 2301
rect 13909 2261 13921 2295
rect 13955 2292 13967 2295
rect 14550 2292 14556 2304
rect 13955 2264 14556 2292
rect 13955 2261 13967 2264
rect 13909 2255 13967 2261
rect 14550 2252 14556 2264
rect 14608 2252 14614 2304
rect 16546 2292 16574 2332
rect 20714 2320 20720 2332
rect 20772 2320 20778 2372
rect 17494 2292 17500 2304
rect 16546 2264 17500 2292
rect 17494 2252 17500 2264
rect 17552 2252 17558 2304
rect 1104 2202 21804 2224
rect 1104 2150 4432 2202
rect 4484 2150 4496 2202
rect 4548 2150 4560 2202
rect 4612 2150 4624 2202
rect 4676 2150 11332 2202
rect 11384 2150 11396 2202
rect 11448 2150 11460 2202
rect 11512 2150 11524 2202
rect 11576 2150 18232 2202
rect 18284 2150 18296 2202
rect 18348 2150 18360 2202
rect 18412 2150 18424 2202
rect 18476 2150 21804 2202
rect 1104 2128 21804 2150
<< via1 >>
rect 4432 22822 4484 22874
rect 4496 22822 4548 22874
rect 4560 22822 4612 22874
rect 4624 22822 4676 22874
rect 11332 22822 11384 22874
rect 11396 22822 11448 22874
rect 11460 22822 11512 22874
rect 11524 22822 11576 22874
rect 18232 22822 18284 22874
rect 18296 22822 18348 22874
rect 18360 22822 18412 22874
rect 18424 22822 18476 22874
rect 1492 22763 1544 22772
rect 1492 22729 1501 22763
rect 1501 22729 1535 22763
rect 1535 22729 1544 22763
rect 1492 22720 1544 22729
rect 5448 22652 5500 22704
rect 11060 22652 11112 22704
rect 940 22516 992 22568
rect 2780 22559 2832 22568
rect 2780 22525 2789 22559
rect 2789 22525 2823 22559
rect 2823 22525 2832 22559
rect 4712 22559 4764 22568
rect 2780 22516 2832 22525
rect 4712 22525 4721 22559
rect 4721 22525 4755 22559
rect 4755 22525 4764 22559
rect 4712 22516 4764 22525
rect 4804 22516 4856 22568
rect 6000 22516 6052 22568
rect 7840 22559 7892 22568
rect 7840 22525 7849 22559
rect 7849 22525 7883 22559
rect 7883 22525 7892 22559
rect 7840 22516 7892 22525
rect 9680 22559 9732 22568
rect 9680 22525 9689 22559
rect 9689 22525 9723 22559
rect 9723 22525 9732 22559
rect 9680 22516 9732 22525
rect 11704 22516 11756 22568
rect 12900 22559 12952 22568
rect 12900 22525 12909 22559
rect 12909 22525 12943 22559
rect 12943 22525 12952 22559
rect 12900 22516 12952 22525
rect 14740 22516 14792 22568
rect 16580 22516 16632 22568
rect 17960 22516 18012 22568
rect 19800 22516 19852 22568
rect 21640 22516 21692 22568
rect 1584 22491 1636 22500
rect 1584 22457 1593 22491
rect 1593 22457 1627 22491
rect 1627 22457 1636 22491
rect 1584 22448 1636 22457
rect 2044 22380 2096 22432
rect 4896 22423 4948 22432
rect 4896 22389 4905 22423
rect 4905 22389 4939 22423
rect 4939 22389 4948 22423
rect 4896 22380 4948 22389
rect 6184 22380 6236 22432
rect 7012 22380 7064 22432
rect 10600 22380 10652 22432
rect 12348 22380 12400 22432
rect 12716 22380 12768 22432
rect 14648 22380 14700 22432
rect 16304 22380 16356 22432
rect 17960 22423 18012 22432
rect 17960 22389 17969 22423
rect 17969 22389 18003 22423
rect 18003 22389 18012 22423
rect 17960 22380 18012 22389
rect 19156 22423 19208 22432
rect 19156 22389 19165 22423
rect 19165 22389 19199 22423
rect 19199 22389 19208 22423
rect 19156 22380 19208 22389
rect 21180 22380 21232 22432
rect 7882 22278 7934 22330
rect 7946 22278 7998 22330
rect 8010 22278 8062 22330
rect 8074 22278 8126 22330
rect 14782 22278 14834 22330
rect 14846 22278 14898 22330
rect 14910 22278 14962 22330
rect 14974 22278 15026 22330
rect 10876 22151 10928 22160
rect 10876 22117 10885 22151
rect 10885 22117 10919 22151
rect 10919 22117 10928 22151
rect 11888 22151 11940 22160
rect 10876 22108 10928 22117
rect 11888 22117 11897 22151
rect 11897 22117 11931 22151
rect 11931 22117 11940 22151
rect 11888 22108 11940 22117
rect 4988 22083 5040 22092
rect 4988 22049 4997 22083
rect 4997 22049 5031 22083
rect 5031 22049 5040 22083
rect 4988 22040 5040 22049
rect 5080 22083 5132 22092
rect 5080 22049 5089 22083
rect 5089 22049 5123 22083
rect 5123 22049 5132 22083
rect 5080 22040 5132 22049
rect 5540 22040 5592 22092
rect 4712 21972 4764 22024
rect 10324 22040 10376 22092
rect 11704 22083 11756 22092
rect 11704 22049 11713 22083
rect 11713 22049 11747 22083
rect 11747 22049 11756 22083
rect 11704 22040 11756 22049
rect 11980 22083 12032 22092
rect 11980 22049 11989 22083
rect 11989 22049 12023 22083
rect 12023 22049 12032 22083
rect 11980 22040 12032 22049
rect 12164 22040 12216 22092
rect 12900 22083 12952 22092
rect 12900 22049 12909 22083
rect 12909 22049 12943 22083
rect 12943 22049 12952 22083
rect 12900 22040 12952 22049
rect 17500 22040 17552 22092
rect 20536 22040 20588 22092
rect 21088 22083 21140 22092
rect 21088 22049 21097 22083
rect 21097 22049 21131 22083
rect 21131 22049 21140 22083
rect 21088 22040 21140 22049
rect 15292 21904 15344 21956
rect 4160 21836 4212 21888
rect 5264 21879 5316 21888
rect 5264 21845 5273 21879
rect 5273 21845 5307 21879
rect 5307 21845 5316 21879
rect 5264 21836 5316 21845
rect 7748 21879 7800 21888
rect 7748 21845 7757 21879
rect 7757 21845 7791 21879
rect 7791 21845 7800 21879
rect 7748 21836 7800 21845
rect 10048 21879 10100 21888
rect 10048 21845 10057 21879
rect 10057 21845 10091 21879
rect 10091 21845 10100 21879
rect 10048 21836 10100 21845
rect 10692 21879 10744 21888
rect 10692 21845 10701 21879
rect 10701 21845 10735 21879
rect 10735 21845 10744 21879
rect 10692 21836 10744 21845
rect 12256 21879 12308 21888
rect 12256 21845 12265 21879
rect 12265 21845 12299 21879
rect 12299 21845 12308 21879
rect 12256 21836 12308 21845
rect 12808 21836 12860 21888
rect 15200 21879 15252 21888
rect 15200 21845 15209 21879
rect 15209 21845 15243 21879
rect 15243 21845 15252 21879
rect 15200 21836 15252 21845
rect 18696 21836 18748 21888
rect 20076 21836 20128 21888
rect 4432 21734 4484 21786
rect 4496 21734 4548 21786
rect 4560 21734 4612 21786
rect 4624 21734 4676 21786
rect 11332 21734 11384 21786
rect 11396 21734 11448 21786
rect 11460 21734 11512 21786
rect 11524 21734 11576 21786
rect 18232 21734 18284 21786
rect 18296 21734 18348 21786
rect 18360 21734 18412 21786
rect 18424 21734 18476 21786
rect 1584 21632 1636 21684
rect 10876 21675 10928 21684
rect 10876 21641 10885 21675
rect 10885 21641 10919 21675
rect 10919 21641 10928 21675
rect 10876 21632 10928 21641
rect 8208 21564 8260 21616
rect 20168 21564 20220 21616
rect 4160 21539 4212 21548
rect 4160 21505 4169 21539
rect 4169 21505 4203 21539
rect 4203 21505 4212 21539
rect 4160 21496 4212 21505
rect 9128 21539 9180 21548
rect 2504 21428 2556 21480
rect 9128 21505 9137 21539
rect 9137 21505 9171 21539
rect 9171 21505 9180 21539
rect 9128 21496 9180 21505
rect 10692 21496 10744 21548
rect 12256 21496 12308 21548
rect 16212 21496 16264 21548
rect 19064 21496 19116 21548
rect 4896 21360 4948 21412
rect 20168 21471 20220 21480
rect 7196 21360 7248 21412
rect 7748 21360 7800 21412
rect 10048 21360 10100 21412
rect 5540 21292 5592 21344
rect 9128 21292 9180 21344
rect 12072 21335 12124 21344
rect 12072 21301 12081 21335
rect 12081 21301 12115 21335
rect 12115 21301 12124 21335
rect 12072 21292 12124 21301
rect 12808 21360 12860 21412
rect 20168 21437 20177 21471
rect 20177 21437 20211 21471
rect 20211 21437 20220 21471
rect 20168 21428 20220 21437
rect 15200 21360 15252 21412
rect 15752 21403 15804 21412
rect 15752 21369 15761 21403
rect 15761 21369 15795 21403
rect 15795 21369 15804 21403
rect 15752 21360 15804 21369
rect 17960 21360 18012 21412
rect 18696 21360 18748 21412
rect 14280 21335 14332 21344
rect 14280 21301 14289 21335
rect 14289 21301 14323 21335
rect 14323 21301 14332 21335
rect 14280 21292 14332 21301
rect 15476 21292 15528 21344
rect 21088 21428 21140 21480
rect 19340 21292 19392 21344
rect 7882 21190 7934 21242
rect 7946 21190 7998 21242
rect 8010 21190 8062 21242
rect 8074 21190 8126 21242
rect 14782 21190 14834 21242
rect 14846 21190 14898 21242
rect 14910 21190 14962 21242
rect 14974 21190 15026 21242
rect 4988 21088 5040 21140
rect 7196 21131 7248 21140
rect 7196 21097 7205 21131
rect 7205 21097 7239 21131
rect 7239 21097 7248 21131
rect 7196 21088 7248 21097
rect 11704 21088 11756 21140
rect 11980 21088 12032 21140
rect 12164 21088 12216 21140
rect 7472 21063 7524 21072
rect 7472 21029 7481 21063
rect 7481 21029 7515 21063
rect 7515 21029 7524 21063
rect 7472 21020 7524 21029
rect 7656 21020 7708 21072
rect 8208 21020 8260 21072
rect 12072 21063 12124 21072
rect 12072 21029 12081 21063
rect 12081 21029 12115 21063
rect 12115 21029 12124 21063
rect 12072 21020 12124 21029
rect 5540 20952 5592 21004
rect 7380 20995 7432 21004
rect 7380 20961 7389 20995
rect 7389 20961 7423 20995
rect 7423 20961 7432 20995
rect 7380 20952 7432 20961
rect 8484 20952 8536 21004
rect 11980 20995 12032 21004
rect 11980 20961 11989 20995
rect 11989 20961 12023 20995
rect 12023 20961 12032 20995
rect 11980 20952 12032 20961
rect 12164 20995 12216 21004
rect 12164 20961 12173 20995
rect 12173 20961 12207 20995
rect 12207 20961 12216 20995
rect 14280 21020 14332 21072
rect 15752 21088 15804 21140
rect 17224 21020 17276 21072
rect 12164 20952 12216 20961
rect 5080 20816 5132 20868
rect 15476 20952 15528 21004
rect 16212 20995 16264 21004
rect 16212 20961 16221 20995
rect 16221 20961 16255 20995
rect 16255 20961 16264 20995
rect 16212 20952 16264 20961
rect 20812 20952 20864 21004
rect 15660 20884 15712 20936
rect 16488 20927 16540 20936
rect 16488 20893 16497 20927
rect 16497 20893 16531 20927
rect 16531 20893 16540 20927
rect 16488 20884 16540 20893
rect 15384 20816 15436 20868
rect 4988 20748 5040 20800
rect 5264 20748 5316 20800
rect 11796 20791 11848 20800
rect 11796 20757 11805 20791
rect 11805 20757 11839 20791
rect 11839 20757 11848 20791
rect 11796 20748 11848 20757
rect 15660 20748 15712 20800
rect 20628 20748 20680 20800
rect 4432 20646 4484 20698
rect 4496 20646 4548 20698
rect 4560 20646 4612 20698
rect 4624 20646 4676 20698
rect 11332 20646 11384 20698
rect 11396 20646 11448 20698
rect 11460 20646 11512 20698
rect 11524 20646 11576 20698
rect 18232 20646 18284 20698
rect 18296 20646 18348 20698
rect 18360 20646 18412 20698
rect 18424 20646 18476 20698
rect 7380 20544 7432 20596
rect 12072 20544 12124 20596
rect 12164 20476 12216 20528
rect 12532 20519 12584 20528
rect 2504 20451 2556 20460
rect 2504 20417 2513 20451
rect 2513 20417 2547 20451
rect 2547 20417 2556 20451
rect 2504 20408 2556 20417
rect 9128 20408 9180 20460
rect 11796 20408 11848 20460
rect 1400 20383 1452 20392
rect 1400 20349 1409 20383
rect 1409 20349 1443 20383
rect 1443 20349 1452 20383
rect 1400 20340 1452 20349
rect 5264 20383 5316 20392
rect 5264 20349 5273 20383
rect 5273 20349 5307 20383
rect 5307 20349 5316 20383
rect 5264 20340 5316 20349
rect 5540 20340 5592 20392
rect 6000 20340 6052 20392
rect 7656 20383 7708 20392
rect 7656 20349 7665 20383
rect 7665 20349 7699 20383
rect 7699 20349 7708 20383
rect 7656 20340 7708 20349
rect 7748 20340 7800 20392
rect 11888 20340 11940 20392
rect 12532 20485 12541 20519
rect 12541 20485 12575 20519
rect 12575 20485 12584 20519
rect 12532 20476 12584 20485
rect 17224 20544 17276 20596
rect 14280 20476 14332 20528
rect 14556 20408 14608 20460
rect 14280 20383 14332 20392
rect 1492 20204 1544 20256
rect 3332 20272 3384 20324
rect 10416 20272 10468 20324
rect 11980 20272 12032 20324
rect 14280 20349 14289 20383
rect 14289 20349 14323 20383
rect 14323 20349 14332 20383
rect 14280 20340 14332 20349
rect 14924 20408 14976 20460
rect 16212 20408 16264 20460
rect 19340 20451 19392 20460
rect 19340 20417 19349 20451
rect 19349 20417 19383 20451
rect 19383 20417 19392 20451
rect 19340 20408 19392 20417
rect 15660 20340 15712 20392
rect 17500 20383 17552 20392
rect 17500 20349 17509 20383
rect 17509 20349 17543 20383
rect 17543 20349 17552 20383
rect 17500 20340 17552 20349
rect 19064 20383 19116 20392
rect 19064 20349 19073 20383
rect 19073 20349 19107 20383
rect 19107 20349 19116 20383
rect 19064 20340 19116 20349
rect 14464 20272 14516 20324
rect 14924 20315 14976 20324
rect 14924 20281 14933 20315
rect 14933 20281 14967 20315
rect 14967 20281 14976 20315
rect 14924 20272 14976 20281
rect 20076 20272 20128 20324
rect 4160 20204 4212 20256
rect 5172 20204 5224 20256
rect 5356 20247 5408 20256
rect 5356 20213 5365 20247
rect 5365 20213 5399 20247
rect 5399 20213 5408 20247
rect 5356 20204 5408 20213
rect 14280 20204 14332 20256
rect 15200 20204 15252 20256
rect 19616 20204 19668 20256
rect 20168 20204 20220 20256
rect 7882 20102 7934 20154
rect 7946 20102 7998 20154
rect 8010 20102 8062 20154
rect 8074 20102 8126 20154
rect 14782 20102 14834 20154
rect 14846 20102 14898 20154
rect 14910 20102 14962 20154
rect 14974 20102 15026 20154
rect 3332 20043 3384 20052
rect 3332 20009 3341 20043
rect 3341 20009 3375 20043
rect 3375 20009 3384 20043
rect 3332 20000 3384 20009
rect 4160 20000 4212 20052
rect 4804 19864 4856 19916
rect 7472 20000 7524 20052
rect 8208 20000 8260 20052
rect 10416 20000 10468 20052
rect 16212 20043 16264 20052
rect 16212 20009 16221 20043
rect 16221 20009 16255 20043
rect 16255 20009 16264 20043
rect 16212 20000 16264 20009
rect 5356 19932 5408 19984
rect 6000 19975 6052 19984
rect 6000 19941 6009 19975
rect 6009 19941 6043 19975
rect 6043 19941 6052 19975
rect 6000 19932 6052 19941
rect 14464 19932 14516 19984
rect 15384 19932 15436 19984
rect 4988 19796 5040 19848
rect 5172 19907 5224 19916
rect 5172 19873 5207 19907
rect 5207 19873 5224 19907
rect 5172 19864 5224 19873
rect 7748 19907 7800 19916
rect 5080 19728 5132 19780
rect 5264 19728 5316 19780
rect 7748 19873 7757 19907
rect 7757 19873 7791 19907
rect 7791 19873 7800 19907
rect 7748 19864 7800 19873
rect 10324 19907 10376 19916
rect 7472 19796 7524 19848
rect 7656 19796 7708 19848
rect 10324 19873 10333 19907
rect 10333 19873 10367 19907
rect 10367 19873 10376 19907
rect 10324 19864 10376 19873
rect 12900 19864 12952 19916
rect 15108 19864 15160 19916
rect 15752 19864 15804 19916
rect 20536 19864 20588 19916
rect 15200 19796 15252 19848
rect 15384 19839 15436 19848
rect 15384 19805 15393 19839
rect 15393 19805 15427 19839
rect 15427 19805 15436 19839
rect 15384 19796 15436 19805
rect 16488 19728 16540 19780
rect 14648 19660 14700 19712
rect 20352 19660 20404 19712
rect 4432 19558 4484 19610
rect 4496 19558 4548 19610
rect 4560 19558 4612 19610
rect 4624 19558 4676 19610
rect 11332 19558 11384 19610
rect 11396 19558 11448 19610
rect 11460 19558 11512 19610
rect 11524 19558 11576 19610
rect 18232 19558 18284 19610
rect 18296 19558 18348 19610
rect 18360 19558 18412 19610
rect 18424 19558 18476 19610
rect 5264 19456 5316 19508
rect 15384 19456 15436 19508
rect 21088 19499 21140 19508
rect 21088 19465 21097 19499
rect 21097 19465 21131 19499
rect 21131 19465 21140 19499
rect 21088 19456 21140 19465
rect 14648 19363 14700 19372
rect 5172 19252 5224 19304
rect 5540 19252 5592 19304
rect 5632 19184 5684 19236
rect 5908 19252 5960 19304
rect 7380 19295 7432 19304
rect 7380 19261 7389 19295
rect 7389 19261 7423 19295
rect 7423 19261 7432 19295
rect 7380 19252 7432 19261
rect 6644 19184 6696 19236
rect 8484 19295 8536 19304
rect 8484 19261 8493 19295
rect 8493 19261 8527 19295
rect 8527 19261 8536 19295
rect 8484 19252 8536 19261
rect 7288 19116 7340 19168
rect 7656 19227 7708 19236
rect 7656 19193 7665 19227
rect 7665 19193 7699 19227
rect 7699 19193 7708 19227
rect 7656 19184 7708 19193
rect 7748 19116 7800 19168
rect 8944 19295 8996 19304
rect 8944 19261 8958 19295
rect 8958 19261 8992 19295
rect 8992 19261 8996 19295
rect 8944 19252 8996 19261
rect 8760 19227 8812 19236
rect 8760 19193 8769 19227
rect 8769 19193 8803 19227
rect 8803 19193 8812 19227
rect 8760 19184 8812 19193
rect 8852 19227 8904 19236
rect 8852 19193 8861 19227
rect 8861 19193 8895 19227
rect 8895 19193 8904 19227
rect 8852 19184 8904 19193
rect 13636 19252 13688 19304
rect 14648 19329 14657 19363
rect 14657 19329 14691 19363
rect 14691 19329 14700 19363
rect 14648 19320 14700 19329
rect 19616 19363 19668 19372
rect 14280 19252 14332 19304
rect 14556 19295 14608 19304
rect 14556 19261 14565 19295
rect 14565 19261 14599 19295
rect 14599 19261 14608 19295
rect 14556 19252 14608 19261
rect 14740 19295 14792 19304
rect 14740 19261 14749 19295
rect 14749 19261 14783 19295
rect 14783 19261 14792 19295
rect 14740 19252 14792 19261
rect 19616 19329 19625 19363
rect 19625 19329 19659 19363
rect 19659 19329 19668 19363
rect 19616 19320 19668 19329
rect 15200 19252 15252 19304
rect 17500 19252 17552 19304
rect 17776 19252 17828 19304
rect 19064 19252 19116 19304
rect 12808 19184 12860 19236
rect 9496 19116 9548 19168
rect 12624 19159 12676 19168
rect 12624 19125 12633 19159
rect 12633 19125 12667 19159
rect 12667 19125 12676 19159
rect 12624 19116 12676 19125
rect 12992 19116 13044 19168
rect 13636 19116 13688 19168
rect 15108 19184 15160 19236
rect 20352 19184 20404 19236
rect 17684 19116 17736 19168
rect 7882 19014 7934 19066
rect 7946 19014 7998 19066
rect 8010 19014 8062 19066
rect 8074 19014 8126 19066
rect 14782 19014 14834 19066
rect 14846 19014 14898 19066
rect 14910 19014 14962 19066
rect 14974 19014 15026 19066
rect 5540 18912 5592 18964
rect 5816 18912 5868 18964
rect 6644 18955 6696 18964
rect 6644 18921 6653 18955
rect 6653 18921 6687 18955
rect 6687 18921 6696 18955
rect 6644 18912 6696 18921
rect 8852 18912 8904 18964
rect 7288 18844 7340 18896
rect 5632 18819 5684 18828
rect 5632 18785 5641 18819
rect 5641 18785 5675 18819
rect 5675 18785 5684 18819
rect 5632 18776 5684 18785
rect 5356 18751 5408 18760
rect 5356 18717 5365 18751
rect 5365 18717 5399 18751
rect 5399 18717 5408 18751
rect 5356 18708 5408 18717
rect 5908 18708 5960 18760
rect 6736 18776 6788 18828
rect 7380 18776 7432 18828
rect 8944 18844 8996 18896
rect 12808 18844 12860 18896
rect 12992 18887 13044 18896
rect 12992 18853 13001 18887
rect 13001 18853 13035 18887
rect 13035 18853 13044 18887
rect 12992 18844 13044 18853
rect 8668 18776 8720 18828
rect 8760 18776 8812 18828
rect 12532 18819 12584 18828
rect 12532 18785 12541 18819
rect 12541 18785 12575 18819
rect 12575 18785 12584 18819
rect 12532 18776 12584 18785
rect 17684 18844 17736 18896
rect 19984 18844 20036 18896
rect 13728 18819 13780 18828
rect 13728 18785 13737 18819
rect 13737 18785 13771 18819
rect 13771 18785 13780 18819
rect 15476 18819 15528 18828
rect 13728 18776 13780 18785
rect 15476 18785 15485 18819
rect 15485 18785 15519 18819
rect 15519 18785 15528 18819
rect 15476 18776 15528 18785
rect 15660 18819 15712 18828
rect 15660 18785 15669 18819
rect 15669 18785 15703 18819
rect 15703 18785 15712 18819
rect 15660 18776 15712 18785
rect 16488 18776 16540 18828
rect 20352 18819 20404 18828
rect 8208 18708 8260 18760
rect 15752 18751 15804 18760
rect 15752 18717 15761 18751
rect 15761 18717 15795 18751
rect 15795 18717 15804 18751
rect 15752 18708 15804 18717
rect 16580 18708 16632 18760
rect 20352 18785 20361 18819
rect 20361 18785 20395 18819
rect 20395 18785 20404 18819
rect 20352 18776 20404 18785
rect 20536 18844 20588 18896
rect 16948 18708 17000 18760
rect 17316 18708 17368 18760
rect 5724 18640 5776 18692
rect 8484 18640 8536 18692
rect 9036 18640 9088 18692
rect 12532 18640 12584 18692
rect 16672 18640 16724 18692
rect 19156 18640 19208 18692
rect 7380 18572 7432 18624
rect 8576 18572 8628 18624
rect 13544 18615 13596 18624
rect 13544 18581 13553 18615
rect 13553 18581 13587 18615
rect 13587 18581 13596 18615
rect 13544 18572 13596 18581
rect 19064 18572 19116 18624
rect 20260 18572 20312 18624
rect 4432 18470 4484 18522
rect 4496 18470 4548 18522
rect 4560 18470 4612 18522
rect 4624 18470 4676 18522
rect 11332 18470 11384 18522
rect 11396 18470 11448 18522
rect 11460 18470 11512 18522
rect 11524 18470 11576 18522
rect 18232 18470 18284 18522
rect 18296 18470 18348 18522
rect 18360 18470 18412 18522
rect 18424 18470 18476 18522
rect 6644 18368 6696 18420
rect 15752 18368 15804 18420
rect 19064 18411 19116 18420
rect 19064 18377 19073 18411
rect 19073 18377 19107 18411
rect 19107 18377 19116 18411
rect 19064 18368 19116 18377
rect 2504 18232 2556 18284
rect 8576 18232 8628 18284
rect 9496 18275 9548 18284
rect 5724 18164 5776 18216
rect 6828 18164 6880 18216
rect 9496 18241 9505 18275
rect 9505 18241 9539 18275
rect 9539 18241 9548 18275
rect 9496 18232 9548 18241
rect 12992 18300 13044 18352
rect 13728 18300 13780 18352
rect 9680 18207 9732 18216
rect 3240 18096 3292 18148
rect 4252 18139 4304 18148
rect 4252 18105 4261 18139
rect 4261 18105 4295 18139
rect 4295 18105 4304 18139
rect 4252 18096 4304 18105
rect 5080 18096 5132 18148
rect 5632 18139 5684 18148
rect 5632 18105 5641 18139
rect 5641 18105 5675 18139
rect 5675 18105 5684 18139
rect 5632 18096 5684 18105
rect 8852 18096 8904 18148
rect 9680 18173 9689 18207
rect 9689 18173 9723 18207
rect 9723 18173 9732 18207
rect 9680 18164 9732 18173
rect 10324 18207 10376 18216
rect 10324 18173 10333 18207
rect 10333 18173 10367 18207
rect 10367 18173 10376 18207
rect 10324 18164 10376 18173
rect 10968 18164 11020 18216
rect 12624 18207 12676 18216
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 12624 18164 12676 18173
rect 16580 18232 16632 18284
rect 17224 18232 17276 18284
rect 20536 18300 20588 18352
rect 12992 18207 13044 18216
rect 12992 18173 13001 18207
rect 13001 18173 13035 18207
rect 13035 18173 13044 18207
rect 12992 18164 13044 18173
rect 13176 18207 13228 18216
rect 13176 18173 13185 18207
rect 13185 18173 13219 18207
rect 13219 18173 13228 18207
rect 13176 18164 13228 18173
rect 13544 18207 13596 18216
rect 13544 18173 13553 18207
rect 13553 18173 13587 18207
rect 13587 18173 13596 18207
rect 13544 18164 13596 18173
rect 17132 18164 17184 18216
rect 17316 18207 17368 18216
rect 17316 18173 17325 18207
rect 17325 18173 17359 18207
rect 17359 18173 17368 18207
rect 17316 18164 17368 18173
rect 19984 18232 20036 18284
rect 10232 18096 10284 18148
rect 19156 18164 19208 18216
rect 19616 18207 19668 18216
rect 19616 18173 19625 18207
rect 19625 18173 19659 18207
rect 19659 18173 19668 18207
rect 19616 18164 19668 18173
rect 20260 18164 20312 18216
rect 20628 18164 20680 18216
rect 4804 18028 4856 18080
rect 8484 18071 8536 18080
rect 8484 18037 8493 18071
rect 8493 18037 8527 18071
rect 8527 18037 8536 18071
rect 8484 18028 8536 18037
rect 8760 18028 8812 18080
rect 9772 18028 9824 18080
rect 10508 18071 10560 18080
rect 10508 18037 10517 18071
rect 10517 18037 10551 18071
rect 10551 18037 10560 18071
rect 10508 18028 10560 18037
rect 15660 18028 15712 18080
rect 17316 18028 17368 18080
rect 19616 18028 19668 18080
rect 20352 18028 20404 18080
rect 20996 18028 21048 18080
rect 7882 17926 7934 17978
rect 7946 17926 7998 17978
rect 8010 17926 8062 17978
rect 8074 17926 8126 17978
rect 14782 17926 14834 17978
rect 14846 17926 14898 17978
rect 14910 17926 14962 17978
rect 14974 17926 15026 17978
rect 3240 17824 3292 17876
rect 4252 17824 4304 17876
rect 13176 17824 13228 17876
rect 6092 17756 6144 17808
rect 7104 17756 7156 17808
rect 9772 17799 9824 17808
rect 9772 17765 9781 17799
rect 9781 17765 9815 17799
rect 9815 17765 9824 17799
rect 9772 17756 9824 17765
rect 10508 17756 10560 17808
rect 14648 17756 14700 17808
rect 15200 17756 15252 17808
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 4804 17731 4856 17740
rect 4804 17697 4813 17731
rect 4813 17697 4847 17731
rect 4847 17697 4856 17731
rect 4804 17688 4856 17697
rect 4988 17731 5040 17740
rect 4988 17697 4997 17731
rect 4997 17697 5031 17731
rect 5031 17697 5040 17731
rect 4988 17688 5040 17697
rect 5080 17731 5132 17740
rect 5080 17697 5115 17731
rect 5115 17697 5132 17731
rect 5080 17688 5132 17697
rect 5540 17688 5592 17740
rect 6644 17688 6696 17740
rect 6828 17731 6880 17740
rect 6828 17697 6837 17731
rect 6837 17697 6871 17731
rect 6871 17697 6880 17731
rect 6828 17688 6880 17697
rect 7748 17688 7800 17740
rect 8576 17688 8628 17740
rect 8944 17688 8996 17740
rect 9128 17688 9180 17740
rect 12164 17688 12216 17740
rect 12624 17688 12676 17740
rect 14464 17688 14516 17740
rect 15476 17688 15528 17740
rect 20904 17731 20956 17740
rect 20904 17697 20913 17731
rect 20913 17697 20947 17731
rect 20947 17697 20956 17731
rect 20904 17688 20956 17697
rect 4896 17620 4948 17672
rect 5264 17663 5316 17672
rect 5264 17629 5273 17663
rect 5273 17629 5307 17663
rect 5307 17629 5316 17663
rect 5264 17620 5316 17629
rect 7472 17620 7524 17672
rect 8392 17620 8444 17672
rect 12440 17620 12492 17672
rect 8484 17552 8536 17604
rect 1584 17527 1636 17536
rect 1584 17493 1593 17527
rect 1593 17493 1627 17527
rect 1627 17493 1636 17527
rect 1584 17484 1636 17493
rect 8300 17484 8352 17536
rect 8852 17484 8904 17536
rect 10140 17484 10192 17536
rect 12808 17552 12860 17604
rect 15936 17484 15988 17536
rect 20720 17527 20772 17536
rect 20720 17493 20729 17527
rect 20729 17493 20763 17527
rect 20763 17493 20772 17527
rect 20720 17484 20772 17493
rect 4432 17382 4484 17434
rect 4496 17382 4548 17434
rect 4560 17382 4612 17434
rect 4624 17382 4676 17434
rect 11332 17382 11384 17434
rect 11396 17382 11448 17434
rect 11460 17382 11512 17434
rect 11524 17382 11576 17434
rect 18232 17382 18284 17434
rect 18296 17382 18348 17434
rect 18360 17382 18412 17434
rect 18424 17382 18476 17434
rect 5816 17280 5868 17332
rect 7472 17323 7524 17332
rect 7472 17289 7481 17323
rect 7481 17289 7515 17323
rect 7515 17289 7524 17323
rect 7472 17280 7524 17289
rect 10232 17323 10284 17332
rect 10232 17289 10241 17323
rect 10241 17289 10275 17323
rect 10275 17289 10284 17323
rect 10232 17280 10284 17289
rect 12440 17280 12492 17332
rect 5540 17119 5592 17128
rect 5540 17085 5549 17119
rect 5549 17085 5583 17119
rect 5583 17085 5592 17119
rect 5540 17076 5592 17085
rect 5908 17212 5960 17264
rect 5724 17076 5776 17128
rect 5816 17008 5868 17060
rect 6736 17076 6788 17128
rect 7380 17212 7432 17264
rect 12532 17212 12584 17264
rect 7104 17187 7156 17196
rect 7104 17153 7113 17187
rect 7113 17153 7147 17187
rect 7147 17153 7156 17187
rect 7104 17144 7156 17153
rect 11060 17144 11112 17196
rect 12256 17144 12308 17196
rect 12624 17187 12676 17196
rect 7196 17119 7248 17128
rect 7196 17085 7205 17119
rect 7205 17085 7239 17119
rect 7239 17085 7248 17119
rect 7196 17076 7248 17085
rect 6644 17008 6696 17060
rect 8484 17076 8536 17128
rect 10140 17119 10192 17128
rect 10140 17085 10149 17119
rect 10149 17085 10183 17119
rect 10183 17085 10192 17119
rect 10140 17076 10192 17085
rect 12164 17076 12216 17128
rect 12624 17153 12633 17187
rect 12633 17153 12667 17187
rect 12667 17153 12676 17187
rect 12624 17144 12676 17153
rect 12808 17187 12860 17196
rect 12808 17153 12817 17187
rect 12817 17153 12851 17187
rect 12851 17153 12860 17187
rect 12808 17144 12860 17153
rect 15200 17280 15252 17332
rect 15936 17187 15988 17196
rect 15936 17153 15945 17187
rect 15945 17153 15979 17187
rect 15979 17153 15988 17187
rect 15936 17144 15988 17153
rect 16672 17144 16724 17196
rect 17040 17144 17092 17196
rect 17776 17144 17828 17196
rect 20720 17076 20772 17128
rect 10968 17008 11020 17060
rect 19616 17051 19668 17060
rect 5632 16940 5684 16992
rect 6552 16940 6604 16992
rect 8576 16940 8628 16992
rect 19616 17017 19625 17051
rect 19625 17017 19659 17051
rect 19659 17017 19668 17051
rect 19616 17008 19668 17017
rect 16212 16940 16264 16992
rect 17868 16940 17920 16992
rect 20260 16940 20312 16992
rect 7882 16838 7934 16890
rect 7946 16838 7998 16890
rect 8010 16838 8062 16890
rect 8074 16838 8126 16890
rect 14782 16838 14834 16890
rect 14846 16838 14898 16890
rect 14910 16838 14962 16890
rect 14974 16838 15026 16890
rect 6644 16779 6696 16788
rect 6644 16745 6653 16779
rect 6653 16745 6687 16779
rect 6687 16745 6696 16779
rect 6644 16736 6696 16745
rect 12440 16736 12492 16788
rect 14464 16736 14516 16788
rect 6920 16668 6972 16720
rect 5816 16643 5868 16652
rect 5816 16609 5825 16643
rect 5825 16609 5859 16643
rect 5859 16609 5868 16643
rect 5816 16600 5868 16609
rect 5908 16643 5960 16652
rect 5908 16609 5917 16643
rect 5917 16609 5951 16643
rect 5951 16609 5960 16643
rect 6552 16643 6604 16652
rect 5908 16600 5960 16609
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 6552 16600 6604 16609
rect 8300 16668 8352 16720
rect 14648 16668 14700 16720
rect 8852 16600 8904 16652
rect 12256 16600 12308 16652
rect 14924 16643 14976 16652
rect 14924 16609 14933 16643
rect 14933 16609 14967 16643
rect 14967 16609 14976 16643
rect 14924 16600 14976 16609
rect 15016 16600 15068 16652
rect 15200 16643 15252 16652
rect 15200 16609 15209 16643
rect 15209 16609 15243 16643
rect 15243 16609 15252 16643
rect 19248 16736 19300 16788
rect 19616 16736 19668 16788
rect 17224 16711 17276 16720
rect 17224 16677 17233 16711
rect 17233 16677 17267 16711
rect 17267 16677 17276 16711
rect 17224 16668 17276 16677
rect 15200 16600 15252 16609
rect 17132 16643 17184 16652
rect 6092 16575 6144 16584
rect 6092 16541 6101 16575
rect 6101 16541 6135 16575
rect 6135 16541 6144 16575
rect 6092 16532 6144 16541
rect 17132 16609 17141 16643
rect 17141 16609 17175 16643
rect 17175 16609 17184 16643
rect 17132 16600 17184 16609
rect 17316 16643 17368 16652
rect 17316 16609 17325 16643
rect 17325 16609 17359 16643
rect 17359 16609 17368 16643
rect 17316 16600 17368 16609
rect 17868 16600 17920 16652
rect 19524 16668 19576 16720
rect 20260 16711 20312 16720
rect 20260 16677 20269 16711
rect 20269 16677 20303 16711
rect 20303 16677 20312 16711
rect 20260 16668 20312 16677
rect 20168 16643 20220 16652
rect 19892 16532 19944 16584
rect 20168 16609 20177 16643
rect 20177 16609 20211 16643
rect 20211 16609 20220 16643
rect 20168 16600 20220 16609
rect 20076 16532 20128 16584
rect 20812 16532 20864 16584
rect 21180 16532 21232 16584
rect 13912 16396 13964 16448
rect 17592 16396 17644 16448
rect 18052 16396 18104 16448
rect 4432 16294 4484 16346
rect 4496 16294 4548 16346
rect 4560 16294 4612 16346
rect 4624 16294 4676 16346
rect 11332 16294 11384 16346
rect 11396 16294 11448 16346
rect 11460 16294 11512 16346
rect 11524 16294 11576 16346
rect 18232 16294 18284 16346
rect 18296 16294 18348 16346
rect 18360 16294 18412 16346
rect 18424 16294 18476 16346
rect 9680 16192 9732 16244
rect 12164 16235 12216 16244
rect 12164 16201 12173 16235
rect 12173 16201 12207 16235
rect 12207 16201 12216 16235
rect 12164 16192 12216 16201
rect 1952 15988 2004 16040
rect 2872 15988 2924 16040
rect 6828 16056 6880 16108
rect 6920 15988 6972 16040
rect 7196 16031 7248 16040
rect 7196 15997 7205 16031
rect 7205 15997 7239 16031
rect 7239 15997 7248 16031
rect 7196 15988 7248 15997
rect 7288 16031 7340 16040
rect 9036 16056 9088 16108
rect 12992 16056 13044 16108
rect 14924 16192 14976 16244
rect 19984 16235 20036 16244
rect 19984 16201 19993 16235
rect 19993 16201 20027 16235
rect 20027 16201 20036 16235
rect 19984 16192 20036 16201
rect 15108 16167 15160 16176
rect 15108 16133 15117 16167
rect 15117 16133 15151 16167
rect 15151 16133 15160 16167
rect 15108 16124 15160 16133
rect 19340 16124 19392 16176
rect 20168 16124 20220 16176
rect 7288 15997 7333 16031
rect 7333 15997 7340 16031
rect 7288 15988 7340 15997
rect 8576 16031 8628 16040
rect 8576 15997 8586 16031
rect 8586 15997 8620 16031
rect 8620 15997 8628 16031
rect 8852 16031 8904 16040
rect 8576 15988 8628 15997
rect 8852 15997 8861 16031
rect 8861 15997 8895 16031
rect 8895 15997 8904 16031
rect 8852 15988 8904 15997
rect 2688 15920 2740 15972
rect 8300 15920 8352 15972
rect 6276 15852 6328 15904
rect 8484 15852 8536 15904
rect 9864 16031 9916 16040
rect 9864 15997 9873 16031
rect 9873 15997 9907 16031
rect 9907 15997 9916 16031
rect 10968 16031 11020 16040
rect 9864 15988 9916 15997
rect 10968 15997 10977 16031
rect 10977 15997 11011 16031
rect 11011 15997 11020 16031
rect 10968 15988 11020 15997
rect 12348 16031 12400 16040
rect 12348 15997 12357 16031
rect 12357 15997 12391 16031
rect 12391 15997 12400 16031
rect 12348 15988 12400 15997
rect 12532 15988 12584 16040
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 15016 16056 15068 16108
rect 15200 15988 15252 16040
rect 17040 16056 17092 16108
rect 17592 16099 17644 16108
rect 17592 16065 17601 16099
rect 17601 16065 17635 16099
rect 17635 16065 17644 16099
rect 17592 16056 17644 16065
rect 19248 16056 19300 16108
rect 17132 15988 17184 16040
rect 19524 16031 19576 16040
rect 19524 15997 19533 16031
rect 19533 15997 19567 16031
rect 19567 15997 19576 16031
rect 19524 15988 19576 15997
rect 19800 16031 19852 16040
rect 19800 15997 19809 16031
rect 19809 15997 19843 16031
rect 19843 15997 19852 16031
rect 19800 15988 19852 15997
rect 18052 15920 18104 15972
rect 10232 15852 10284 15904
rect 11244 15852 11296 15904
rect 15200 15852 15252 15904
rect 19248 15852 19300 15904
rect 20536 15895 20588 15904
rect 20536 15861 20545 15895
rect 20545 15861 20579 15895
rect 20579 15861 20588 15895
rect 20536 15852 20588 15861
rect 7882 15750 7934 15802
rect 7946 15750 7998 15802
rect 8010 15750 8062 15802
rect 8074 15750 8126 15802
rect 14782 15750 14834 15802
rect 14846 15750 14898 15802
rect 14910 15750 14962 15802
rect 14974 15750 15026 15802
rect 7288 15648 7340 15700
rect 8484 15648 8536 15700
rect 5724 15580 5776 15632
rect 7196 15580 7248 15632
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 3240 15555 3292 15564
rect 3240 15521 3249 15555
rect 3249 15521 3283 15555
rect 3283 15521 3292 15555
rect 3240 15512 3292 15521
rect 1952 15444 2004 15496
rect 2872 15444 2924 15496
rect 6276 15487 6328 15496
rect 6276 15453 6285 15487
rect 6285 15453 6319 15487
rect 6319 15453 6328 15487
rect 6276 15444 6328 15453
rect 6920 15512 6972 15564
rect 7288 15512 7340 15564
rect 7472 15444 7524 15496
rect 8944 15580 8996 15632
rect 10232 15623 10284 15632
rect 10232 15589 10241 15623
rect 10241 15589 10275 15623
rect 10275 15589 10284 15623
rect 10232 15580 10284 15589
rect 11244 15580 11296 15632
rect 12348 15623 12400 15632
rect 12348 15589 12357 15623
rect 12357 15589 12391 15623
rect 12391 15589 12400 15623
rect 12348 15580 12400 15589
rect 12992 15580 13044 15632
rect 8300 15555 8352 15564
rect 8300 15521 8309 15555
rect 8309 15521 8343 15555
rect 8343 15521 8352 15555
rect 8300 15512 8352 15521
rect 9864 15512 9916 15564
rect 12532 15555 12584 15564
rect 12532 15521 12541 15555
rect 12541 15521 12575 15555
rect 12575 15521 12584 15555
rect 12532 15512 12584 15521
rect 17316 15648 17368 15700
rect 20444 15648 20496 15700
rect 19800 15580 19852 15632
rect 9128 15444 9180 15496
rect 13912 15512 13964 15564
rect 17132 15512 17184 15564
rect 17224 15512 17276 15564
rect 17684 15512 17736 15564
rect 19984 15555 20036 15564
rect 19984 15521 19993 15555
rect 19993 15521 20027 15555
rect 20027 15521 20036 15555
rect 19984 15512 20036 15521
rect 20168 15555 20220 15564
rect 20168 15521 20177 15555
rect 20177 15521 20211 15555
rect 20211 15521 20220 15555
rect 20168 15512 20220 15521
rect 20536 15555 20588 15564
rect 20536 15521 20545 15555
rect 20545 15521 20579 15555
rect 20579 15521 20588 15555
rect 20536 15512 20588 15521
rect 14556 15444 14608 15496
rect 2688 15376 2740 15428
rect 4988 15376 5040 15428
rect 9680 15376 9732 15428
rect 1860 15308 1912 15360
rect 4252 15351 4304 15360
rect 4252 15317 4261 15351
rect 4261 15317 4295 15351
rect 4295 15317 4304 15351
rect 4252 15308 4304 15317
rect 6368 15351 6420 15360
rect 6368 15317 6377 15351
rect 6377 15317 6411 15351
rect 6411 15317 6420 15351
rect 6368 15308 6420 15317
rect 10416 15308 10468 15360
rect 17776 15308 17828 15360
rect 4432 15206 4484 15258
rect 4496 15206 4548 15258
rect 4560 15206 4612 15258
rect 4624 15206 4676 15258
rect 11332 15206 11384 15258
rect 11396 15206 11448 15258
rect 11460 15206 11512 15258
rect 11524 15206 11576 15258
rect 18232 15206 18284 15258
rect 18296 15206 18348 15258
rect 18360 15206 18412 15258
rect 18424 15206 18476 15258
rect 1952 15104 2004 15156
rect 6828 15147 6880 15156
rect 6828 15113 6837 15147
rect 6837 15113 6871 15147
rect 6871 15113 6880 15147
rect 6828 15104 6880 15113
rect 7196 15104 7248 15156
rect 9864 15104 9916 15156
rect 12624 15104 12676 15156
rect 18880 15104 18932 15156
rect 19248 15104 19300 15156
rect 20352 15104 20404 15156
rect 4252 15079 4304 15088
rect 4252 15045 4261 15079
rect 4261 15045 4295 15079
rect 4295 15045 4304 15079
rect 4252 15036 4304 15045
rect 2044 15011 2096 15020
rect 2044 14977 2053 15011
rect 2053 14977 2087 15011
rect 2087 14977 2096 15011
rect 2044 14968 2096 14977
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 2872 14943 2924 14952
rect 2872 14909 2881 14943
rect 2881 14909 2915 14943
rect 2915 14909 2924 14943
rect 2872 14900 2924 14909
rect 4896 14900 4948 14952
rect 6828 14900 6880 14952
rect 8300 14968 8352 15020
rect 10232 14968 10284 15020
rect 7472 14900 7524 14952
rect 10416 14900 10468 14952
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 7564 14832 7616 14884
rect 12072 14832 12124 14884
rect 14648 14900 14700 14952
rect 15016 14943 15068 14952
rect 15016 14909 15025 14943
rect 15025 14909 15059 14943
rect 15059 14909 15068 14943
rect 15016 14900 15068 14909
rect 15384 14832 15436 14884
rect 19340 14900 19392 14952
rect 20260 14968 20312 15020
rect 19984 14943 20036 14952
rect 19984 14909 19993 14943
rect 19993 14909 20027 14943
rect 20027 14909 20036 14943
rect 19984 14900 20036 14909
rect 20168 14943 20220 14952
rect 20168 14909 20177 14943
rect 20177 14909 20211 14943
rect 20211 14909 20220 14943
rect 20168 14900 20220 14909
rect 21088 14943 21140 14952
rect 21088 14909 21097 14943
rect 21097 14909 21131 14943
rect 21131 14909 21140 14943
rect 21088 14900 21140 14909
rect 20444 14832 20496 14884
rect 3240 14764 3292 14816
rect 4804 14764 4856 14816
rect 12256 14764 12308 14816
rect 15200 14764 15252 14816
rect 16028 14764 16080 14816
rect 7882 14662 7934 14714
rect 7946 14662 7998 14714
rect 8010 14662 8062 14714
rect 8074 14662 8126 14714
rect 14782 14662 14834 14714
rect 14846 14662 14898 14714
rect 14910 14662 14962 14714
rect 14974 14662 15026 14714
rect 5540 14560 5592 14612
rect 6092 14560 6144 14612
rect 4804 14492 4856 14544
rect 6368 14492 6420 14544
rect 14556 14560 14608 14612
rect 8300 14492 8352 14544
rect 9128 14492 9180 14544
rect 14464 14492 14516 14544
rect 17224 14560 17276 14612
rect 20168 14603 20220 14612
rect 20168 14569 20177 14603
rect 20177 14569 20211 14603
rect 20211 14569 20220 14603
rect 20168 14560 20220 14569
rect 20260 14560 20312 14612
rect 6828 14424 6880 14476
rect 7196 14356 7248 14408
rect 8760 14356 8812 14408
rect 6828 14288 6880 14340
rect 5816 14220 5868 14272
rect 6644 14263 6696 14272
rect 6644 14229 6653 14263
rect 6653 14229 6687 14263
rect 6687 14229 6696 14263
rect 6644 14220 6696 14229
rect 6736 14220 6788 14272
rect 10324 14288 10376 14340
rect 14556 14424 14608 14476
rect 15200 14424 15252 14476
rect 15384 14467 15436 14476
rect 15384 14433 15393 14467
rect 15393 14433 15427 14467
rect 15427 14433 15436 14467
rect 15384 14424 15436 14433
rect 16028 14467 16080 14476
rect 16028 14433 16037 14467
rect 16037 14433 16071 14467
rect 16071 14433 16080 14467
rect 16028 14424 16080 14433
rect 18052 14424 18104 14476
rect 20444 14424 20496 14476
rect 14280 14288 14332 14340
rect 15476 14288 15528 14340
rect 17684 14288 17736 14340
rect 7472 14263 7524 14272
rect 7472 14229 7481 14263
rect 7481 14229 7515 14263
rect 7515 14229 7524 14263
rect 7472 14220 7524 14229
rect 17408 14263 17460 14272
rect 17408 14229 17417 14263
rect 17417 14229 17451 14263
rect 17451 14229 17460 14263
rect 17408 14220 17460 14229
rect 18696 14220 18748 14272
rect 20260 14220 20312 14272
rect 4432 14118 4484 14170
rect 4496 14118 4548 14170
rect 4560 14118 4612 14170
rect 4624 14118 4676 14170
rect 11332 14118 11384 14170
rect 11396 14118 11448 14170
rect 11460 14118 11512 14170
rect 11524 14118 11576 14170
rect 18232 14118 18284 14170
rect 18296 14118 18348 14170
rect 18360 14118 18412 14170
rect 18424 14118 18476 14170
rect 1952 14016 2004 14068
rect 8668 14016 8720 14068
rect 2872 13948 2924 14000
rect 6644 13948 6696 14000
rect 7288 13923 7340 13932
rect 7288 13889 7297 13923
rect 7297 13889 7331 13923
rect 7331 13889 7340 13923
rect 7288 13880 7340 13889
rect 5540 13812 5592 13864
rect 6736 13812 6788 13864
rect 6920 13812 6972 13864
rect 3332 13787 3384 13796
rect 3332 13753 3341 13787
rect 3341 13753 3375 13787
rect 3375 13753 3384 13787
rect 3332 13744 3384 13753
rect 7196 13855 7248 13864
rect 7196 13821 7205 13855
rect 7205 13821 7239 13855
rect 7239 13821 7248 13855
rect 7196 13812 7248 13821
rect 7656 13880 7708 13932
rect 10232 14059 10284 14068
rect 10232 14025 10241 14059
rect 10241 14025 10275 14059
rect 10275 14025 10284 14059
rect 10232 14016 10284 14025
rect 10324 14016 10376 14068
rect 9956 13948 10008 14000
rect 10140 13948 10192 14000
rect 7472 13812 7524 13864
rect 8576 13812 8628 13864
rect 9680 13880 9732 13932
rect 14464 13880 14516 13932
rect 9772 13855 9824 13864
rect 9772 13821 9781 13855
rect 9781 13821 9815 13855
rect 9815 13821 9824 13855
rect 9772 13812 9824 13821
rect 9404 13744 9456 13796
rect 10140 13812 10192 13864
rect 12164 13855 12216 13864
rect 12164 13821 12173 13855
rect 12173 13821 12207 13855
rect 12207 13821 12216 13855
rect 12164 13812 12216 13821
rect 12256 13855 12308 13864
rect 12256 13821 12265 13855
rect 12265 13821 12299 13855
rect 12299 13821 12308 13855
rect 14280 13855 14332 13864
rect 12256 13812 12308 13821
rect 14280 13821 14289 13855
rect 14289 13821 14323 13855
rect 14323 13821 14332 13855
rect 14280 13812 14332 13821
rect 14556 13812 14608 13864
rect 18144 13880 18196 13932
rect 18972 13923 19024 13932
rect 18972 13889 18981 13923
rect 18981 13889 19015 13923
rect 19015 13889 19024 13923
rect 18972 13880 19024 13889
rect 15200 13812 15252 13864
rect 17500 13855 17552 13864
rect 17500 13821 17509 13855
rect 17509 13821 17543 13855
rect 17543 13821 17552 13855
rect 17500 13812 17552 13821
rect 17684 13855 17736 13864
rect 17684 13821 17693 13855
rect 17693 13821 17727 13855
rect 17727 13821 17736 13855
rect 17684 13812 17736 13821
rect 17776 13855 17828 13864
rect 17776 13821 17785 13855
rect 17785 13821 17819 13855
rect 17819 13821 17828 13855
rect 17776 13812 17828 13821
rect 18052 13812 18104 13864
rect 18696 13855 18748 13864
rect 18696 13821 18705 13855
rect 18705 13821 18739 13855
rect 18739 13821 18748 13855
rect 18696 13812 18748 13821
rect 18880 13855 18932 13864
rect 18880 13821 18889 13855
rect 18889 13821 18923 13855
rect 18923 13821 18932 13855
rect 18880 13812 18932 13821
rect 20444 13880 20496 13932
rect 20628 13812 20680 13864
rect 20076 13744 20128 13796
rect 7656 13676 7708 13728
rect 12440 13719 12492 13728
rect 12440 13685 12449 13719
rect 12449 13685 12483 13719
rect 12483 13685 12492 13719
rect 14096 13719 14148 13728
rect 12440 13676 12492 13685
rect 14096 13685 14105 13719
rect 14105 13685 14139 13719
rect 14139 13685 14148 13719
rect 14096 13676 14148 13685
rect 17316 13719 17368 13728
rect 17316 13685 17325 13719
rect 17325 13685 17359 13719
rect 17359 13685 17368 13719
rect 17316 13676 17368 13685
rect 18604 13676 18656 13728
rect 7882 13574 7934 13626
rect 7946 13574 7998 13626
rect 8010 13574 8062 13626
rect 8074 13574 8126 13626
rect 14782 13574 14834 13626
rect 14846 13574 14898 13626
rect 14910 13574 14962 13626
rect 14974 13574 15026 13626
rect 1584 13472 1636 13524
rect 7104 13472 7156 13524
rect 7380 13515 7432 13524
rect 7380 13481 7389 13515
rect 7389 13481 7423 13515
rect 7423 13481 7432 13515
rect 7380 13472 7432 13481
rect 8392 13472 8444 13524
rect 18144 13515 18196 13524
rect 18144 13481 18153 13515
rect 18153 13481 18187 13515
rect 18187 13481 18196 13515
rect 18144 13472 18196 13481
rect 6092 13447 6144 13456
rect 6092 13413 6101 13447
rect 6101 13413 6135 13447
rect 6135 13413 6144 13447
rect 6092 13404 6144 13413
rect 6920 13404 6972 13456
rect 4896 13336 4948 13388
rect 6828 13336 6880 13388
rect 10048 13404 10100 13456
rect 12072 13447 12124 13456
rect 12072 13413 12081 13447
rect 12081 13413 12115 13447
rect 12115 13413 12124 13447
rect 12072 13404 12124 13413
rect 8208 13379 8260 13388
rect 8208 13345 8217 13379
rect 8217 13345 8251 13379
rect 8251 13345 8260 13379
rect 8208 13336 8260 13345
rect 8576 13336 8628 13388
rect 9496 13379 9548 13388
rect 9496 13345 9505 13379
rect 9505 13345 9539 13379
rect 9539 13345 9548 13379
rect 9496 13336 9548 13345
rect 9680 13379 9732 13388
rect 9680 13345 9689 13379
rect 9689 13345 9723 13379
rect 9723 13345 9732 13379
rect 9680 13336 9732 13345
rect 10232 13336 10284 13388
rect 2136 13268 2188 13320
rect 6184 13268 6236 13320
rect 12440 13404 12492 13456
rect 15200 13404 15252 13456
rect 17316 13404 17368 13456
rect 19892 13404 19944 13456
rect 16396 13336 16448 13388
rect 18052 13336 18104 13388
rect 13820 13268 13872 13320
rect 17040 13268 17092 13320
rect 17684 13311 17736 13320
rect 17684 13277 17693 13311
rect 17693 13277 17727 13311
rect 17727 13277 17736 13311
rect 17684 13268 17736 13277
rect 20076 13336 20128 13388
rect 20260 13379 20312 13388
rect 20260 13345 20269 13379
rect 20269 13345 20303 13379
rect 20303 13345 20312 13379
rect 20260 13336 20312 13345
rect 20444 13336 20496 13388
rect 13084 13200 13136 13252
rect 16304 13200 16356 13252
rect 2136 13132 2188 13184
rect 8668 13132 8720 13184
rect 9312 13132 9364 13184
rect 11060 13132 11112 13184
rect 11796 13132 11848 13184
rect 14188 13132 14240 13184
rect 17408 13132 17460 13184
rect 18880 13132 18932 13184
rect 19616 13132 19668 13184
rect 4432 13030 4484 13082
rect 4496 13030 4548 13082
rect 4560 13030 4612 13082
rect 4624 13030 4676 13082
rect 11332 13030 11384 13082
rect 11396 13030 11448 13082
rect 11460 13030 11512 13082
rect 11524 13030 11576 13082
rect 18232 13030 18284 13082
rect 18296 13030 18348 13082
rect 18360 13030 18412 13082
rect 18424 13030 18476 13082
rect 1492 12971 1544 12980
rect 1492 12937 1501 12971
rect 1501 12937 1535 12971
rect 1535 12937 1544 12971
rect 1492 12928 1544 12937
rect 3332 12928 3384 12980
rect 4896 12971 4948 12980
rect 4896 12937 4905 12971
rect 4905 12937 4939 12971
rect 4939 12937 4948 12971
rect 4896 12928 4948 12937
rect 9772 12928 9824 12980
rect 10048 12971 10100 12980
rect 10048 12937 10057 12971
rect 10057 12937 10091 12971
rect 10091 12937 10100 12971
rect 10048 12928 10100 12937
rect 10324 12928 10376 12980
rect 11704 12928 11756 12980
rect 12256 12928 12308 12980
rect 14556 12928 14608 12980
rect 16396 12971 16448 12980
rect 16396 12937 16405 12971
rect 16405 12937 16439 12971
rect 16439 12937 16448 12971
rect 16396 12928 16448 12937
rect 17500 12928 17552 12980
rect 20260 12928 20312 12980
rect 6828 12860 6880 12912
rect 9404 12860 9456 12912
rect 17684 12860 17736 12912
rect 2136 12767 2188 12776
rect 2136 12733 2145 12767
rect 2145 12733 2179 12767
rect 2179 12733 2188 12767
rect 2136 12724 2188 12733
rect 2780 12724 2832 12776
rect 3332 12724 3384 12776
rect 5172 12767 5224 12776
rect 5172 12733 5181 12767
rect 5181 12733 5215 12767
rect 5215 12733 5224 12767
rect 5172 12724 5224 12733
rect 3240 12656 3292 12708
rect 4988 12656 5040 12708
rect 7196 12724 7248 12776
rect 7380 12724 7432 12776
rect 8392 12724 8444 12776
rect 8944 12767 8996 12776
rect 8944 12733 8953 12767
rect 8953 12733 8987 12767
rect 8987 12733 8996 12767
rect 8944 12724 8996 12733
rect 9680 12767 9732 12776
rect 9680 12733 9689 12767
rect 9689 12733 9723 12767
rect 9723 12733 9732 12767
rect 9680 12724 9732 12733
rect 9956 12724 10008 12776
rect 10140 12767 10192 12776
rect 10140 12733 10149 12767
rect 10149 12733 10183 12767
rect 10183 12733 10192 12767
rect 10140 12724 10192 12733
rect 10600 12724 10652 12776
rect 12072 12792 12124 12844
rect 12348 12792 12400 12844
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 17408 12792 17460 12844
rect 18880 12792 18932 12844
rect 19616 12835 19668 12844
rect 19616 12801 19625 12835
rect 19625 12801 19659 12835
rect 19659 12801 19668 12835
rect 19616 12792 19668 12801
rect 11060 12767 11112 12776
rect 11060 12733 11069 12767
rect 11069 12733 11103 12767
rect 11103 12733 11112 12767
rect 11060 12724 11112 12733
rect 13084 12767 13136 12776
rect 13084 12733 13093 12767
rect 13093 12733 13127 12767
rect 13127 12733 13136 12767
rect 13084 12724 13136 12733
rect 16212 12767 16264 12776
rect 16212 12733 16221 12767
rect 16221 12733 16255 12767
rect 16255 12733 16264 12767
rect 16212 12724 16264 12733
rect 18052 12724 18104 12776
rect 18604 12724 18656 12776
rect 6920 12656 6972 12708
rect 7656 12656 7708 12708
rect 8208 12588 8260 12640
rect 9220 12588 9272 12640
rect 12624 12631 12676 12640
rect 12624 12597 12633 12631
rect 12633 12597 12667 12631
rect 12667 12597 12676 12631
rect 12624 12588 12676 12597
rect 12992 12631 13044 12640
rect 12992 12597 13001 12631
rect 13001 12597 13035 12631
rect 13035 12597 13044 12631
rect 12992 12588 13044 12597
rect 15108 12656 15160 12708
rect 17776 12656 17828 12708
rect 20628 12656 20680 12708
rect 17960 12588 18012 12640
rect 18880 12631 18932 12640
rect 18880 12597 18889 12631
rect 18889 12597 18923 12631
rect 18923 12597 18932 12631
rect 18880 12588 18932 12597
rect 7882 12486 7934 12538
rect 7946 12486 7998 12538
rect 8010 12486 8062 12538
rect 8074 12486 8126 12538
rect 14782 12486 14834 12538
rect 14846 12486 14898 12538
rect 14910 12486 14962 12538
rect 14974 12486 15026 12538
rect 5540 12427 5592 12436
rect 5540 12393 5549 12427
rect 5549 12393 5583 12427
rect 5583 12393 5592 12427
rect 5540 12384 5592 12393
rect 11060 12384 11112 12436
rect 12164 12384 12216 12436
rect 12992 12384 13044 12436
rect 15108 12384 15160 12436
rect 20628 12427 20680 12436
rect 20628 12393 20637 12427
rect 20637 12393 20671 12427
rect 20671 12393 20680 12427
rect 20628 12384 20680 12393
rect 3332 12359 3384 12368
rect 3332 12325 3341 12359
rect 3341 12325 3375 12359
rect 3375 12325 3384 12359
rect 3332 12316 3384 12325
rect 11796 12359 11848 12368
rect 11796 12325 11805 12359
rect 11805 12325 11839 12359
rect 11839 12325 11848 12359
rect 11796 12316 11848 12325
rect 2964 12248 3016 12300
rect 5172 12248 5224 12300
rect 5724 12248 5776 12300
rect 6920 12248 6972 12300
rect 7564 12291 7616 12300
rect 7564 12257 7573 12291
rect 7573 12257 7607 12291
rect 7607 12257 7616 12291
rect 7564 12248 7616 12257
rect 5908 12180 5960 12232
rect 6828 12180 6880 12232
rect 8208 12180 8260 12232
rect 10416 12180 10468 12232
rect 16212 12248 16264 12300
rect 20076 12248 20128 12300
rect 20904 12248 20956 12300
rect 5080 12087 5132 12096
rect 5080 12053 5089 12087
rect 5089 12053 5123 12087
rect 5123 12053 5132 12087
rect 5080 12044 5132 12053
rect 5632 12044 5684 12096
rect 6736 12112 6788 12164
rect 7472 12112 7524 12164
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 4432 11942 4484 11994
rect 4496 11942 4548 11994
rect 4560 11942 4612 11994
rect 4624 11942 4676 11994
rect 11332 11942 11384 11994
rect 11396 11942 11448 11994
rect 11460 11942 11512 11994
rect 11524 11942 11576 11994
rect 18232 11942 18284 11994
rect 18296 11942 18348 11994
rect 18360 11942 18412 11994
rect 18424 11942 18476 11994
rect 2964 11883 3016 11892
rect 2964 11849 2973 11883
rect 2973 11849 3007 11883
rect 3007 11849 3016 11883
rect 2964 11840 3016 11849
rect 5724 11747 5776 11756
rect 5724 11713 5733 11747
rect 5733 11713 5767 11747
rect 5767 11713 5776 11747
rect 5724 11704 5776 11713
rect 6000 11704 6052 11756
rect 6828 11747 6880 11756
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 2780 11636 2832 11688
rect 3516 11679 3568 11688
rect 3516 11645 3525 11679
rect 3525 11645 3559 11679
rect 3559 11645 3568 11679
rect 3516 11636 3568 11645
rect 5632 11679 5684 11688
rect 5632 11645 5641 11679
rect 5641 11645 5675 11679
rect 5675 11645 5684 11679
rect 7380 11840 7432 11892
rect 8208 11840 8260 11892
rect 9220 11840 9272 11892
rect 7656 11704 7708 11756
rect 8944 11704 8996 11756
rect 5632 11636 5684 11645
rect 9312 11679 9364 11688
rect 4068 11568 4120 11620
rect 5264 11568 5316 11620
rect 7288 11568 7340 11620
rect 7748 11568 7800 11620
rect 9312 11645 9321 11679
rect 9321 11645 9355 11679
rect 9355 11645 9364 11679
rect 9312 11636 9364 11645
rect 10324 11704 10376 11756
rect 4988 11500 5040 11552
rect 9680 11568 9732 11620
rect 9772 11543 9824 11552
rect 9772 11509 9781 11543
rect 9781 11509 9815 11543
rect 9815 11509 9824 11543
rect 9772 11500 9824 11509
rect 18420 11500 18472 11552
rect 7882 11398 7934 11450
rect 7946 11398 7998 11450
rect 8010 11398 8062 11450
rect 8074 11398 8126 11450
rect 14782 11398 14834 11450
rect 14846 11398 14898 11450
rect 14910 11398 14962 11450
rect 14974 11398 15026 11450
rect 1860 11296 1912 11348
rect 2964 11339 3016 11348
rect 2964 11305 2973 11339
rect 2973 11305 3007 11339
rect 3007 11305 3016 11339
rect 2964 11296 3016 11305
rect 4252 11228 4304 11280
rect 9772 11296 9824 11348
rect 12716 11296 12768 11348
rect 5632 11228 5684 11280
rect 2228 11135 2280 11144
rect 2228 11101 2237 11135
rect 2237 11101 2271 11135
rect 2271 11101 2280 11135
rect 2228 11092 2280 11101
rect 3516 11092 3568 11144
rect 4068 11092 4120 11144
rect 5540 11160 5592 11212
rect 5908 11160 5960 11212
rect 9680 11228 9732 11280
rect 10048 11271 10100 11280
rect 10048 11237 10057 11271
rect 10057 11237 10091 11271
rect 10091 11237 10100 11271
rect 10048 11228 10100 11237
rect 10416 11228 10468 11280
rect 11704 11228 11756 11280
rect 6828 11160 6880 11212
rect 7104 11160 7156 11212
rect 7656 11160 7708 11212
rect 8208 11160 8260 11212
rect 6000 11092 6052 11144
rect 7380 11092 7432 11144
rect 15016 11203 15068 11212
rect 15016 11169 15025 11203
rect 15025 11169 15059 11203
rect 15059 11169 15068 11203
rect 15016 11160 15068 11169
rect 7288 11024 7340 11076
rect 10416 11067 10468 11076
rect 10416 11033 10425 11067
rect 10425 11033 10459 11067
rect 10459 11033 10468 11067
rect 10416 11024 10468 11033
rect 10600 11024 10652 11076
rect 12348 11092 12400 11144
rect 18144 11228 18196 11280
rect 20996 11296 21048 11348
rect 20904 11228 20956 11280
rect 16948 11203 17000 11212
rect 16948 11169 16957 11203
rect 16957 11169 16991 11203
rect 16991 11169 17000 11203
rect 16948 11160 17000 11169
rect 18420 11203 18472 11212
rect 16488 11092 16540 11144
rect 18420 11169 18429 11203
rect 18429 11169 18463 11203
rect 18463 11169 18472 11203
rect 18420 11160 18472 11169
rect 20076 11203 20128 11212
rect 20076 11169 20085 11203
rect 20085 11169 20119 11203
rect 20119 11169 20128 11203
rect 20076 11160 20128 11169
rect 18328 11092 18380 11144
rect 18604 11135 18656 11144
rect 18604 11101 18613 11135
rect 18613 11101 18647 11135
rect 18647 11101 18656 11135
rect 18604 11092 18656 11101
rect 14832 11024 14884 11076
rect 15200 11067 15252 11076
rect 15200 11033 15209 11067
rect 15209 11033 15243 11067
rect 15243 11033 15252 11067
rect 15200 11024 15252 11033
rect 18052 11067 18104 11076
rect 1584 10999 1636 11008
rect 1584 10965 1593 10999
rect 1593 10965 1627 10999
rect 1627 10965 1636 10999
rect 1584 10956 1636 10965
rect 5908 10999 5960 11008
rect 5908 10965 5917 10999
rect 5917 10965 5951 10999
rect 5951 10965 5960 10999
rect 5908 10956 5960 10965
rect 9864 10956 9916 11008
rect 10232 10999 10284 11008
rect 10232 10965 10241 10999
rect 10241 10965 10275 10999
rect 10275 10965 10284 10999
rect 10232 10956 10284 10965
rect 16856 10999 16908 11008
rect 16856 10965 16865 10999
rect 16865 10965 16899 10999
rect 16899 10965 16908 10999
rect 16856 10956 16908 10965
rect 18052 11033 18061 11067
rect 18061 11033 18095 11067
rect 18095 11033 18104 11067
rect 18052 11024 18104 11033
rect 20168 11024 20220 11076
rect 18696 10956 18748 11008
rect 4432 10854 4484 10906
rect 4496 10854 4548 10906
rect 4560 10854 4612 10906
rect 4624 10854 4676 10906
rect 11332 10854 11384 10906
rect 11396 10854 11448 10906
rect 11460 10854 11512 10906
rect 11524 10854 11576 10906
rect 18232 10854 18284 10906
rect 18296 10854 18348 10906
rect 18360 10854 18412 10906
rect 18424 10854 18476 10906
rect 4252 10752 4304 10804
rect 4896 10752 4948 10804
rect 7564 10795 7616 10804
rect 7564 10761 7573 10795
rect 7573 10761 7607 10795
rect 7607 10761 7616 10795
rect 7564 10752 7616 10761
rect 13820 10752 13872 10804
rect 15016 10752 15068 10804
rect 20444 10752 20496 10804
rect 7656 10684 7708 10736
rect 16856 10684 16908 10736
rect 5632 10616 5684 10668
rect 2688 10591 2740 10600
rect 2688 10557 2697 10591
rect 2697 10557 2731 10591
rect 2731 10557 2740 10591
rect 2688 10548 2740 10557
rect 5264 10548 5316 10600
rect 7748 10548 7800 10600
rect 9680 10616 9732 10668
rect 12624 10616 12676 10668
rect 18604 10616 18656 10668
rect 18880 10616 18932 10668
rect 9496 10548 9548 10600
rect 13452 10591 13504 10600
rect 13452 10557 13461 10591
rect 13461 10557 13495 10591
rect 13495 10557 13504 10591
rect 13452 10548 13504 10557
rect 14832 10591 14884 10600
rect 14832 10557 14841 10591
rect 14841 10557 14875 10591
rect 14875 10557 14884 10591
rect 14832 10548 14884 10557
rect 15200 10548 15252 10600
rect 17684 10548 17736 10600
rect 17960 10548 18012 10600
rect 2044 10480 2096 10532
rect 2872 10523 2924 10532
rect 2872 10489 2881 10523
rect 2881 10489 2915 10523
rect 2915 10489 2924 10523
rect 2872 10480 2924 10489
rect 8484 10523 8536 10532
rect 8484 10489 8493 10523
rect 8493 10489 8527 10523
rect 8527 10489 8536 10523
rect 8484 10480 8536 10489
rect 1492 10455 1544 10464
rect 1492 10421 1501 10455
rect 1501 10421 1535 10455
rect 1535 10421 1544 10455
rect 1492 10412 1544 10421
rect 7656 10412 7708 10464
rect 8576 10412 8628 10464
rect 9588 10412 9640 10464
rect 17408 10480 17460 10532
rect 20168 10480 20220 10532
rect 17316 10412 17368 10464
rect 17776 10412 17828 10464
rect 18788 10412 18840 10464
rect 7882 10310 7934 10362
rect 7946 10310 7998 10362
rect 8010 10310 8062 10362
rect 8074 10310 8126 10362
rect 14782 10310 14834 10362
rect 14846 10310 14898 10362
rect 14910 10310 14962 10362
rect 14974 10310 15026 10362
rect 2228 10251 2280 10260
rect 2228 10217 2237 10251
rect 2237 10217 2271 10251
rect 2271 10217 2280 10251
rect 2228 10208 2280 10217
rect 5356 10208 5408 10260
rect 7012 10208 7064 10260
rect 7380 10208 7432 10260
rect 12440 10208 12492 10260
rect 20904 10251 20956 10260
rect 5908 10140 5960 10192
rect 1584 10072 1636 10124
rect 8208 10072 8260 10124
rect 9220 10140 9272 10192
rect 8576 10115 8628 10124
rect 8576 10081 8585 10115
rect 8585 10081 8619 10115
rect 8619 10081 8628 10115
rect 8576 10072 8628 10081
rect 9404 10072 9456 10124
rect 13820 10140 13872 10192
rect 16948 10140 17000 10192
rect 20904 10217 20913 10251
rect 20913 10217 20947 10251
rect 20947 10217 20956 10251
rect 20904 10208 20956 10217
rect 12624 10072 12676 10124
rect 12992 10072 13044 10124
rect 16488 10072 16540 10124
rect 17776 10115 17828 10124
rect 17776 10081 17785 10115
rect 17785 10081 17819 10115
rect 17819 10081 17828 10115
rect 17776 10072 17828 10081
rect 21088 10115 21140 10124
rect 21088 10081 21097 10115
rect 21097 10081 21131 10115
rect 21131 10081 21140 10115
rect 21088 10072 21140 10081
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 9772 10047 9824 10056
rect 9772 10013 9781 10047
rect 9781 10013 9815 10047
rect 9815 10013 9824 10047
rect 9772 10004 9824 10013
rect 11152 10004 11204 10056
rect 18696 10004 18748 10056
rect 2780 9936 2832 9988
rect 10232 9936 10284 9988
rect 11888 9979 11940 9988
rect 11888 9945 11897 9979
rect 11897 9945 11931 9979
rect 11931 9945 11940 9979
rect 11888 9936 11940 9945
rect 6184 9868 6236 9920
rect 8760 9868 8812 9920
rect 13360 9868 13412 9920
rect 4432 9766 4484 9818
rect 4496 9766 4548 9818
rect 4560 9766 4612 9818
rect 4624 9766 4676 9818
rect 11332 9766 11384 9818
rect 11396 9766 11448 9818
rect 11460 9766 11512 9818
rect 11524 9766 11576 9818
rect 18232 9766 18284 9818
rect 18296 9766 18348 9818
rect 18360 9766 18412 9818
rect 18424 9766 18476 9818
rect 2228 9664 2280 9716
rect 13452 9664 13504 9716
rect 2780 9639 2832 9648
rect 2780 9605 2789 9639
rect 2789 9605 2823 9639
rect 2823 9605 2832 9639
rect 2780 9596 2832 9605
rect 11152 9596 11204 9648
rect 7196 9528 7248 9580
rect 1584 9460 1636 9512
rect 2872 9460 2924 9512
rect 4988 9503 5040 9512
rect 4988 9469 4997 9503
rect 4997 9469 5031 9503
rect 5031 9469 5040 9503
rect 4988 9460 5040 9469
rect 7564 9503 7616 9512
rect 7564 9469 7573 9503
rect 7573 9469 7607 9503
rect 7607 9469 7616 9503
rect 7564 9460 7616 9469
rect 2412 9392 2464 9444
rect 5172 9392 5224 9444
rect 5448 9392 5500 9444
rect 8484 9460 8536 9512
rect 10508 9528 10560 9580
rect 12440 9571 12492 9580
rect 12440 9537 12449 9571
rect 12449 9537 12483 9571
rect 12483 9537 12492 9571
rect 12440 9528 12492 9537
rect 12992 9460 13044 9512
rect 14280 9503 14332 9512
rect 14280 9469 14289 9503
rect 14289 9469 14323 9503
rect 14323 9469 14332 9503
rect 14280 9460 14332 9469
rect 9680 9392 9732 9444
rect 12348 9392 12400 9444
rect 4804 9367 4856 9376
rect 4804 9333 4813 9367
rect 4813 9333 4847 9367
rect 4847 9333 4856 9367
rect 4804 9324 4856 9333
rect 9956 9324 10008 9376
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10140 9324 10192 9333
rect 15200 9324 15252 9376
rect 7882 9222 7934 9274
rect 7946 9222 7998 9274
rect 8010 9222 8062 9274
rect 8074 9222 8126 9274
rect 14782 9222 14834 9274
rect 14846 9222 14898 9274
rect 14910 9222 14962 9274
rect 14974 9222 15026 9274
rect 2228 9120 2280 9172
rect 9956 9163 10008 9172
rect 1400 9052 1452 9104
rect 5540 9052 5592 9104
rect 5816 9095 5868 9104
rect 5816 9061 5825 9095
rect 5825 9061 5859 9095
rect 5859 9061 5868 9095
rect 5816 9052 5868 9061
rect 6000 9095 6052 9104
rect 6000 9061 6009 9095
rect 6009 9061 6043 9095
rect 6043 9061 6052 9095
rect 6000 9052 6052 9061
rect 2504 8848 2556 8900
rect 4988 9027 5040 9036
rect 4988 8993 4997 9027
rect 4997 8993 5031 9027
rect 5031 8993 5040 9027
rect 4988 8984 5040 8993
rect 6920 8984 6972 9036
rect 9956 9129 9965 9163
rect 9965 9129 9999 9163
rect 9999 9129 10008 9163
rect 9956 9120 10008 9129
rect 11888 9120 11940 9172
rect 15200 9163 15252 9172
rect 15200 9129 15209 9163
rect 15209 9129 15243 9163
rect 15243 9129 15252 9163
rect 15200 9120 15252 9129
rect 15292 9163 15344 9172
rect 15292 9129 15301 9163
rect 15301 9129 15335 9163
rect 15335 9129 15344 9163
rect 18604 9163 18656 9172
rect 15292 9120 15344 9129
rect 18604 9129 18613 9163
rect 18613 9129 18647 9163
rect 18647 9129 18656 9163
rect 18604 9120 18656 9129
rect 17316 9095 17368 9104
rect 17316 9061 17325 9095
rect 17325 9061 17359 9095
rect 17359 9061 17368 9095
rect 17316 9052 17368 9061
rect 8392 8984 8444 9036
rect 9588 9027 9640 9036
rect 9588 8993 9597 9027
rect 9597 8993 9631 9027
rect 9631 8993 9640 9027
rect 9588 8984 9640 8993
rect 10048 8984 10100 9036
rect 10692 8984 10744 9036
rect 12992 8984 13044 9036
rect 14464 8984 14516 9036
rect 5724 8959 5776 8968
rect 5724 8925 5733 8959
rect 5733 8925 5767 8959
rect 5767 8925 5776 8959
rect 5724 8916 5776 8925
rect 7564 8916 7616 8968
rect 12624 8916 12676 8968
rect 16580 8959 16632 8968
rect 16580 8925 16589 8959
rect 16589 8925 16623 8959
rect 16623 8925 16632 8959
rect 16580 8916 16632 8925
rect 18052 8984 18104 9036
rect 18696 8916 18748 8968
rect 7656 8848 7708 8900
rect 9772 8848 9824 8900
rect 19156 8848 19208 8900
rect 3884 8780 3936 8832
rect 6276 8823 6328 8832
rect 6276 8789 6285 8823
rect 6285 8789 6319 8823
rect 6319 8789 6328 8823
rect 6276 8780 6328 8789
rect 7748 8780 7800 8832
rect 14648 8780 14700 8832
rect 4432 8678 4484 8730
rect 4496 8678 4548 8730
rect 4560 8678 4612 8730
rect 4624 8678 4676 8730
rect 11332 8678 11384 8730
rect 11396 8678 11448 8730
rect 11460 8678 11512 8730
rect 11524 8678 11576 8730
rect 18232 8678 18284 8730
rect 18296 8678 18348 8730
rect 18360 8678 18412 8730
rect 18424 8678 18476 8730
rect 2136 8619 2188 8628
rect 2136 8585 2145 8619
rect 2145 8585 2179 8619
rect 2179 8585 2188 8619
rect 2136 8576 2188 8585
rect 4988 8576 5040 8628
rect 9588 8619 9640 8628
rect 9588 8585 9597 8619
rect 9597 8585 9631 8619
rect 9631 8585 9640 8619
rect 9588 8576 9640 8585
rect 16580 8576 16632 8628
rect 18604 8576 18656 8628
rect 19156 8619 19208 8628
rect 19156 8585 19165 8619
rect 19165 8585 19199 8619
rect 19199 8585 19208 8619
rect 19156 8576 19208 8585
rect 6276 8508 6328 8560
rect 14464 8508 14516 8560
rect 3884 8483 3936 8492
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 2504 8415 2556 8424
rect 2504 8381 2513 8415
rect 2513 8381 2547 8415
rect 2547 8381 2556 8415
rect 2504 8372 2556 8381
rect 2412 8304 2464 8356
rect 3884 8449 3893 8483
rect 3893 8449 3927 8483
rect 3927 8449 3936 8483
rect 3884 8440 3936 8449
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 9772 8440 9824 8492
rect 14188 8483 14240 8492
rect 10048 8372 10100 8424
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 3792 8347 3844 8356
rect 3792 8313 3801 8347
rect 3801 8313 3835 8347
rect 3835 8313 3844 8347
rect 3792 8304 3844 8313
rect 8392 8304 8444 8356
rect 9220 8304 9272 8356
rect 14280 8372 14332 8424
rect 15292 8372 15344 8424
rect 18052 8372 18104 8424
rect 18144 8415 18196 8424
rect 18144 8381 18153 8415
rect 18153 8381 18187 8415
rect 18187 8381 18196 8415
rect 18696 8415 18748 8424
rect 18144 8372 18196 8381
rect 18696 8381 18705 8415
rect 18705 8381 18739 8415
rect 18739 8381 18748 8415
rect 18696 8372 18748 8381
rect 21088 8415 21140 8424
rect 21088 8381 21097 8415
rect 21097 8381 21131 8415
rect 21131 8381 21140 8415
rect 21088 8372 21140 8381
rect 12348 8304 12400 8356
rect 12624 8304 12676 8356
rect 9864 8279 9916 8288
rect 9864 8245 9873 8279
rect 9873 8245 9907 8279
rect 9907 8245 9916 8279
rect 9864 8236 9916 8245
rect 12440 8279 12492 8288
rect 12440 8245 12449 8279
rect 12449 8245 12483 8279
rect 12483 8245 12492 8279
rect 14556 8279 14608 8288
rect 12440 8236 12492 8245
rect 14556 8245 14565 8279
rect 14565 8245 14599 8279
rect 14599 8245 14608 8279
rect 14556 8236 14608 8245
rect 20904 8279 20956 8288
rect 20904 8245 20913 8279
rect 20913 8245 20947 8279
rect 20947 8245 20956 8279
rect 20904 8236 20956 8245
rect 7882 8134 7934 8186
rect 7946 8134 7998 8186
rect 8010 8134 8062 8186
rect 8074 8134 8126 8186
rect 14782 8134 14834 8186
rect 14846 8134 14898 8186
rect 14910 8134 14962 8186
rect 14974 8134 15026 8186
rect 12440 8032 12492 8084
rect 18604 8032 18656 8084
rect 8300 7964 8352 8016
rect 14556 7964 14608 8016
rect 16580 7964 16632 8016
rect 18052 7964 18104 8016
rect 2136 7939 2188 7948
rect 2136 7905 2145 7939
rect 2145 7905 2179 7939
rect 2179 7905 2188 7939
rect 2136 7896 2188 7905
rect 2688 7939 2740 7948
rect 2688 7905 2697 7939
rect 2697 7905 2731 7939
rect 2731 7905 2740 7939
rect 2688 7896 2740 7905
rect 7748 7939 7800 7948
rect 7748 7905 7757 7939
rect 7757 7905 7791 7939
rect 7791 7905 7800 7939
rect 7748 7896 7800 7905
rect 10324 7896 10376 7948
rect 14188 7896 14240 7948
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 12624 7871 12676 7880
rect 12624 7837 12633 7871
rect 12633 7837 12667 7871
rect 12667 7837 12676 7871
rect 12624 7828 12676 7837
rect 20904 7828 20956 7880
rect 3792 7692 3844 7744
rect 9496 7692 9548 7744
rect 13268 7692 13320 7744
rect 4432 7590 4484 7642
rect 4496 7590 4548 7642
rect 4560 7590 4612 7642
rect 4624 7590 4676 7642
rect 11332 7590 11384 7642
rect 11396 7590 11448 7642
rect 11460 7590 11512 7642
rect 11524 7590 11576 7642
rect 18232 7590 18284 7642
rect 18296 7590 18348 7642
rect 18360 7590 18412 7642
rect 18424 7590 18476 7642
rect 4068 7488 4120 7540
rect 13452 7488 13504 7540
rect 4252 7352 4304 7404
rect 5080 7352 5132 7404
rect 13268 7395 13320 7404
rect 7748 7327 7800 7336
rect 7748 7293 7757 7327
rect 7757 7293 7791 7327
rect 7791 7293 7800 7327
rect 7748 7284 7800 7293
rect 9496 7327 9548 7336
rect 9496 7293 9505 7327
rect 9505 7293 9539 7327
rect 9539 7293 9548 7327
rect 9496 7284 9548 7293
rect 10692 7327 10744 7336
rect 10692 7293 10701 7327
rect 10701 7293 10735 7327
rect 10735 7293 10744 7327
rect 10692 7284 10744 7293
rect 13268 7361 13277 7395
rect 13277 7361 13311 7395
rect 13311 7361 13320 7395
rect 13268 7352 13320 7361
rect 15292 7352 15344 7404
rect 14556 7284 14608 7336
rect 3884 7259 3936 7268
rect 3884 7225 3893 7259
rect 3893 7225 3927 7259
rect 3927 7225 3936 7259
rect 3884 7216 3936 7225
rect 7564 7216 7616 7268
rect 9220 7259 9272 7268
rect 9220 7225 9229 7259
rect 9229 7225 9263 7259
rect 9263 7225 9272 7259
rect 9220 7216 9272 7225
rect 10968 7216 11020 7268
rect 5908 7191 5960 7200
rect 5908 7157 5917 7191
rect 5917 7157 5951 7191
rect 5951 7157 5960 7191
rect 5908 7148 5960 7157
rect 7882 7046 7934 7098
rect 7946 7046 7998 7098
rect 8010 7046 8062 7098
rect 8074 7046 8126 7098
rect 14782 7046 14834 7098
rect 14846 7046 14898 7098
rect 14910 7046 14962 7098
rect 14974 7046 15026 7098
rect 7748 6944 7800 6996
rect 10876 6987 10928 6996
rect 10876 6953 10885 6987
rect 10885 6953 10919 6987
rect 10919 6953 10928 6987
rect 10876 6944 10928 6953
rect 17776 6987 17828 6996
rect 17776 6953 17785 6987
rect 17785 6953 17819 6987
rect 17819 6953 17828 6987
rect 17776 6944 17828 6953
rect 3884 6876 3936 6928
rect 5908 6876 5960 6928
rect 7656 6876 7708 6928
rect 10324 6919 10376 6928
rect 10324 6885 10333 6919
rect 10333 6885 10367 6919
rect 10367 6885 10376 6919
rect 10324 6876 10376 6885
rect 4252 6851 4304 6860
rect 4252 6817 4261 6851
rect 4261 6817 4295 6851
rect 4295 6817 4304 6851
rect 4252 6808 4304 6817
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 6184 6851 6236 6860
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 10140 6808 10192 6860
rect 10968 6808 11020 6860
rect 15936 6851 15988 6860
rect 15936 6817 15945 6851
rect 15945 6817 15979 6851
rect 15979 6817 15988 6851
rect 15936 6808 15988 6817
rect 17408 6808 17460 6860
rect 16212 6783 16264 6792
rect 9680 6672 9732 6724
rect 16212 6749 16221 6783
rect 16221 6749 16255 6783
rect 16255 6749 16264 6783
rect 16212 6740 16264 6749
rect 17500 6740 17552 6792
rect 17868 6808 17920 6860
rect 18696 6740 18748 6792
rect 20904 6672 20956 6724
rect 2044 6604 2096 6656
rect 4432 6502 4484 6554
rect 4496 6502 4548 6554
rect 4560 6502 4612 6554
rect 4624 6502 4676 6554
rect 11332 6502 11384 6554
rect 11396 6502 11448 6554
rect 11460 6502 11512 6554
rect 11524 6502 11576 6554
rect 18232 6502 18284 6554
rect 18296 6502 18348 6554
rect 18360 6502 18412 6554
rect 18424 6502 18476 6554
rect 10876 6332 10928 6384
rect 6184 6264 6236 6316
rect 10140 6264 10192 6316
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 16212 6264 16264 6316
rect 3884 6196 3936 6248
rect 5632 6196 5684 6248
rect 6828 6196 6880 6248
rect 15108 6196 15160 6248
rect 17500 6239 17552 6248
rect 17500 6205 17509 6239
rect 17509 6205 17543 6239
rect 17543 6205 17552 6239
rect 17500 6196 17552 6205
rect 17684 6239 17736 6248
rect 17684 6205 17693 6239
rect 17693 6205 17727 6239
rect 17727 6205 17736 6239
rect 17684 6196 17736 6205
rect 17868 6239 17920 6248
rect 17868 6205 17877 6239
rect 17877 6205 17911 6239
rect 17911 6205 17920 6239
rect 17868 6196 17920 6205
rect 18696 6239 18748 6248
rect 18696 6205 18705 6239
rect 18705 6205 18739 6239
rect 18739 6205 18748 6239
rect 18696 6196 18748 6205
rect 18880 6239 18932 6248
rect 18880 6205 18889 6239
rect 18889 6205 18923 6239
rect 18923 6205 18932 6239
rect 18880 6196 18932 6205
rect 2780 6060 2832 6112
rect 5908 6103 5960 6112
rect 5908 6069 5917 6103
rect 5917 6069 5951 6103
rect 5951 6069 5960 6103
rect 5908 6060 5960 6069
rect 10324 6060 10376 6112
rect 15200 6060 15252 6112
rect 18604 6060 18656 6112
rect 7882 5958 7934 6010
rect 7946 5958 7998 6010
rect 8010 5958 8062 6010
rect 8074 5958 8126 6010
rect 14782 5958 14834 6010
rect 14846 5958 14898 6010
rect 14910 5958 14962 6010
rect 14974 5958 15026 6010
rect 6828 5856 6880 5908
rect 15936 5856 15988 5908
rect 18696 5856 18748 5908
rect 20904 5899 20956 5908
rect 20904 5865 20913 5899
rect 20913 5865 20947 5899
rect 20947 5865 20956 5899
rect 20904 5856 20956 5865
rect 4988 5788 5040 5840
rect 13452 5831 13504 5840
rect 13452 5797 13461 5831
rect 13461 5797 13495 5831
rect 13495 5797 13504 5831
rect 13452 5788 13504 5797
rect 14832 5788 14884 5840
rect 15200 5831 15252 5840
rect 15200 5797 15209 5831
rect 15209 5797 15243 5831
rect 15243 5797 15252 5831
rect 15200 5788 15252 5797
rect 17684 5788 17736 5840
rect 2780 5763 2832 5772
rect 2780 5729 2789 5763
rect 2789 5729 2823 5763
rect 2823 5729 2832 5763
rect 2780 5720 2832 5729
rect 8300 5720 8352 5772
rect 12716 5763 12768 5772
rect 12716 5729 12725 5763
rect 12725 5729 12759 5763
rect 12759 5729 12768 5763
rect 12716 5720 12768 5729
rect 14648 5720 14700 5772
rect 15292 5763 15344 5772
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 17316 5720 17368 5772
rect 17868 5720 17920 5772
rect 20812 5720 20864 5772
rect 21088 5763 21140 5772
rect 21088 5729 21097 5763
rect 21097 5729 21131 5763
rect 21131 5729 21140 5763
rect 21088 5720 21140 5729
rect 15200 5652 15252 5704
rect 18880 5652 18932 5704
rect 9680 5584 9732 5636
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 2688 5559 2740 5568
rect 2688 5525 2697 5559
rect 2697 5525 2731 5559
rect 2731 5525 2740 5559
rect 2688 5516 2740 5525
rect 12624 5559 12676 5568
rect 12624 5525 12633 5559
rect 12633 5525 12667 5559
rect 12667 5525 12676 5559
rect 12624 5516 12676 5525
rect 4432 5414 4484 5466
rect 4496 5414 4548 5466
rect 4560 5414 4612 5466
rect 4624 5414 4676 5466
rect 11332 5414 11384 5466
rect 11396 5414 11448 5466
rect 11460 5414 11512 5466
rect 11524 5414 11576 5466
rect 18232 5414 18284 5466
rect 18296 5414 18348 5466
rect 18360 5414 18412 5466
rect 18424 5414 18476 5466
rect 8300 5312 8352 5364
rect 12716 5312 12768 5364
rect 15108 5355 15160 5364
rect 15108 5321 15117 5355
rect 15117 5321 15151 5355
rect 15151 5321 15160 5355
rect 15108 5312 15160 5321
rect 17316 5355 17368 5364
rect 17316 5321 17325 5355
rect 17325 5321 17359 5355
rect 17359 5321 17368 5355
rect 17316 5312 17368 5321
rect 18880 5312 18932 5364
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3240 5176 3292 5185
rect 2044 5108 2096 5160
rect 2688 5108 2740 5160
rect 15200 5244 15252 5296
rect 7012 5108 7064 5160
rect 7564 5151 7616 5160
rect 7564 5117 7573 5151
rect 7573 5117 7607 5151
rect 7607 5117 7616 5151
rect 7564 5108 7616 5117
rect 9680 5108 9732 5160
rect 10232 5151 10284 5160
rect 10232 5117 10241 5151
rect 10241 5117 10275 5151
rect 10275 5117 10284 5151
rect 10232 5108 10284 5117
rect 11060 5108 11112 5160
rect 17776 5176 17828 5228
rect 6276 5040 6328 5092
rect 10968 5083 11020 5092
rect 10968 5049 10977 5083
rect 10977 5049 11011 5083
rect 11011 5049 11020 5083
rect 10968 5040 11020 5049
rect 12624 5040 12676 5092
rect 14832 5108 14884 5160
rect 15292 5151 15344 5160
rect 15292 5117 15301 5151
rect 15301 5117 15335 5151
rect 15335 5117 15344 5151
rect 15292 5108 15344 5117
rect 17500 5108 17552 5160
rect 17684 5015 17736 5024
rect 17684 4981 17693 5015
rect 17693 4981 17727 5015
rect 17727 4981 17736 5015
rect 17684 4972 17736 4981
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 7882 4870 7934 4922
rect 7946 4870 7998 4922
rect 8010 4870 8062 4922
rect 8074 4870 8126 4922
rect 14782 4870 14834 4922
rect 14846 4870 14898 4922
rect 14910 4870 14962 4922
rect 14974 4870 15026 4922
rect 7564 4768 7616 4820
rect 17684 4768 17736 4820
rect 19616 4768 19668 4820
rect 20720 4768 20772 4820
rect 6276 4700 6328 4752
rect 6736 4700 6788 4752
rect 7472 4700 7524 4752
rect 10968 4700 11020 4752
rect 4988 4675 5040 4684
rect 4988 4641 4997 4675
rect 4997 4641 5031 4675
rect 5031 4641 5040 4675
rect 4988 4632 5040 4641
rect 7012 4675 7064 4684
rect 7012 4641 7021 4675
rect 7021 4641 7055 4675
rect 7055 4641 7064 4675
rect 7012 4632 7064 4641
rect 10232 4632 10284 4684
rect 12164 4632 12216 4684
rect 19432 4632 19484 4684
rect 8208 4564 8260 4616
rect 8484 4607 8536 4616
rect 8484 4573 8493 4607
rect 8493 4573 8527 4607
rect 8527 4573 8536 4607
rect 8484 4564 8536 4573
rect 9772 4564 9824 4616
rect 18604 4607 18656 4616
rect 18604 4573 18613 4607
rect 18613 4573 18647 4607
rect 18647 4573 18656 4607
rect 18604 4564 18656 4573
rect 17316 4428 17368 4480
rect 17776 4428 17828 4480
rect 4432 4326 4484 4378
rect 4496 4326 4548 4378
rect 4560 4326 4612 4378
rect 4624 4326 4676 4378
rect 11332 4326 11384 4378
rect 11396 4326 11448 4378
rect 11460 4326 11512 4378
rect 11524 4326 11576 4378
rect 18232 4326 18284 4378
rect 18296 4326 18348 4378
rect 18360 4326 18412 4378
rect 18424 4326 18476 4378
rect 8300 4267 8352 4276
rect 8300 4233 8309 4267
rect 8309 4233 8343 4267
rect 8343 4233 8352 4267
rect 8300 4224 8352 4233
rect 12164 4267 12216 4276
rect 12164 4233 12173 4267
rect 12173 4233 12207 4267
rect 12207 4233 12216 4267
rect 12164 4224 12216 4233
rect 19432 4224 19484 4276
rect 20168 4224 20220 4276
rect 15292 4156 15344 4208
rect 7564 4088 7616 4140
rect 9772 4088 9824 4140
rect 10508 4088 10560 4140
rect 19616 4088 19668 4140
rect 9864 4063 9916 4072
rect 9864 4029 9873 4063
rect 9873 4029 9907 4063
rect 9907 4029 9916 4063
rect 9864 4020 9916 4029
rect 1676 3952 1728 4004
rect 11704 3952 11756 4004
rect 15568 3995 15620 4004
rect 15568 3961 15577 3995
rect 15577 3961 15611 3995
rect 15611 3961 15620 3995
rect 15568 3952 15620 3961
rect 18052 3952 18104 4004
rect 8944 3927 8996 3936
rect 8944 3893 8953 3927
rect 8953 3893 8987 3927
rect 8987 3893 8996 3927
rect 8944 3884 8996 3893
rect 9772 3927 9824 3936
rect 9772 3893 9781 3927
rect 9781 3893 9815 3927
rect 9815 3893 9824 3927
rect 9772 3884 9824 3893
rect 11060 3884 11112 3936
rect 11152 3884 11204 3936
rect 14648 3884 14700 3936
rect 15384 3884 15436 3936
rect 20168 3927 20220 3936
rect 20168 3893 20177 3927
rect 20177 3893 20211 3927
rect 20211 3893 20220 3927
rect 20168 3884 20220 3893
rect 7882 3782 7934 3834
rect 7946 3782 7998 3834
rect 8010 3782 8062 3834
rect 8074 3782 8126 3834
rect 14782 3782 14834 3834
rect 14846 3782 14898 3834
rect 14910 3782 14962 3834
rect 14974 3782 15026 3834
rect 8944 3680 8996 3732
rect 10048 3680 10100 3732
rect 10416 3680 10468 3732
rect 3792 3612 3844 3664
rect 10508 3612 10560 3664
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 6920 3587 6972 3596
rect 6920 3553 6929 3587
rect 6929 3553 6963 3587
rect 6963 3553 6972 3587
rect 6920 3544 6972 3553
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 9036 3476 9088 3528
rect 13176 3612 13228 3664
rect 15568 3680 15620 3732
rect 15384 3612 15436 3664
rect 12624 3544 12676 3596
rect 11980 3476 12032 3528
rect 13912 3544 13964 3596
rect 21088 3587 21140 3596
rect 21088 3553 21097 3587
rect 21097 3553 21131 3587
rect 21131 3553 21140 3587
rect 21088 3544 21140 3553
rect 15568 3476 15620 3528
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 6644 3340 6696 3392
rect 6736 3383 6788 3392
rect 6736 3349 6745 3383
rect 6745 3349 6779 3383
rect 6779 3349 6788 3383
rect 6736 3340 6788 3349
rect 8208 3340 8260 3392
rect 20812 3408 20864 3460
rect 10876 3383 10928 3392
rect 10876 3349 10885 3383
rect 10885 3349 10919 3383
rect 10919 3349 10928 3383
rect 10876 3340 10928 3349
rect 12072 3383 12124 3392
rect 12072 3349 12081 3383
rect 12081 3349 12115 3383
rect 12115 3349 12124 3383
rect 12072 3340 12124 3349
rect 16028 3340 16080 3392
rect 4432 3238 4484 3290
rect 4496 3238 4548 3290
rect 4560 3238 4612 3290
rect 4624 3238 4676 3290
rect 11332 3238 11384 3290
rect 11396 3238 11448 3290
rect 11460 3238 11512 3290
rect 11524 3238 11576 3290
rect 18232 3238 18284 3290
rect 18296 3238 18348 3290
rect 18360 3238 18412 3290
rect 18424 3238 18476 3290
rect 6644 3136 6696 3188
rect 9036 3179 9088 3188
rect 1584 3068 1636 3120
rect 9036 3145 9045 3179
rect 9045 3145 9079 3179
rect 9079 3145 9088 3179
rect 9036 3136 9088 3145
rect 10048 3179 10100 3188
rect 10048 3145 10057 3179
rect 10057 3145 10091 3179
rect 10091 3145 10100 3179
rect 10048 3136 10100 3145
rect 11152 3179 11204 3188
rect 11152 3145 11161 3179
rect 11161 3145 11195 3179
rect 11195 3145 11204 3179
rect 11152 3136 11204 3145
rect 12532 3136 12584 3188
rect 14648 3179 14700 3188
rect 14648 3145 14657 3179
rect 14657 3145 14691 3179
rect 14691 3145 14700 3179
rect 14648 3136 14700 3145
rect 15568 3179 15620 3188
rect 15568 3145 15577 3179
rect 15577 3145 15611 3179
rect 15611 3145 15620 3179
rect 15568 3136 15620 3145
rect 20812 3136 20864 3188
rect 480 2932 532 2984
rect 13912 3068 13964 3120
rect 8484 3043 8536 3052
rect 8484 3009 8493 3043
rect 8493 3009 8527 3043
rect 8527 3009 8536 3043
rect 8484 3000 8536 3009
rect 8760 2932 8812 2984
rect 9036 2932 9088 2984
rect 9680 2932 9732 2984
rect 10876 2932 10928 2984
rect 12624 3000 12676 3052
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 16028 3043 16080 3052
rect 13176 3000 13228 3009
rect 11704 2932 11756 2984
rect 14280 2975 14332 2984
rect 6736 2864 6788 2916
rect 14280 2941 14289 2975
rect 14289 2941 14323 2975
rect 14323 2941 14332 2975
rect 14280 2932 14332 2941
rect 14648 2975 14700 2984
rect 14648 2941 14657 2975
rect 14657 2941 14691 2975
rect 14691 2941 14700 2975
rect 14648 2932 14700 2941
rect 16028 3009 16037 3043
rect 16037 3009 16071 3043
rect 16071 3009 16080 3043
rect 16028 3000 16080 3009
rect 16120 3043 16172 3052
rect 16120 3009 16129 3043
rect 16129 3009 16163 3043
rect 16163 3009 16172 3043
rect 17316 3043 17368 3052
rect 16120 3000 16172 3009
rect 17316 3009 17325 3043
rect 17325 3009 17359 3043
rect 17359 3009 17368 3043
rect 17316 3000 17368 3009
rect 1676 2796 1728 2848
rect 7288 2796 7340 2848
rect 12900 2796 12952 2848
rect 13452 2839 13504 2848
rect 13452 2805 13461 2839
rect 13461 2805 13495 2839
rect 13495 2805 13504 2839
rect 13820 2839 13872 2848
rect 13452 2796 13504 2805
rect 13820 2805 13829 2839
rect 13829 2805 13863 2839
rect 13863 2805 13872 2839
rect 13820 2796 13872 2805
rect 19616 2932 19668 2984
rect 22100 2932 22152 2984
rect 18052 2864 18104 2916
rect 7882 2694 7934 2746
rect 7946 2694 7998 2746
rect 8010 2694 8062 2746
rect 8074 2694 8126 2746
rect 14782 2694 14834 2746
rect 14846 2694 14898 2746
rect 14910 2694 14962 2746
rect 14974 2694 15026 2746
rect 4804 2592 4856 2644
rect 5816 2592 5868 2644
rect 6920 2592 6972 2644
rect 9772 2635 9824 2644
rect 9772 2601 9781 2635
rect 9781 2601 9815 2635
rect 9815 2601 9824 2635
rect 9772 2592 9824 2601
rect 11152 2592 11204 2644
rect 12900 2635 12952 2644
rect 12900 2601 12909 2635
rect 12909 2601 12943 2635
rect 12943 2601 12952 2635
rect 12900 2592 12952 2601
rect 14648 2592 14700 2644
rect 18788 2592 18840 2644
rect 2044 2567 2096 2576
rect 2044 2533 2053 2567
rect 2053 2533 2087 2567
rect 2087 2533 2096 2567
rect 2044 2524 2096 2533
rect 3700 2456 3752 2508
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 6920 2456 6972 2508
rect 8760 2456 8812 2508
rect 10600 2456 10652 2508
rect 10876 2456 10928 2508
rect 12072 2456 12124 2508
rect 13820 2524 13872 2576
rect 14280 2524 14332 2576
rect 17868 2567 17920 2576
rect 17868 2533 17877 2567
rect 17877 2533 17911 2567
rect 17911 2533 17920 2567
rect 17868 2524 17920 2533
rect 20168 2524 20220 2576
rect 13912 2499 13964 2508
rect 13912 2465 13921 2499
rect 13921 2465 13955 2499
rect 13955 2465 13964 2499
rect 13912 2456 13964 2465
rect 15660 2499 15712 2508
rect 15660 2465 15669 2499
rect 15669 2465 15703 2499
rect 15703 2465 15712 2499
rect 15660 2456 15712 2465
rect 17040 2456 17092 2508
rect 18880 2456 18932 2508
rect 13820 2388 13872 2440
rect 16120 2431 16172 2440
rect 16120 2397 16129 2431
rect 16129 2397 16163 2431
rect 16163 2397 16172 2431
rect 16120 2388 16172 2397
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 20720 2363 20772 2372
rect 14556 2252 14608 2304
rect 20720 2329 20729 2363
rect 20729 2329 20763 2363
rect 20763 2329 20772 2363
rect 20720 2320 20772 2329
rect 17500 2252 17552 2304
rect 4432 2150 4484 2202
rect 4496 2150 4548 2202
rect 4560 2150 4612 2202
rect 4624 2150 4676 2202
rect 11332 2150 11384 2202
rect 11396 2150 11448 2202
rect 11460 2150 11512 2202
rect 11524 2150 11576 2202
rect 18232 2150 18284 2202
rect 18296 2150 18348 2202
rect 18360 2150 18412 2202
rect 18424 2150 18476 2202
<< metal2 >>
rect 938 24323 994 25123
rect 2778 24323 2834 25123
rect 4618 24323 4674 25123
rect 5998 24323 6054 25123
rect 7838 24323 7894 25123
rect 9678 24323 9734 25123
rect 11518 24323 11574 25123
rect 12898 24323 12954 25123
rect 14738 24323 14794 25123
rect 16578 24323 16634 25123
rect 17958 24323 18014 25123
rect 19798 24323 19854 25123
rect 21638 24323 21694 25123
rect 952 22574 980 24323
rect 1490 23216 1546 23225
rect 1490 23151 1546 23160
rect 1504 22778 1532 23151
rect 1492 22772 1544 22778
rect 1492 22714 1544 22720
rect 2792 22574 2820 24323
rect 4632 23066 4660 24323
rect 4632 23038 4844 23066
rect 4406 22876 4702 22896
rect 4462 22874 4486 22876
rect 4542 22874 4566 22876
rect 4622 22874 4646 22876
rect 4484 22822 4486 22874
rect 4548 22822 4560 22874
rect 4622 22822 4624 22874
rect 4462 22820 4486 22822
rect 4542 22820 4566 22822
rect 4622 22820 4646 22822
rect 4406 22800 4702 22820
rect 4816 22574 4844 23038
rect 5448 22704 5500 22710
rect 5448 22646 5500 22652
rect 940 22568 992 22574
rect 940 22510 992 22516
rect 2780 22568 2832 22574
rect 2780 22510 2832 22516
rect 4712 22568 4764 22574
rect 4712 22510 4764 22516
rect 4804 22568 4856 22574
rect 4804 22510 4856 22516
rect 1584 22500 1636 22506
rect 1584 22442 1636 22448
rect 1596 21690 1624 22442
rect 2044 22432 2096 22438
rect 2044 22374 2096 22380
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1398 20496 1454 20505
rect 1398 20431 1454 20440
rect 1412 20398 1440 20431
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1492 20256 1544 20262
rect 1492 20198 1544 20204
rect 1398 17776 1454 17785
rect 1398 17711 1400 17720
rect 1452 17711 1454 17720
rect 1400 17682 1452 17688
rect 1398 15736 1454 15745
rect 1398 15671 1454 15680
rect 1412 15570 1440 15671
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1504 13138 1532 20198
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 1596 13530 1624 17478
rect 1952 16040 2004 16046
rect 1952 15982 2004 15988
rect 1964 15502 1992 15982
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1412 13110 1532 13138
rect 1412 9110 1440 13110
rect 1490 13016 1546 13025
rect 1490 12951 1492 12960
rect 1544 12951 1546 12960
rect 1492 12922 1544 12928
rect 1872 11354 1900 15302
rect 1964 15162 1992 15438
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 2056 15026 2084 22374
rect 4724 22030 4752 22510
rect 4896 22432 4948 22438
rect 4896 22374 4948 22380
rect 4712 22024 4764 22030
rect 4712 21966 4764 21972
rect 4160 21888 4212 21894
rect 4724 21876 4752 21966
rect 4724 21848 4844 21876
rect 4160 21830 4212 21836
rect 4172 21554 4200 21830
rect 4406 21788 4702 21808
rect 4462 21786 4486 21788
rect 4542 21786 4566 21788
rect 4622 21786 4646 21788
rect 4484 21734 4486 21786
rect 4548 21734 4560 21786
rect 4622 21734 4624 21786
rect 4462 21732 4486 21734
rect 4542 21732 4566 21734
rect 4622 21732 4646 21734
rect 4406 21712 4702 21732
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 2504 21480 2556 21486
rect 2504 21422 2556 21428
rect 2516 20466 2544 21422
rect 4406 20700 4702 20720
rect 4462 20698 4486 20700
rect 4542 20698 4566 20700
rect 4622 20698 4646 20700
rect 4484 20646 4486 20698
rect 4548 20646 4560 20698
rect 4622 20646 4624 20698
rect 4462 20644 4486 20646
rect 4542 20644 4566 20646
rect 4622 20644 4646 20646
rect 4406 20624 4702 20644
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 2516 18290 2544 20402
rect 3332 20324 3384 20330
rect 3332 20266 3384 20272
rect 3344 20058 3372 20266
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 4172 20058 4200 20198
rect 3332 20052 3384 20058
rect 3332 19994 3384 20000
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4816 19922 4844 21848
rect 4908 21418 4936 22374
rect 4988 22092 5040 22098
rect 4988 22034 5040 22040
rect 5080 22092 5132 22098
rect 5080 22034 5132 22040
rect 4896 21412 4948 21418
rect 4896 21354 4948 21360
rect 5000 21146 5028 22034
rect 4988 21140 5040 21146
rect 4988 21082 5040 21088
rect 5092 20874 5120 22034
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 5080 20868 5132 20874
rect 5080 20810 5132 20816
rect 4988 20800 5040 20806
rect 4988 20742 5040 20748
rect 4804 19916 4856 19922
rect 4804 19858 4856 19864
rect 4406 19612 4702 19632
rect 4462 19610 4486 19612
rect 4542 19610 4566 19612
rect 4622 19610 4646 19612
rect 4484 19558 4486 19610
rect 4548 19558 4560 19610
rect 4622 19558 4624 19610
rect 4462 19556 4486 19558
rect 4542 19556 4566 19558
rect 4622 19556 4646 19558
rect 4406 19536 4702 19556
rect 4406 18524 4702 18544
rect 4462 18522 4486 18524
rect 4542 18522 4566 18524
rect 4622 18522 4646 18524
rect 4484 18470 4486 18522
rect 4548 18470 4560 18522
rect 4622 18470 4624 18522
rect 4462 18468 4486 18470
rect 4542 18468 4566 18470
rect 4622 18468 4646 18470
rect 4406 18448 4702 18468
rect 4816 18442 4844 19858
rect 5000 19854 5028 20742
rect 4988 19848 5040 19854
rect 4988 19790 5040 19796
rect 4816 18414 4936 18442
rect 2504 18284 2556 18290
rect 2504 18226 2556 18232
rect 3240 18148 3292 18154
rect 3240 18090 3292 18096
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 3252 17882 3280 18090
rect 4264 17882 4292 18090
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 3240 17876 3292 17882
rect 3240 17818 3292 17824
rect 4252 17876 4304 17882
rect 4252 17818 4304 17824
rect 4816 17746 4844 18022
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4908 17678 4936 18414
rect 5000 17746 5028 19790
rect 5092 19786 5120 20810
rect 5276 20806 5304 21830
rect 5264 20800 5316 20806
rect 5264 20742 5316 20748
rect 5264 20392 5316 20398
rect 5264 20334 5316 20340
rect 5172 20256 5224 20262
rect 5172 20198 5224 20204
rect 5184 19922 5212 20198
rect 5172 19916 5224 19922
rect 5172 19858 5224 19864
rect 5080 19780 5132 19786
rect 5080 19722 5132 19728
rect 5092 18306 5120 19722
rect 5184 19310 5212 19858
rect 5276 19786 5304 20334
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5368 19990 5396 20198
rect 5356 19984 5408 19990
rect 5356 19926 5408 19932
rect 5264 19780 5316 19786
rect 5264 19722 5316 19728
rect 5276 19514 5304 19722
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5368 18766 5396 19926
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 5092 18278 5212 18306
rect 5080 18148 5132 18154
rect 5080 18090 5132 18096
rect 5092 17746 5120 18090
rect 4988 17740 5040 17746
rect 4988 17682 5040 17688
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4406 17436 4702 17456
rect 4462 17434 4486 17436
rect 4542 17434 4566 17436
rect 4622 17434 4646 17436
rect 4484 17382 4486 17434
rect 4548 17382 4560 17434
rect 4622 17382 4624 17434
rect 4462 17380 4486 17382
rect 4542 17380 4566 17382
rect 4622 17380 4646 17382
rect 4406 17360 4702 17380
rect 4406 16348 4702 16368
rect 4462 16346 4486 16348
rect 4542 16346 4566 16348
rect 4622 16346 4646 16348
rect 4484 16294 4486 16346
rect 4548 16294 4560 16346
rect 4622 16294 4624 16346
rect 4462 16292 4486 16294
rect 4542 16292 4566 16294
rect 4622 16292 4646 16294
rect 4406 16272 4702 16292
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 2700 15434 2728 15914
rect 2884 15502 2912 15982
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2688 15428 2740 15434
rect 2688 15370 2740 15376
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1964 14074 1992 14758
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2148 13326 2176 14962
rect 2136 13320 2188 13326
rect 2188 13268 2268 13274
rect 2136 13262 2268 13268
rect 2148 13246 2268 13262
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2148 12782 2176 13126
rect 2136 12776 2188 12782
rect 2136 12718 2188 12724
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 2240 11150 2268 13246
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 1584 11008 1636 11014
rect 1584 10950 1636 10956
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 1504 10305 1532 10406
rect 1490 10296 1546 10305
rect 1490 10231 1546 10240
rect 1596 10130 1624 10950
rect 2044 10532 2096 10538
rect 2044 10474 2096 10480
rect 1584 10124 1636 10130
rect 1584 10066 1636 10072
rect 1596 9518 1624 10066
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1400 9104 1452 9110
rect 1400 9046 1452 9052
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 8265 1440 8366
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 2056 6662 2084 10474
rect 2240 10418 2268 11086
rect 2700 10606 2728 15370
rect 2884 14958 2912 15438
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2884 14006 2912 14894
rect 3252 14822 3280 15506
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 4264 15094 4292 15302
rect 4406 15260 4702 15280
rect 4462 15258 4486 15260
rect 4542 15258 4566 15260
rect 4622 15258 4646 15260
rect 4484 15206 4486 15258
rect 4548 15206 4560 15258
rect 4622 15206 4624 15258
rect 4462 15204 4486 15206
rect 4542 15204 4566 15206
rect 4622 15204 4646 15206
rect 4406 15184 4702 15204
rect 4252 15088 4304 15094
rect 4252 15030 4304 15036
rect 4908 14958 4936 17614
rect 5000 15434 5028 17682
rect 5184 17660 5212 18278
rect 5264 17672 5316 17678
rect 5184 17632 5264 17660
rect 5264 17614 5316 17620
rect 4988 15428 5040 15434
rect 4988 15370 5040 15376
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4816 14550 4844 14758
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4406 14172 4702 14192
rect 4462 14170 4486 14172
rect 4542 14170 4566 14172
rect 4622 14170 4646 14172
rect 4484 14118 4486 14170
rect 4548 14118 4560 14170
rect 4622 14118 4624 14170
rect 4462 14116 4486 14118
rect 4542 14116 4566 14118
rect 4622 14116 4646 14118
rect 4406 14096 4702 14116
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 3332 13796 3384 13802
rect 3332 13738 3384 13744
rect 3344 12986 3372 13738
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 4406 13084 4702 13104
rect 4462 13082 4486 13084
rect 4542 13082 4566 13084
rect 4622 13082 4646 13084
rect 4484 13030 4486 13082
rect 4548 13030 4560 13082
rect 4622 13030 4624 13082
rect 4462 13028 4486 13030
rect 4542 13028 4566 13030
rect 4622 13028 4646 13030
rect 4406 13008 4702 13028
rect 4908 12986 4936 13330
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 2792 11694 2820 12718
rect 3240 12708 3292 12714
rect 3240 12650 3292 12656
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 2976 11898 3004 12242
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2976 11354 3004 11834
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2872 10532 2924 10538
rect 2872 10474 2924 10480
rect 2240 10390 2452 10418
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2240 9722 2268 10202
rect 2228 9716 2280 9722
rect 2228 9658 2280 9664
rect 2240 9178 2268 9658
rect 2424 9450 2452 10390
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2792 9654 2820 9930
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2884 9518 2912 10474
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2412 9444 2464 9450
rect 2412 9386 2464 9392
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2148 7954 2176 8570
rect 2424 8362 2452 9386
rect 2884 9058 2912 9454
rect 2700 9030 2912 9058
rect 2504 8900 2556 8906
rect 2504 8842 2556 8848
rect 2516 8430 2544 8842
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2412 8356 2464 8362
rect 2412 8298 2464 8304
rect 2700 7954 2728 9030
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2792 5778 2820 6054
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 1492 5568 1544 5574
rect 1490 5536 1492 5545
rect 2688 5568 2740 5574
rect 1544 5536 1546 5545
rect 2688 5510 2740 5516
rect 1490 5471 1546 5480
rect 2700 5166 2728 5510
rect 3252 5234 3280 12650
rect 3344 12374 3372 12718
rect 4988 12708 5040 12714
rect 4988 12650 5040 12656
rect 5000 12434 5028 12650
rect 4908 12406 5028 12434
rect 5184 12434 5212 12718
rect 5184 12406 5304 12434
rect 3332 12368 3384 12374
rect 3332 12310 3384 12316
rect 4406 11996 4702 12016
rect 4462 11994 4486 11996
rect 4542 11994 4566 11996
rect 4622 11994 4646 11996
rect 4484 11942 4486 11994
rect 4548 11942 4560 11994
rect 4622 11942 4624 11994
rect 4462 11940 4486 11942
rect 4542 11940 4566 11942
rect 4622 11940 4646 11942
rect 4406 11920 4702 11940
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3528 11150 3556 11630
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 4080 11150 4108 11562
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3896 8498 3924 8774
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3804 7750 3832 8298
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 1676 4004 1728 4010
rect 1676 3946 1728 3952
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 480 2984 532 2990
rect 480 2926 532 2932
rect 492 800 520 2926
rect 1412 2825 1440 3538
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1596 3126 1624 3334
rect 1584 3120 1636 3126
rect 1584 3062 1636 3068
rect 1688 2854 1716 3946
rect 1676 2848 1728 2854
rect 1398 2816 1454 2825
rect 1676 2790 1728 2796
rect 1398 2751 1454 2760
rect 2056 2582 2084 5102
rect 3804 3670 3832 7686
rect 4080 7546 4108 11086
rect 4264 10810 4292 11222
rect 4406 10908 4702 10928
rect 4462 10906 4486 10908
rect 4542 10906 4566 10908
rect 4622 10906 4646 10908
rect 4484 10854 4486 10906
rect 4548 10854 4560 10906
rect 4622 10854 4624 10906
rect 4462 10852 4486 10854
rect 4542 10852 4566 10854
rect 4622 10852 4646 10854
rect 4406 10832 4702 10852
rect 4908 10810 4936 12406
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4406 9820 4702 9840
rect 4462 9818 4486 9820
rect 4542 9818 4566 9820
rect 4622 9818 4646 9820
rect 4484 9766 4486 9818
rect 4548 9766 4560 9818
rect 4622 9766 4624 9818
rect 4462 9764 4486 9766
rect 4542 9764 4566 9766
rect 4622 9764 4646 9766
rect 4406 9744 4702 9764
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4908 9330 4936 10746
rect 5000 9518 5028 11494
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 4406 8732 4702 8752
rect 4462 8730 4486 8732
rect 4542 8730 4566 8732
rect 4622 8730 4646 8732
rect 4484 8678 4486 8730
rect 4548 8678 4560 8730
rect 4622 8678 4624 8730
rect 4462 8676 4486 8678
rect 4542 8676 4566 8678
rect 4622 8676 4646 8678
rect 4406 8656 4702 8676
rect 4406 7644 4702 7664
rect 4462 7642 4486 7644
rect 4542 7642 4566 7644
rect 4622 7642 4646 7644
rect 4484 7590 4486 7642
rect 4548 7590 4560 7642
rect 4622 7590 4624 7642
rect 4462 7588 4486 7590
rect 4542 7588 4566 7590
rect 4622 7588 4646 7590
rect 4406 7568 4702 7588
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 3896 6934 3924 7210
rect 3884 6928 3936 6934
rect 3884 6870 3936 6876
rect 3896 6254 3924 6870
rect 4264 6866 4292 7346
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4406 6556 4702 6576
rect 4462 6554 4486 6556
rect 4542 6554 4566 6556
rect 4622 6554 4646 6556
rect 4484 6502 4486 6554
rect 4548 6502 4560 6554
rect 4622 6502 4624 6554
rect 4462 6500 4486 6502
rect 4542 6500 4566 6502
rect 4622 6500 4646 6502
rect 4406 6480 4702 6500
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 4406 5468 4702 5488
rect 4462 5466 4486 5468
rect 4542 5466 4566 5468
rect 4622 5466 4646 5468
rect 4484 5414 4486 5466
rect 4548 5414 4560 5466
rect 4622 5414 4624 5466
rect 4462 5412 4486 5414
rect 4542 5412 4566 5414
rect 4622 5412 4646 5414
rect 4406 5392 4702 5412
rect 4406 4380 4702 4400
rect 4462 4378 4486 4380
rect 4542 4378 4566 4380
rect 4622 4378 4646 4380
rect 4484 4326 4486 4378
rect 4548 4326 4560 4378
rect 4622 4326 4624 4378
rect 4462 4324 4486 4326
rect 4542 4324 4566 4326
rect 4622 4324 4646 4326
rect 4406 4304 4702 4324
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 4406 3292 4702 3312
rect 4462 3290 4486 3292
rect 4542 3290 4566 3292
rect 4622 3290 4646 3292
rect 4484 3238 4486 3290
rect 4548 3238 4560 3290
rect 4622 3238 4624 3290
rect 4462 3236 4486 3238
rect 4542 3236 4566 3238
rect 4622 3236 4646 3238
rect 4406 3216 4702 3236
rect 4816 2650 4844 9318
rect 4908 9302 5028 9330
rect 5000 9042 5028 9302
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 5000 8634 5028 8978
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5092 7410 5120 12038
rect 5184 10062 5212 12242
rect 5276 11626 5304 12406
rect 5264 11620 5316 11626
rect 5264 11562 5316 11568
rect 5276 10606 5304 11562
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5356 10260 5408 10266
rect 5460 10248 5488 22646
rect 6012 22574 6040 24323
rect 7852 22574 7880 24323
rect 9692 22574 9720 24323
rect 11532 23066 11560 24323
rect 11532 23038 11744 23066
rect 11306 22876 11602 22896
rect 11362 22874 11386 22876
rect 11442 22874 11466 22876
rect 11522 22874 11546 22876
rect 11384 22822 11386 22874
rect 11448 22822 11460 22874
rect 11522 22822 11524 22874
rect 11362 22820 11386 22822
rect 11442 22820 11466 22822
rect 11522 22820 11546 22822
rect 11306 22800 11602 22820
rect 11060 22704 11112 22710
rect 11060 22646 11112 22652
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 7840 22568 7892 22574
rect 7840 22510 7892 22516
rect 9680 22568 9732 22574
rect 9680 22510 9732 22516
rect 6184 22432 6236 22438
rect 6184 22374 6236 22380
rect 7012 22432 7064 22438
rect 7012 22374 7064 22380
rect 10600 22432 10652 22438
rect 10600 22374 10652 22380
rect 5540 22092 5592 22098
rect 5540 22034 5592 22040
rect 5552 21350 5580 22034
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 5552 21010 5580 21286
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 5552 20398 5580 20946
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 6000 20392 6052 20398
rect 6000 20334 6052 20340
rect 6012 19990 6040 20334
rect 6000 19984 6052 19990
rect 6000 19926 6052 19932
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 5552 18970 5580 19246
rect 5632 19236 5684 19242
rect 5632 19178 5684 19184
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5644 18834 5672 19178
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5724 18692 5776 18698
rect 5724 18634 5776 18640
rect 5736 18222 5764 18634
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5632 18148 5684 18154
rect 5632 18090 5684 18096
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5552 17134 5580 17682
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5552 14618 5580 17070
rect 5644 16998 5672 18090
rect 5828 17338 5856 18906
rect 5920 18766 5948 19246
rect 5908 18760 5960 18766
rect 5908 18702 5960 18708
rect 6092 17808 6144 17814
rect 6092 17750 6144 17756
rect 5816 17332 5868 17338
rect 5816 17274 5868 17280
rect 5908 17264 5960 17270
rect 5908 17206 5960 17212
rect 5724 17128 5776 17134
rect 5724 17070 5776 17076
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5736 15638 5764 17070
rect 5816 17060 5868 17066
rect 5816 17002 5868 17008
rect 5828 16658 5856 17002
rect 5920 16658 5948 17206
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 5724 15632 5776 15638
rect 5724 15574 5776 15580
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 5828 14278 5856 16594
rect 6104 16590 6132 17750
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5552 12442 5580 13806
rect 6104 13462 6132 14554
rect 6092 13456 6144 13462
rect 6092 13398 6144 13404
rect 5540 12436 5592 12442
rect 6104 12434 6132 13398
rect 6196 13326 6224 22374
rect 6644 19236 6696 19242
rect 6644 19178 6696 19184
rect 6656 18970 6684 19178
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 6656 18426 6684 18906
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 6656 17066 6684 17682
rect 6748 17134 6776 18770
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6840 17746 6868 18158
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6736 17128 6788 17134
rect 6736 17070 6788 17076
rect 6644 17060 6696 17066
rect 6644 17002 6696 17008
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6564 16658 6592 16934
rect 6656 16794 6684 17002
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6288 15502 6316 15846
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6380 14550 6408 15302
rect 6840 15162 6868 16050
rect 6932 16046 6960 16662
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6932 15570 6960 15982
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6368 14544 6420 14550
rect 6368 14486 6420 14492
rect 6840 14482 6868 14894
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6840 14346 6868 14418
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6656 14006 6684 14214
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6748 13870 6776 14214
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6840 13394 6868 14282
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6932 13462 6960 13806
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6840 12918 6868 13330
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6840 12434 6868 12854
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 5540 12378 5592 12384
rect 5920 12406 6132 12434
rect 6748 12406 6868 12434
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5644 11694 5672 12038
rect 5736 11762 5764 12242
rect 5920 12238 5948 12406
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5644 11286 5672 11630
rect 5632 11280 5684 11286
rect 5632 11222 5684 11228
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5408 10220 5488 10248
rect 5356 10202 5408 10208
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5184 9450 5212 9998
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 5460 8956 5488 9386
rect 5552 9110 5580 11154
rect 5644 10674 5672 11222
rect 5920 11218 5948 12174
rect 6748 12170 6776 12406
rect 6932 12306 6960 12650
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6840 11762 6868 12174
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 6012 11150 6040 11698
rect 6840 11218 6868 11698
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5920 10198 5948 10950
rect 5908 10192 5960 10198
rect 5908 10134 5960 10140
rect 6012 9110 6040 11086
rect 7024 10266 7052 22374
rect 7856 22332 8152 22352
rect 7912 22330 7936 22332
rect 7992 22330 8016 22332
rect 8072 22330 8096 22332
rect 7934 22278 7936 22330
rect 7998 22278 8010 22330
rect 8072 22278 8074 22330
rect 7912 22276 7936 22278
rect 7992 22276 8016 22278
rect 8072 22276 8096 22278
rect 7856 22256 8152 22276
rect 10324 22092 10376 22098
rect 10324 22034 10376 22040
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 7760 21418 7788 21830
rect 8208 21616 8260 21622
rect 8208 21558 8260 21564
rect 7196 21412 7248 21418
rect 7196 21354 7248 21360
rect 7748 21412 7800 21418
rect 7748 21354 7800 21360
rect 7208 21146 7236 21354
rect 7856 21244 8152 21264
rect 7912 21242 7936 21244
rect 7992 21242 8016 21244
rect 8072 21242 8096 21244
rect 7934 21190 7936 21242
rect 7998 21190 8010 21242
rect 8072 21190 8074 21242
rect 7912 21188 7936 21190
rect 7992 21188 8016 21190
rect 8072 21188 8096 21190
rect 7856 21168 8152 21188
rect 7196 21140 7248 21146
rect 7196 21082 7248 21088
rect 8220 21078 8248 21558
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 9140 21350 9168 21490
rect 10060 21418 10088 21830
rect 10048 21412 10100 21418
rect 10048 21354 10100 21360
rect 9128 21344 9180 21350
rect 9128 21286 9180 21292
rect 7472 21072 7524 21078
rect 7472 21014 7524 21020
rect 7656 21072 7708 21078
rect 7656 21014 7708 21020
rect 8208 21072 8260 21078
rect 8208 21014 8260 21020
rect 7380 21004 7432 21010
rect 7380 20946 7432 20952
rect 7392 20602 7420 20946
rect 7380 20596 7432 20602
rect 7380 20538 7432 20544
rect 7484 20058 7512 21014
rect 7668 20482 7696 21014
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 7576 20454 7696 20482
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7300 18902 7328 19110
rect 7288 18896 7340 18902
rect 7288 18838 7340 18844
rect 7392 18834 7420 19246
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7392 18630 7420 18770
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7104 17808 7156 17814
rect 7104 17750 7156 17756
rect 7116 17202 7144 17750
rect 7484 17678 7512 19790
rect 7576 19394 7604 20454
rect 7656 20392 7708 20398
rect 7656 20334 7708 20340
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 7668 19854 7696 20334
rect 7760 19922 7788 20334
rect 7856 20156 8152 20176
rect 7912 20154 7936 20156
rect 7992 20154 8016 20156
rect 8072 20154 8096 20156
rect 7934 20102 7936 20154
rect 7998 20102 8010 20154
rect 8072 20102 8074 20154
rect 7912 20100 7936 20102
rect 7992 20100 8016 20102
rect 8072 20100 8096 20102
rect 7856 20080 8152 20100
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7656 19848 7708 19854
rect 7656 19790 7708 19796
rect 7576 19366 7696 19394
rect 7668 19242 7696 19366
rect 7656 19236 7708 19242
rect 7656 19178 7708 19184
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7484 17338 7512 17614
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 7380 17264 7432 17270
rect 7380 17206 7432 17212
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 7208 16046 7236 17070
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7300 15706 7328 15982
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7196 15632 7248 15638
rect 7196 15574 7248 15580
rect 7208 15162 7236 15574
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7208 13870 7236 14350
rect 7300 13938 7328 15506
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7116 11218 7144 13466
rect 7208 12782 7236 13806
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7194 12608 7250 12617
rect 7194 12543 7250 12552
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 5724 8968 5776 8974
rect 5460 8928 5724 8956
rect 5724 8910 5776 8916
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5644 6254 5672 6802
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 4988 5840 5040 5846
rect 4988 5782 5040 5788
rect 5000 4690 5028 5782
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 5828 2650 5856 9046
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5920 6934 5948 7142
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5920 6118 5948 6870
rect 6196 6866 6224 9862
rect 7208 9586 7236 12543
rect 7300 11626 7328 13874
rect 7392 13530 7420 17206
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7484 14958 7512 15438
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7484 14278 7512 14894
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7484 13870 7512 14214
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7392 11898 7420 12718
rect 7484 12434 7512 13806
rect 7576 12617 7604 14826
rect 7668 13938 7696 19178
rect 7760 19174 7788 19858
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7760 17746 7788 19110
rect 7856 19068 8152 19088
rect 7912 19066 7936 19068
rect 7992 19066 8016 19068
rect 8072 19066 8096 19068
rect 7934 19014 7936 19066
rect 7998 19014 8010 19066
rect 8072 19014 8074 19066
rect 7912 19012 7936 19014
rect 7992 19012 8016 19014
rect 8072 19012 8096 19014
rect 7856 18992 8152 19012
rect 8220 18766 8248 19994
rect 8496 19310 8524 20946
rect 9140 20466 9168 21286
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 8484 19304 8536 19310
rect 8484 19246 8536 19252
rect 8944 19304 8996 19310
rect 8944 19246 8996 19252
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8496 18698 8524 19246
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8852 19236 8904 19242
rect 8852 19178 8904 19184
rect 8772 18834 8800 19178
rect 8864 18970 8892 19178
rect 8852 18964 8904 18970
rect 8852 18906 8904 18912
rect 8956 18902 8984 19246
rect 8944 18896 8996 18902
rect 8944 18838 8996 18844
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8484 18692 8536 18698
rect 8484 18634 8536 18640
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8588 18290 8616 18566
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 7856 17980 8152 18000
rect 7912 17978 7936 17980
rect 7992 17978 8016 17980
rect 8072 17978 8096 17980
rect 7934 17926 7936 17978
rect 7998 17926 8010 17978
rect 8072 17926 8074 17978
rect 7912 17924 7936 17926
rect 7992 17924 8016 17926
rect 8072 17924 8096 17926
rect 7856 17904 8152 17924
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 7856 16892 8152 16912
rect 7912 16890 7936 16892
rect 7992 16890 8016 16892
rect 8072 16890 8096 16892
rect 7934 16838 7936 16890
rect 7998 16838 8010 16890
rect 8072 16838 8074 16890
rect 7912 16836 7936 16838
rect 7992 16836 8016 16838
rect 8072 16836 8096 16838
rect 7856 16816 8152 16836
rect 8312 16726 8340 17478
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8312 15978 8340 16662
rect 8300 15972 8352 15978
rect 8300 15914 8352 15920
rect 7856 15804 8152 15824
rect 7912 15802 7936 15804
rect 7992 15802 8016 15804
rect 8072 15802 8096 15804
rect 7934 15750 7936 15802
rect 7998 15750 8010 15802
rect 8072 15750 8074 15802
rect 7912 15748 7936 15750
rect 7992 15748 8016 15750
rect 8072 15748 8096 15750
rect 7856 15728 8152 15748
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8312 15026 8340 15506
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 7856 14716 8152 14736
rect 7912 14714 7936 14716
rect 7992 14714 8016 14716
rect 8072 14714 8096 14716
rect 7934 14662 7936 14714
rect 7998 14662 8010 14714
rect 8072 14662 8074 14714
rect 7912 14660 7936 14662
rect 7992 14660 8016 14662
rect 8072 14660 8096 14662
rect 7856 14640 8152 14660
rect 8300 14544 8352 14550
rect 8300 14486 8352 14492
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7668 13734 7696 13874
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7668 12714 7696 13670
rect 7856 13628 8152 13648
rect 7912 13626 7936 13628
rect 7992 13626 8016 13628
rect 8072 13626 8096 13628
rect 7934 13574 7936 13626
rect 7998 13574 8010 13626
rect 8072 13574 8074 13626
rect 7912 13572 7936 13574
rect 7992 13572 8016 13574
rect 8072 13572 8096 13574
rect 7856 13552 8152 13572
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 8220 12646 8248 13330
rect 8208 12640 8260 12646
rect 7562 12608 7618 12617
rect 8208 12582 8260 12588
rect 7562 12543 7618 12552
rect 7856 12540 8152 12560
rect 7912 12538 7936 12540
rect 7992 12538 8016 12540
rect 8072 12538 8096 12540
rect 7934 12486 7936 12538
rect 7998 12486 8010 12538
rect 8072 12486 8074 12538
rect 7912 12484 7936 12486
rect 7992 12484 8016 12486
rect 8072 12484 8096 12486
rect 7856 12464 8152 12484
rect 7484 12406 7604 12434
rect 7576 12306 7604 12406
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6288 8566 6316 8774
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6196 6322 6224 6802
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 6840 5914 6868 6190
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6276 5092 6328 5098
rect 6276 5034 6328 5040
rect 6288 4758 6316 5034
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6736 4752 6788 4758
rect 6736 4694 6788 4700
rect 6748 3398 6776 4694
rect 6932 3602 6960 8978
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 7024 4690 7052 5102
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6656 3194 6684 3334
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6748 2922 6776 3334
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6932 2650 6960 3538
rect 7300 2854 7328 11018
rect 7392 10266 7420 11086
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7484 4758 7512 12106
rect 7576 10810 7604 12242
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7668 11762 7696 12038
rect 8220 11898 8248 12174
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7668 11218 7696 11698
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7668 10742 7696 11154
rect 7656 10736 7708 10742
rect 7656 10678 7708 10684
rect 7760 10606 7788 11562
rect 7856 11452 8152 11472
rect 7912 11450 7936 11452
rect 7992 11450 8016 11452
rect 8072 11450 8096 11452
rect 7934 11398 7936 11450
rect 7998 11398 8010 11450
rect 8072 11398 8074 11450
rect 7912 11396 7936 11398
rect 7992 11396 8016 11398
rect 8072 11396 8096 11398
rect 7856 11376 8152 11396
rect 8220 11218 8248 11834
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7576 8974 7604 9454
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7576 8430 7604 8910
rect 7668 8906 7696 10406
rect 7856 10364 8152 10384
rect 7912 10362 7936 10364
rect 7992 10362 8016 10364
rect 8072 10362 8096 10364
rect 7934 10310 7936 10362
rect 7998 10310 8010 10362
rect 8072 10310 8074 10362
rect 7912 10308 7936 10310
rect 7992 10308 8016 10310
rect 8072 10308 8096 10310
rect 7856 10288 8152 10308
rect 8220 10130 8248 11154
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 7856 9276 8152 9296
rect 7912 9274 7936 9276
rect 7992 9274 8016 9276
rect 8072 9274 8096 9276
rect 7934 9222 7936 9274
rect 7998 9222 8010 9274
rect 8072 9222 8074 9274
rect 7912 9220 7936 9222
rect 7992 9220 8016 9222
rect 8072 9220 8096 9222
rect 7856 9200 8152 9220
rect 7656 8900 7708 8906
rect 7656 8842 7708 8848
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7576 7274 7604 8366
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7668 6934 7696 8842
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7760 7954 7788 8774
rect 7856 8188 8152 8208
rect 7912 8186 7936 8188
rect 7992 8186 8016 8188
rect 8072 8186 8096 8188
rect 7934 8134 7936 8186
rect 7998 8134 8010 8186
rect 8072 8134 8074 8186
rect 7912 8132 7936 8134
rect 7992 8132 8016 8134
rect 8072 8132 8096 8134
rect 7856 8112 8152 8132
rect 8312 8022 8340 14486
rect 8404 13530 8432 17614
rect 8496 17610 8524 18022
rect 8588 17746 8616 18226
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8496 15910 8524 17070
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8588 16046 8616 16934
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 8496 15706 8524 15846
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8680 14074 8708 18770
rect 8772 18086 8800 18770
rect 9036 18692 9088 18698
rect 9036 18634 9088 18640
rect 8852 18148 8904 18154
rect 8852 18090 8904 18096
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8864 17542 8892 18090
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 8864 16776 8892 17478
rect 8772 16748 8892 16776
rect 8772 14414 8800 16748
rect 8852 16652 8904 16658
rect 8852 16594 8904 16600
rect 8864 16046 8892 16594
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 8956 15638 8984 17682
rect 9048 16114 9076 18634
rect 9140 17746 9168 20402
rect 10336 19922 10364 22034
rect 10416 20324 10468 20330
rect 10416 20266 10468 20272
rect 10428 20058 10456 20266
rect 10416 20052 10468 20058
rect 10416 19994 10468 20000
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9508 18290 9536 19110
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 10336 18222 10364 19858
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 8944 15632 8996 15638
rect 8944 15574 8996 15580
rect 9140 15502 9168 17682
rect 9692 16250 9720 18158
rect 10232 18148 10284 18154
rect 10232 18090 10284 18096
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9784 17814 9812 18022
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10152 17134 10180 17478
rect 10244 17338 10272 18090
rect 10508 18080 10560 18086
rect 10508 18022 10560 18028
rect 10520 17814 10548 18022
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9140 14550 9168 15438
rect 9692 15434 9720 16186
rect 9864 16040 9916 16046
rect 10244 15994 10272 17274
rect 10612 17252 10640 22374
rect 10876 22160 10928 22166
rect 10876 22102 10928 22108
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10704 21554 10732 21830
rect 10888 21690 10916 22102
rect 10876 21684 10928 21690
rect 10876 21626 10928 21632
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 9864 15982 9916 15988
rect 9876 15570 9904 15982
rect 10152 15966 10272 15994
rect 10520 17224 10640 17252
rect 9864 15564 9916 15570
rect 9864 15506 9916 15512
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9876 15162 9904 15506
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9128 14544 9180 14550
rect 9128 14486 9180 14492
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8404 12782 8432 13466
rect 8588 13394 8616 13806
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8680 13190 8708 14010
rect 9876 13954 9904 15098
rect 10152 14006 10180 15966
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 10244 15638 10272 15846
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10244 14074 10272 14962
rect 10428 14958 10456 15302
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10324 14340 10376 14346
rect 10324 14282 10376 14288
rect 10336 14074 10364 14282
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9784 13926 9904 13954
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8956 11762 8984 12718
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9232 11898 9260 12582
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8484 10532 8536 10538
rect 8484 10474 8536 10480
rect 8496 9518 8524 10474
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8588 10130 8616 10406
rect 9232 10198 9260 11834
rect 9324 11694 9352 13126
rect 9416 12918 9444 13738
rect 9692 13394 9720 13874
rect 9784 13870 9812 13926
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9220 10192 9272 10198
rect 9220 10134 9272 10140
rect 9416 10130 9444 12854
rect 9508 10606 9536 13330
rect 9692 12782 9720 13330
rect 9784 12986 9812 13806
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9968 12782 9996 13942
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 10060 12986 10088 13398
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10152 12782 10180 13806
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9692 11286 9720 11562
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9784 11354 9812 11494
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8404 8362 8432 8978
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7760 7002 7788 7278
rect 7856 7100 8152 7120
rect 7912 7098 7936 7100
rect 7992 7098 8016 7100
rect 8072 7098 8096 7100
rect 7934 7046 7936 7098
rect 7998 7046 8010 7098
rect 8072 7046 8074 7098
rect 7912 7044 7936 7046
rect 7992 7044 8016 7046
rect 8072 7044 8096 7046
rect 7856 7024 8152 7044
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7856 6012 8152 6032
rect 7912 6010 7936 6012
rect 7992 6010 8016 6012
rect 8072 6010 8096 6012
rect 7934 5958 7936 6010
rect 7998 5958 8010 6010
rect 8072 5958 8074 6010
rect 7912 5956 7936 5958
rect 7992 5956 8016 5958
rect 8072 5956 8096 5958
rect 7856 5936 8152 5956
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8312 5370 8340 5714
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7576 4826 7604 5102
rect 7856 4924 8152 4944
rect 7912 4922 7936 4924
rect 7992 4922 8016 4924
rect 8072 4922 8096 4924
rect 7934 4870 7936 4922
rect 7998 4870 8010 4922
rect 8072 4870 8074 4922
rect 7912 4868 7936 4870
rect 7992 4868 8016 4870
rect 8072 4868 8096 4870
rect 7856 4848 8152 4868
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7472 4752 7524 4758
rect 7472 4694 7524 4700
rect 7576 4146 7604 4762
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7856 3836 8152 3856
rect 7912 3834 7936 3836
rect 7992 3834 8016 3836
rect 8072 3834 8096 3836
rect 7934 3782 7936 3834
rect 7998 3782 8010 3834
rect 8072 3782 8074 3834
rect 7912 3780 7936 3782
rect 7992 3780 8016 3782
rect 8072 3780 8096 3782
rect 7856 3760 8152 3780
rect 8220 3398 8248 4558
rect 8312 4282 8340 5306
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8496 3058 8524 4558
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8772 2990 8800 9862
rect 9600 9042 9628 10406
rect 9692 9450 9720 10610
rect 9784 10062 9812 11290
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9600 8634 9628 8978
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 9232 7274 9260 8298
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7342 9536 7686
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 9692 6730 9720 9386
rect 9772 8900 9824 8906
rect 9876 8888 9904 10950
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9968 9178 9996 9318
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 10060 9042 10088 11222
rect 10244 11014 10272 13330
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10336 11762 10364 12922
rect 10428 12238 10456 14894
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10428 11286 10456 12174
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10232 9988 10284 9994
rect 10232 9930 10284 9936
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9824 8860 9904 8888
rect 9772 8842 9824 8848
rect 9784 8498 9812 8842
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 10060 8430 10088 8978
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9692 5794 9720 6666
rect 9692 5766 9812 5794
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9692 5166 9720 5578
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8956 3738 8984 3878
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9692 3602 9720 5102
rect 9784 4622 9812 5766
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9784 4146 9812 4558
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9876 4078 9904 8230
rect 10152 6866 10180 9318
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10152 6322 10180 6802
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10244 5166 10272 9930
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10336 6934 10364 7890
rect 10324 6928 10376 6934
rect 10324 6870 10376 6876
rect 10336 6118 10364 6870
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10244 4690 10272 5102
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9048 3194 9076 3470
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 9048 2990 9076 3130
rect 9692 2990 9720 3538
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7856 2748 8152 2768
rect 7912 2746 7936 2748
rect 7992 2746 8016 2748
rect 8072 2746 8096 2748
rect 7934 2694 7936 2746
rect 7998 2694 8010 2746
rect 8072 2694 8074 2746
rect 7912 2692 7936 2694
rect 7992 2692 8016 2694
rect 8072 2692 8096 2694
rect 7856 2672 8152 2692
rect 9784 2650 9812 3878
rect 10428 3738 10456 11018
rect 10520 9586 10548 17224
rect 10980 17066 11008 18158
rect 11072 17202 11100 22646
rect 11716 22574 11744 23038
rect 12912 22574 12940 24323
rect 14752 22574 14780 24323
rect 16592 22574 16620 24323
rect 17972 22574 18000 24323
rect 18206 22876 18502 22896
rect 18262 22874 18286 22876
rect 18342 22874 18366 22876
rect 18422 22874 18446 22876
rect 18284 22822 18286 22874
rect 18348 22822 18360 22874
rect 18422 22822 18424 22874
rect 18262 22820 18286 22822
rect 18342 22820 18366 22822
rect 18422 22820 18446 22822
rect 18206 22800 18502 22820
rect 19812 22574 19840 24323
rect 21086 23216 21142 23225
rect 21086 23151 21142 23160
rect 11704 22568 11756 22574
rect 11704 22510 11756 22516
rect 12900 22568 12952 22574
rect 12900 22510 12952 22516
rect 14740 22568 14792 22574
rect 14740 22510 14792 22516
rect 16580 22568 16632 22574
rect 16580 22510 16632 22516
rect 17960 22568 18012 22574
rect 17960 22510 18012 22516
rect 19800 22568 19852 22574
rect 19800 22510 19852 22516
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 12716 22432 12768 22438
rect 12716 22374 12768 22380
rect 14648 22432 14700 22438
rect 14648 22374 14700 22380
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 19156 22432 19208 22438
rect 19156 22374 19208 22380
rect 11888 22160 11940 22166
rect 11888 22102 11940 22108
rect 11704 22092 11756 22098
rect 11704 22034 11756 22040
rect 11306 21788 11602 21808
rect 11362 21786 11386 21788
rect 11442 21786 11466 21788
rect 11522 21786 11546 21788
rect 11384 21734 11386 21786
rect 11448 21734 11460 21786
rect 11522 21734 11524 21786
rect 11362 21732 11386 21734
rect 11442 21732 11466 21734
rect 11522 21732 11546 21734
rect 11306 21712 11602 21732
rect 11716 21146 11744 22034
rect 11704 21140 11756 21146
rect 11704 21082 11756 21088
rect 11796 20800 11848 20806
rect 11796 20742 11848 20748
rect 11306 20700 11602 20720
rect 11362 20698 11386 20700
rect 11442 20698 11466 20700
rect 11522 20698 11546 20700
rect 11384 20646 11386 20698
rect 11448 20646 11460 20698
rect 11522 20646 11524 20698
rect 11362 20644 11386 20646
rect 11442 20644 11466 20646
rect 11522 20644 11546 20646
rect 11306 20624 11602 20644
rect 11808 20466 11836 20742
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11900 20398 11928 22102
rect 11980 22092 12032 22098
rect 12164 22092 12216 22098
rect 12032 22052 12112 22080
rect 11980 22034 12032 22040
rect 12084 21350 12112 22052
rect 12164 22034 12216 22040
rect 12072 21344 12124 21350
rect 12072 21286 12124 21292
rect 11980 21140 12032 21146
rect 11980 21082 12032 21088
rect 11992 21010 12020 21082
rect 12084 21078 12112 21286
rect 12176 21146 12204 22034
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12268 21554 12296 21830
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 12072 21072 12124 21078
rect 12072 21014 12124 21020
rect 11980 21004 12032 21010
rect 11980 20946 12032 20952
rect 11888 20392 11940 20398
rect 11888 20334 11940 20340
rect 11992 20330 12020 20946
rect 12084 20602 12112 21014
rect 12164 21004 12216 21010
rect 12164 20946 12216 20952
rect 12072 20596 12124 20602
rect 12072 20538 12124 20544
rect 12176 20534 12204 20946
rect 12164 20528 12216 20534
rect 12164 20470 12216 20476
rect 11980 20324 12032 20330
rect 11980 20266 12032 20272
rect 11306 19612 11602 19632
rect 11362 19610 11386 19612
rect 11442 19610 11466 19612
rect 11522 19610 11546 19612
rect 11384 19558 11386 19610
rect 11448 19558 11460 19610
rect 11522 19558 11524 19610
rect 11362 19556 11386 19558
rect 11442 19556 11466 19558
rect 11522 19556 11546 19558
rect 11306 19536 11602 19556
rect 11306 18524 11602 18544
rect 11362 18522 11386 18524
rect 11442 18522 11466 18524
rect 11522 18522 11546 18524
rect 11384 18470 11386 18522
rect 11448 18470 11460 18522
rect 11522 18470 11524 18522
rect 11362 18468 11386 18470
rect 11442 18468 11466 18470
rect 11522 18468 11546 18470
rect 11306 18448 11602 18468
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 11306 17436 11602 17456
rect 11362 17434 11386 17436
rect 11442 17434 11466 17436
rect 11522 17434 11546 17436
rect 11384 17382 11386 17434
rect 11448 17382 11460 17434
rect 11522 17382 11524 17434
rect 11362 17380 11386 17382
rect 11442 17380 11466 17382
rect 11522 17380 11546 17382
rect 11306 17360 11602 17380
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 12176 17134 12204 17682
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10980 16046 11008 17002
rect 11306 16348 11602 16368
rect 11362 16346 11386 16348
rect 11442 16346 11466 16348
rect 11522 16346 11546 16348
rect 11384 16294 11386 16346
rect 11448 16294 11460 16346
rect 11522 16294 11524 16346
rect 11362 16292 11386 16294
rect 11442 16292 11466 16294
rect 11522 16292 11546 16294
rect 11306 16272 11602 16292
rect 12176 16250 12204 17070
rect 12268 16658 12296 17138
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12360 16130 12388 22374
rect 12532 20528 12584 20534
rect 12532 20470 12584 20476
rect 12544 18834 12572 20470
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12452 17338 12480 17614
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12452 16794 12480 17274
rect 12544 17270 12572 18634
rect 12636 18222 12664 19110
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12532 17264 12584 17270
rect 12532 17206 12584 17212
rect 12636 17202 12664 17682
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12268 16102 12388 16130
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11256 15638 11284 15846
rect 11244 15632 11296 15638
rect 11244 15574 11296 15580
rect 11306 15260 11602 15280
rect 11362 15258 11386 15260
rect 11442 15258 11466 15260
rect 11522 15258 11546 15260
rect 11384 15206 11386 15258
rect 11448 15206 11460 15258
rect 11522 15206 11524 15258
rect 11362 15204 11386 15206
rect 11442 15204 11466 15206
rect 11522 15204 11546 15206
rect 11306 15184 11602 15204
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 11306 14172 11602 14192
rect 11362 14170 11386 14172
rect 11442 14170 11466 14172
rect 11522 14170 11546 14172
rect 11384 14118 11386 14170
rect 11448 14118 11460 14170
rect 11522 14118 11524 14170
rect 11362 14116 11386 14118
rect 11442 14116 11466 14118
rect 11522 14116 11546 14118
rect 11306 14096 11602 14116
rect 12084 13462 12112 14826
rect 12268 14822 12296 16102
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12360 15638 12388 15982
rect 12348 15632 12400 15638
rect 12348 15574 12400 15580
rect 12544 15570 12572 15982
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11072 12782 11100 13126
rect 11306 13084 11602 13104
rect 11362 13082 11386 13084
rect 11442 13082 11466 13084
rect 11522 13082 11546 13084
rect 11384 13030 11386 13082
rect 11448 13030 11460 13082
rect 11522 13030 11524 13082
rect 11362 13028 11386 13030
rect 11442 13028 11466 13030
rect 11522 13028 11546 13030
rect 11306 13008 11602 13028
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 10612 11082 10640 12718
rect 11072 12442 11100 12718
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 11306 11996 11602 12016
rect 11362 11994 11386 11996
rect 11442 11994 11466 11996
rect 11522 11994 11546 11996
rect 11384 11942 11386 11994
rect 11448 11942 11460 11994
rect 11522 11942 11524 11994
rect 11362 11940 11386 11942
rect 11442 11940 11466 11942
rect 11522 11940 11546 11942
rect 11306 11920 11602 11940
rect 11716 11286 11744 12922
rect 11808 12374 11836 13126
rect 12084 12850 12112 13398
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 12176 12442 12204 13806
rect 12268 12986 12296 13806
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12452 13462 12480 13670
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 12360 11150 12388 12786
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 11306 10908 11602 10928
rect 11362 10906 11386 10908
rect 11442 10906 11466 10908
rect 11522 10906 11546 10908
rect 11384 10854 11386 10906
rect 11448 10854 11460 10906
rect 11522 10854 11524 10906
rect 11362 10852 11386 10854
rect 11442 10852 11466 10854
rect 11522 10852 11546 10854
rect 11306 10832 11602 10852
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11164 9654 11192 9998
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11306 9820 11602 9840
rect 11362 9818 11386 9820
rect 11442 9818 11466 9820
rect 11522 9818 11546 9820
rect 11384 9766 11386 9818
rect 11448 9766 11460 9818
rect 11522 9766 11524 9818
rect 11362 9764 11386 9766
rect 11442 9764 11466 9766
rect 11522 9764 11546 9766
rect 11306 9744 11602 9764
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 11900 9178 11928 9930
rect 12360 9450 12388 11086
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12452 9586 12480 10202
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10704 7342 10732 8978
rect 11306 8732 11602 8752
rect 11362 8730 11386 8732
rect 11442 8730 11466 8732
rect 11522 8730 11546 8732
rect 11384 8678 11386 8730
rect 11448 8678 11460 8730
rect 11522 8678 11524 8730
rect 11362 8676 11386 8678
rect 11442 8676 11466 8678
rect 11522 8676 11546 8678
rect 11306 8656 11602 8676
rect 12360 8362 12388 9386
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12452 8090 12480 8230
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 11306 7644 11602 7664
rect 11362 7642 11386 7644
rect 11442 7642 11466 7644
rect 11522 7642 11546 7644
rect 11384 7590 11386 7642
rect 11448 7590 11460 7642
rect 11522 7590 11524 7642
rect 11362 7588 11386 7590
rect 11442 7588 11466 7590
rect 11522 7588 11546 7590
rect 11306 7568 11602 7588
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10888 6390 10916 6938
rect 10980 6866 11008 7210
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10876 6384 10928 6390
rect 10876 6326 10928 6332
rect 10980 5098 11008 6802
rect 11306 6556 11602 6576
rect 11362 6554 11386 6556
rect 11442 6554 11466 6556
rect 11522 6554 11546 6556
rect 11384 6502 11386 6554
rect 11448 6502 11460 6554
rect 11522 6502 11524 6554
rect 11362 6500 11386 6502
rect 11442 6500 11466 6502
rect 11522 6500 11546 6502
rect 11306 6480 11602 6500
rect 11306 5468 11602 5488
rect 11362 5466 11386 5468
rect 11442 5466 11466 5468
rect 11522 5466 11546 5468
rect 11384 5414 11386 5466
rect 11448 5414 11460 5466
rect 11522 5414 11524 5466
rect 11362 5412 11386 5414
rect 11442 5412 11466 5414
rect 11522 5412 11546 5414
rect 11306 5392 11602 5412
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10980 4758 11008 5034
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 10060 3194 10088 3674
rect 10520 3670 10548 4082
rect 11072 3942 11100 5102
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 11306 4380 11602 4400
rect 11362 4378 11386 4380
rect 11442 4378 11466 4380
rect 11522 4378 11546 4380
rect 11384 4326 11386 4378
rect 11448 4326 11460 4378
rect 11522 4326 11524 4378
rect 11362 4324 11386 4326
rect 11442 4324 11466 4326
rect 11522 4324 11546 4326
rect 11306 4304 11602 4324
rect 12176 4282 12204 4626
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 11704 4004 11756 4010
rect 11704 3946 11756 3952
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10888 2990 10916 3334
rect 11164 3194 11192 3878
rect 11306 3292 11602 3312
rect 11362 3290 11386 3292
rect 11442 3290 11466 3292
rect 11522 3290 11546 3292
rect 11384 3238 11386 3290
rect 11448 3238 11460 3290
rect 11522 3238 11524 3290
rect 11362 3236 11386 3238
rect 11442 3236 11466 3238
rect 11522 3236 11546 3238
rect 11306 3216 11602 3236
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 2044 2576 2096 2582
rect 2044 2518 2096 2524
rect 10888 2514 10916 2926
rect 11164 2650 11192 3130
rect 11716 2990 11744 3946
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 1872 800 1900 2314
rect 3712 800 3740 2450
rect 4406 2204 4702 2224
rect 4462 2202 4486 2204
rect 4542 2202 4566 2204
rect 4622 2202 4646 2204
rect 4484 2150 4486 2202
rect 4548 2150 4560 2202
rect 4622 2150 4624 2202
rect 4462 2148 4486 2150
rect 4542 2148 4566 2150
rect 4622 2148 4646 2150
rect 4406 2128 4702 2148
rect 5552 800 5580 2450
rect 6932 800 6960 2450
rect 8772 800 8800 2450
rect 10612 800 10640 2450
rect 11306 2204 11602 2224
rect 11362 2202 11386 2204
rect 11442 2202 11466 2204
rect 11522 2202 11546 2204
rect 11384 2150 11386 2202
rect 11448 2150 11460 2202
rect 11522 2150 11524 2202
rect 11362 2148 11386 2150
rect 11442 2148 11466 2150
rect 11522 2148 11546 2150
rect 11306 2128 11602 2148
rect 11992 800 12020 3470
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 12084 2514 12112 3334
rect 12544 3194 12572 15506
rect 12636 15162 12664 17138
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12636 10674 12664 12582
rect 12728 11354 12756 22374
rect 12900 22092 12952 22098
rect 12900 22034 12952 22040
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12820 21418 12848 21830
rect 12808 21412 12860 21418
rect 12808 21354 12860 21360
rect 12912 19922 12940 22034
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14292 21078 14320 21286
rect 14280 21072 14332 21078
rect 14280 21014 14332 21020
rect 14292 20534 14320 21014
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 14292 20398 14320 20470
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14464 20324 14516 20330
rect 14464 20266 14516 20272
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 12900 19916 12952 19922
rect 12900 19858 12952 19864
rect 14292 19310 14320 20198
rect 14476 19990 14504 20266
rect 14464 19984 14516 19990
rect 14464 19926 14516 19932
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12820 18902 12848 19178
rect 13648 19174 13676 19246
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13004 18902 13032 19110
rect 12808 18896 12860 18902
rect 12808 18838 12860 18844
rect 12992 18896 13044 18902
rect 12992 18838 13044 18844
rect 13004 18358 13032 18838
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 12992 18352 13044 18358
rect 12992 18294 13044 18300
rect 13556 18222 13584 18566
rect 13740 18358 13768 18770
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 13544 18216 13596 18222
rect 13544 18158 13596 18164
rect 12808 17604 12860 17610
rect 12808 17546 12860 17552
rect 12820 17202 12848 17546
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 13004 16114 13032 18158
rect 13188 17882 13216 18158
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 14476 17746 14504 19926
rect 14568 19310 14596 20402
rect 14660 19938 14688 22374
rect 14756 22332 15052 22352
rect 14812 22330 14836 22332
rect 14892 22330 14916 22332
rect 14972 22330 14996 22332
rect 14834 22278 14836 22330
rect 14898 22278 14910 22330
rect 14972 22278 14974 22330
rect 14812 22276 14836 22278
rect 14892 22276 14916 22278
rect 14972 22276 14996 22278
rect 14756 22256 15052 22276
rect 15292 21956 15344 21962
rect 15292 21898 15344 21904
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 15212 21418 15240 21830
rect 15200 21412 15252 21418
rect 15200 21354 15252 21360
rect 14756 21244 15052 21264
rect 14812 21242 14836 21244
rect 14892 21242 14916 21244
rect 14972 21242 14996 21244
rect 14834 21190 14836 21242
rect 14898 21190 14910 21242
rect 14972 21190 14974 21242
rect 14812 21188 14836 21190
rect 14892 21188 14916 21190
rect 14972 21188 14996 21190
rect 14756 21168 15052 21188
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 14936 20330 14964 20402
rect 14924 20324 14976 20330
rect 14924 20266 14976 20272
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 14756 20156 15052 20176
rect 14812 20154 14836 20156
rect 14892 20154 14916 20156
rect 14972 20154 14996 20156
rect 14834 20102 14836 20154
rect 14898 20102 14910 20154
rect 14972 20102 14974 20154
rect 14812 20100 14836 20102
rect 14892 20100 14916 20102
rect 14972 20100 14996 20102
rect 14756 20080 15052 20100
rect 14660 19910 14780 19938
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14660 19378 14688 19654
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14752 19310 14780 19910
rect 15108 19916 15160 19922
rect 15108 19858 15160 19864
rect 14556 19304 14608 19310
rect 14556 19246 14608 19252
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 15120 19242 15148 19858
rect 15212 19854 15240 20198
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15212 19310 15240 19790
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15108 19236 15160 19242
rect 15108 19178 15160 19184
rect 14756 19068 15052 19088
rect 14812 19066 14836 19068
rect 14892 19066 14916 19068
rect 14972 19066 14996 19068
rect 14834 19014 14836 19066
rect 14898 19014 14910 19066
rect 14972 19014 14974 19066
rect 14812 19012 14836 19014
rect 14892 19012 14916 19014
rect 14972 19012 14996 19014
rect 14756 18992 15052 19012
rect 14756 17980 15052 18000
rect 14812 17978 14836 17980
rect 14892 17978 14916 17980
rect 14972 17978 14996 17980
rect 14834 17926 14836 17978
rect 14898 17926 14910 17978
rect 14972 17926 14974 17978
rect 14812 17924 14836 17926
rect 14892 17924 14916 17926
rect 14972 17924 14996 17926
rect 14756 17904 15052 17924
rect 14648 17808 14700 17814
rect 14648 17750 14700 17756
rect 14464 17740 14516 17746
rect 14464 17682 14516 17688
rect 14476 16794 14504 17682
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 13912 16448 13964 16454
rect 13912 16390 13964 16396
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13004 15638 13032 16050
rect 12992 15632 13044 15638
rect 12992 15574 13044 15580
rect 13924 15570 13952 16390
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 14476 14550 14504 16730
rect 14660 16726 14688 17750
rect 14756 16892 15052 16912
rect 14812 16890 14836 16892
rect 14892 16890 14916 16892
rect 14972 16890 14996 16892
rect 14834 16838 14836 16890
rect 14898 16838 14910 16890
rect 14972 16838 14974 16890
rect 14812 16836 14836 16838
rect 14892 16836 14916 16838
rect 14972 16836 14996 16838
rect 14756 16816 15052 16836
rect 14648 16720 14700 16726
rect 14648 16662 14700 16668
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 14936 16250 14964 16594
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 15028 16114 15056 16594
rect 15120 16182 15148 19178
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 15212 17338 15240 17750
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15212 16658 15240 17274
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15108 16176 15160 16182
rect 15108 16118 15160 16124
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 15212 16046 15240 16594
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 14568 15502 14596 15982
rect 15212 15910 15240 15982
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 14756 15804 15052 15824
rect 14812 15802 14836 15804
rect 14892 15802 14916 15804
rect 14972 15802 14996 15804
rect 14834 15750 14836 15802
rect 14898 15750 14910 15802
rect 14972 15750 14974 15802
rect 14812 15748 14836 15750
rect 14892 15748 14916 15750
rect 14972 15748 14996 15750
rect 14756 15728 15052 15748
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14568 14618 14596 15438
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 15016 14952 15068 14958
rect 15068 14900 15240 14906
rect 15016 14894 15240 14900
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14464 14544 14516 14550
rect 14660 14498 14688 14894
rect 15028 14878 15240 14894
rect 15212 14822 15240 14878
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 14756 14716 15052 14736
rect 14812 14714 14836 14716
rect 14892 14714 14916 14716
rect 14972 14714 14996 14716
rect 14834 14662 14836 14714
rect 14898 14662 14910 14714
rect 14972 14662 14974 14714
rect 14812 14660 14836 14662
rect 14892 14660 14916 14662
rect 14972 14660 14996 14662
rect 14756 14640 15052 14660
rect 14464 14486 14516 14492
rect 14280 14340 14332 14346
rect 14280 14282 14332 14288
rect 14292 13870 14320 14282
rect 14476 13938 14504 14486
rect 14568 14482 14688 14498
rect 15212 14482 15240 14758
rect 14556 14476 14688 14482
rect 14608 14470 14688 14476
rect 15200 14476 15252 14482
rect 14556 14418 14608 14424
rect 15200 14418 15252 14424
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14568 13870 14596 14418
rect 15212 13870 15240 14418
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 14556 13864 14608 13870
rect 14556 13806 14608 13812
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 13096 12782 13124 13194
rect 13832 12850 13860 13262
rect 14108 12850 14136 13670
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 13004 12442 13032 12582
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12636 10130 12664 10610
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 13004 9518 13032 10066
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 13004 9042 13032 9454
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12636 8362 12664 8910
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 12636 7886 12664 8298
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13280 7410 13308 7686
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12636 5098 12664 5510
rect 12728 5370 12756 5714
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12636 3602 12664 5034
rect 13176 3664 13228 3670
rect 13176 3606 13228 3612
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12636 3058 12664 3538
rect 13188 3058 13216 3606
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 13372 2938 13400 9862
rect 13464 9722 13492 10542
rect 13832 10198 13860 10746
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 14200 8498 14228 13126
rect 14568 12986 14596 13806
rect 14756 13628 15052 13648
rect 14812 13626 14836 13628
rect 14892 13626 14916 13628
rect 14972 13626 14996 13628
rect 14834 13574 14836 13626
rect 14898 13574 14910 13626
rect 14972 13574 14974 13626
rect 14812 13572 14836 13574
rect 14892 13572 14916 13574
rect 14972 13572 14996 13574
rect 14756 13552 15052 13572
rect 15212 13462 15240 13806
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 15108 12708 15160 12714
rect 15108 12650 15160 12656
rect 14756 12540 15052 12560
rect 14812 12538 14836 12540
rect 14892 12538 14916 12540
rect 14972 12538 14996 12540
rect 14834 12486 14836 12538
rect 14898 12486 14910 12538
rect 14972 12486 14974 12538
rect 14812 12484 14836 12486
rect 14892 12484 14916 12486
rect 14972 12484 14996 12486
rect 14756 12464 15052 12484
rect 15120 12442 15148 12650
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 14756 11452 15052 11472
rect 14812 11450 14836 11452
rect 14892 11450 14916 11452
rect 14972 11450 14996 11452
rect 14834 11398 14836 11450
rect 14898 11398 14910 11450
rect 14972 11398 14974 11450
rect 14812 11396 14836 11398
rect 14892 11396 14916 11398
rect 14972 11396 14996 11398
rect 14756 11376 15052 11396
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14844 10606 14872 11018
rect 15028 10810 15056 11154
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 15212 10606 15240 11018
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 14756 10364 15052 10384
rect 14812 10362 14836 10364
rect 14892 10362 14916 10364
rect 14972 10362 14996 10364
rect 14834 10310 14836 10362
rect 14898 10310 14910 10362
rect 14972 10310 14974 10362
rect 14812 10308 14836 10310
rect 14892 10308 14916 10310
rect 14972 10308 14996 10310
rect 14756 10288 15052 10308
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14200 7954 14228 8434
rect 14292 8430 14320 9454
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 14756 9276 15052 9296
rect 14812 9274 14836 9276
rect 14892 9274 14916 9276
rect 14972 9274 14996 9276
rect 14834 9222 14836 9274
rect 14898 9222 14910 9274
rect 14972 9222 14974 9274
rect 14812 9220 14836 9222
rect 14892 9220 14916 9222
rect 14972 9220 14996 9222
rect 14756 9200 15052 9220
rect 15212 9178 15240 9318
rect 15304 9178 15332 21898
rect 16212 21548 16264 21554
rect 16212 21490 16264 21496
rect 15752 21412 15804 21418
rect 15752 21354 15804 21360
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15488 21010 15516 21286
rect 15764 21146 15792 21354
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 16224 21010 16252 21490
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 16212 21004 16264 21010
rect 16212 20946 16264 20952
rect 15384 20868 15436 20874
rect 15384 20810 15436 20816
rect 15396 19990 15424 20810
rect 15384 19984 15436 19990
rect 15384 19926 15436 19932
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 15396 19514 15424 19790
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 15488 18834 15516 20946
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15672 20806 15700 20878
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 15672 20398 15700 20742
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 15660 20392 15712 20398
rect 15660 20334 15712 20340
rect 15672 18834 15700 20334
rect 16224 20058 16252 20402
rect 16212 20052 16264 20058
rect 16212 19994 16264 20000
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 15660 18828 15712 18834
rect 15660 18770 15712 18776
rect 15488 17746 15516 18770
rect 15672 18086 15700 18770
rect 15764 18766 15792 19858
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 15764 18426 15792 18702
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15396 14482 15424 14826
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15488 14346 15516 17682
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 15948 17202 15976 17478
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 16040 14482 16068 14758
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 16224 12782 16252 16934
rect 16316 13258 16344 22374
rect 17500 22092 17552 22098
rect 17500 22034 17552 22040
rect 17224 21072 17276 21078
rect 17224 21014 17276 21020
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16500 19786 16528 20878
rect 17236 20602 17264 21014
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 17512 20398 17540 22034
rect 17972 21418 18000 22374
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18206 21788 18502 21808
rect 18262 21786 18286 21788
rect 18342 21786 18366 21788
rect 18422 21786 18446 21788
rect 18284 21734 18286 21786
rect 18348 21734 18360 21786
rect 18422 21734 18424 21786
rect 18262 21732 18286 21734
rect 18342 21732 18366 21734
rect 18422 21732 18446 21734
rect 18206 21712 18502 21732
rect 18708 21418 18736 21830
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 17960 21412 18012 21418
rect 17960 21354 18012 21360
rect 18696 21412 18748 21418
rect 18696 21354 18748 21360
rect 18206 20700 18502 20720
rect 18262 20698 18286 20700
rect 18342 20698 18366 20700
rect 18422 20698 18446 20700
rect 18284 20646 18286 20698
rect 18348 20646 18360 20698
rect 18422 20646 18424 20698
rect 18262 20644 18286 20646
rect 18342 20644 18366 20646
rect 18422 20644 18446 20646
rect 18206 20624 18502 20644
rect 19076 20398 19104 21490
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 16488 19780 16540 19786
rect 16488 19722 16540 19728
rect 17512 19310 17540 20334
rect 18206 19612 18502 19632
rect 18262 19610 18286 19612
rect 18342 19610 18366 19612
rect 18422 19610 18446 19612
rect 18284 19558 18286 19610
rect 18348 19558 18360 19610
rect 18422 19558 18424 19610
rect 18262 19556 18286 19558
rect 18342 19556 18366 19558
rect 18422 19556 18446 19558
rect 18206 19536 18502 19556
rect 19076 19310 19104 20334
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 17696 18902 17724 19110
rect 17684 18896 17736 18902
rect 16500 18834 16988 18850
rect 17684 18838 17736 18844
rect 16488 18828 16988 18834
rect 16540 18822 16988 18828
rect 16488 18770 16540 18776
rect 16960 18766 16988 18822
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 16592 18290 16620 18702
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16684 17202 16712 18634
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17132 18216 17184 18222
rect 17132 18158 17184 18164
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 17052 16114 17080 17138
rect 17144 16658 17172 18158
rect 17236 16726 17264 18226
rect 17328 18222 17356 18702
rect 17316 18216 17368 18222
rect 17316 18158 17368 18164
rect 17316 18080 17368 18086
rect 17316 18022 17368 18028
rect 17224 16720 17276 16726
rect 17224 16662 17276 16668
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16408 12986 16436 13330
rect 17052 13326 17080 16050
rect 17144 16046 17172 16594
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17144 15570 17172 15982
rect 17236 15570 17264 16662
rect 17328 16658 17356 18022
rect 17788 17202 17816 19246
rect 19168 18698 19196 22374
rect 21100 22098 21128 23151
rect 21652 22574 21680 24323
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 21180 22432 21232 22438
rect 21180 22374 21232 22380
rect 20536 22092 20588 22098
rect 20536 22034 20588 22040
rect 21088 22092 21140 22098
rect 21088 22034 21140 22040
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19352 20466 19380 21286
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 20088 20330 20116 21830
rect 20168 21616 20220 21622
rect 20168 21558 20220 21564
rect 20180 21486 20208 21558
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 20076 20324 20128 20330
rect 20076 20266 20128 20272
rect 20180 20262 20208 21422
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 19628 19378 19656 20198
rect 20548 19922 20576 22034
rect 21088 21480 21140 21486
rect 21088 21422 21140 21428
rect 20812 21004 20864 21010
rect 20812 20946 20864 20952
rect 20628 20800 20680 20806
rect 20628 20742 20680 20748
rect 20640 20505 20668 20742
rect 20626 20496 20682 20505
rect 20626 20431 20682 20440
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 20364 19242 20392 19654
rect 20352 19236 20404 19242
rect 20352 19178 20404 19184
rect 19984 18896 20036 18902
rect 19984 18838 20036 18844
rect 20536 18896 20588 18902
rect 20536 18838 20588 18844
rect 19156 18692 19208 18698
rect 19156 18634 19208 18640
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 18206 18524 18502 18544
rect 18262 18522 18286 18524
rect 18342 18522 18366 18524
rect 18422 18522 18446 18524
rect 18284 18470 18286 18522
rect 18348 18470 18360 18522
rect 18422 18470 18424 18522
rect 18262 18468 18286 18470
rect 18342 18468 18366 18470
rect 18422 18468 18446 18470
rect 18206 18448 18502 18468
rect 19076 18426 19104 18566
rect 19064 18420 19116 18426
rect 19064 18362 19116 18368
rect 19168 18222 19196 18634
rect 19996 18290 20024 18838
rect 20352 18828 20404 18834
rect 20352 18770 20404 18776
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19156 18216 19208 18222
rect 19156 18158 19208 18164
rect 19616 18216 19668 18222
rect 19616 18158 19668 18164
rect 19628 18086 19656 18158
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 18206 17436 18502 17456
rect 18262 17434 18286 17436
rect 18342 17434 18366 17436
rect 18422 17434 18446 17436
rect 18284 17382 18286 17434
rect 18348 17382 18360 17434
rect 18422 17382 18424 17434
rect 18262 17380 18286 17382
rect 18342 17380 18366 17382
rect 18422 17380 18446 17382
rect 18206 17360 18502 17380
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 19616 17060 19668 17066
rect 19616 17002 19668 17008
rect 17868 16992 17920 16998
rect 17868 16934 17920 16940
rect 17880 16658 17908 16934
rect 19628 16794 19656 17002
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17328 15706 17356 16594
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 17604 16114 17632 16390
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 18064 15978 18092 16390
rect 18206 16348 18502 16368
rect 18262 16346 18286 16348
rect 18342 16346 18366 16348
rect 18422 16346 18446 16348
rect 18284 16294 18286 16346
rect 18348 16294 18360 16346
rect 18422 16294 18424 16346
rect 18262 16292 18286 16294
rect 18342 16292 18366 16294
rect 18422 16292 18446 16294
rect 18206 16272 18502 16292
rect 19260 16114 19288 16730
rect 19524 16720 19576 16726
rect 19524 16662 19576 16668
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 18052 15972 18104 15978
rect 18052 15914 18104 15920
rect 19260 15910 19288 16050
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17236 14618 17264 15506
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17696 14346 17724 15506
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17328 13462 17356 13670
rect 17316 13456 17368 13462
rect 17316 13398 17368 13404
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17420 13190 17448 14214
rect 17696 13870 17724 14282
rect 17788 13870 17816 15302
rect 18206 15260 18502 15280
rect 18262 15258 18286 15260
rect 18342 15258 18366 15260
rect 18422 15258 18446 15260
rect 18284 15206 18286 15258
rect 18348 15206 18360 15258
rect 18422 15206 18424 15258
rect 18262 15204 18286 15206
rect 18342 15204 18366 15206
rect 18422 15204 18446 15206
rect 18206 15184 18502 15204
rect 19260 15162 19288 15846
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 18064 13954 18092 14418
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18206 14172 18502 14192
rect 18262 14170 18286 14172
rect 18342 14170 18366 14172
rect 18422 14170 18446 14172
rect 18284 14118 18286 14170
rect 18348 14118 18360 14170
rect 18422 14118 18424 14170
rect 18262 14116 18286 14118
rect 18342 14116 18366 14118
rect 18422 14116 18446 14118
rect 18206 14096 18502 14116
rect 18064 13938 18184 13954
rect 18064 13932 18196 13938
rect 18064 13926 18144 13932
rect 18144 13874 18196 13880
rect 17500 13864 17552 13870
rect 17500 13806 17552 13812
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 17420 12850 17448 13126
rect 17512 12986 17540 13806
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17696 12918 17724 13262
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16224 12306 16252 12718
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16500 10130 16528 11086
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16868 10742 16896 10950
rect 16856 10736 16908 10742
rect 16856 10678 16908 10684
rect 16960 10198 16988 11154
rect 17696 10606 17724 12854
rect 17788 12714 17816 13806
rect 18064 13394 18092 13806
rect 18156 13530 18184 13874
rect 18708 13870 18736 14214
rect 18892 13870 18920 15098
rect 19352 14958 19380 16118
rect 19536 16046 19564 16662
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19800 16040 19852 16046
rect 19800 15982 19852 15988
rect 19812 15638 19840 15982
rect 19800 15632 19852 15638
rect 19800 15574 19852 15580
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19352 13954 19380 14894
rect 18984 13938 19380 13954
rect 18972 13932 19380 13938
rect 19024 13926 19380 13932
rect 18972 13874 19024 13880
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18604 13728 18656 13734
rect 18604 13670 18656 13676
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 18064 12782 18092 13330
rect 18206 13084 18502 13104
rect 18262 13082 18286 13084
rect 18342 13082 18366 13084
rect 18422 13082 18446 13084
rect 18284 13030 18286 13082
rect 18348 13030 18360 13082
rect 18422 13030 18424 13082
rect 18262 13028 18286 13030
rect 18342 13028 18366 13030
rect 18422 13028 18446 13030
rect 18206 13008 18502 13028
rect 18616 12782 18644 13670
rect 18892 13190 18920 13806
rect 19904 13462 19932 16526
rect 19996 16250 20024 18226
rect 20272 18222 20300 18566
rect 20260 18216 20312 18222
rect 20260 18158 20312 18164
rect 20364 18086 20392 18770
rect 20548 18358 20576 18838
rect 20536 18352 20588 18358
rect 20536 18294 20588 18300
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 20272 16726 20300 16934
rect 20260 16720 20312 16726
rect 20260 16662 20312 16668
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 20076 16584 20128 16590
rect 20076 16526 20128 16532
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19984 15564 20036 15570
rect 19984 15506 20036 15512
rect 19996 14958 20024 15506
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 20088 13802 20116 16526
rect 20180 16182 20208 16594
rect 20168 16176 20220 16182
rect 20168 16118 20220 16124
rect 20168 15564 20220 15570
rect 20168 15506 20220 15512
rect 20180 14958 20208 15506
rect 20364 15162 20392 18022
rect 20548 15994 20576 18294
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 20640 17785 20668 18158
rect 20626 17776 20682 17785
rect 20626 17711 20682 17720
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20732 17134 20760 17478
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20824 16674 20852 20946
rect 21100 19514 21128 21422
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 20996 18080 21048 18086
rect 20996 18022 21048 18028
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20456 15966 20576 15994
rect 20732 16646 20852 16674
rect 20456 15706 20484 15966
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20548 15570 20576 15846
rect 20536 15564 20588 15570
rect 20536 15506 20588 15512
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20260 15020 20312 15026
rect 20260 14962 20312 14968
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 20180 14618 20208 14894
rect 20272 14618 20300 14962
rect 20444 14884 20496 14890
rect 20444 14826 20496 14832
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 20272 14278 20300 14554
rect 20456 14482 20484 14826
rect 20444 14476 20496 14482
rect 20444 14418 20496 14424
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 20076 13796 20128 13802
rect 20076 13738 20128 13744
rect 19892 13456 19944 13462
rect 19892 13398 19944 13404
rect 20088 13394 20116 13738
rect 20272 13394 20300 14214
rect 20456 13938 20484 14418
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20456 13394 20484 13874
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20076 13388 20128 13394
rect 20076 13330 20128 13336
rect 20260 13388 20312 13394
rect 20260 13330 20312 13336
rect 20444 13388 20496 13394
rect 20444 13330 20496 13336
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 19616 13184 19668 13190
rect 19616 13126 19668 13132
rect 18892 12850 18920 13126
rect 19628 12850 19656 13126
rect 20272 12986 20300 13330
rect 20260 12980 20312 12986
rect 20260 12922 20312 12928
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 17972 10606 18000 12582
rect 18206 11996 18502 12016
rect 18262 11994 18286 11996
rect 18342 11994 18366 11996
rect 18422 11994 18446 11996
rect 18284 11942 18286 11994
rect 18348 11942 18360 11994
rect 18422 11942 18424 11994
rect 18262 11940 18286 11942
rect 18342 11940 18366 11942
rect 18422 11940 18446 11942
rect 18206 11920 18502 11940
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18144 11280 18196 11286
rect 18196 11228 18368 11234
rect 18144 11222 18368 11228
rect 18156 11206 18368 11222
rect 18432 11218 18460 11494
rect 18340 11150 18368 11206
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17408 10532 17460 10538
rect 17408 10474 17460 10480
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 17328 9110 17356 10406
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14476 8566 14504 8978
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14464 8560 14516 8566
rect 14464 8502 14516 8508
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 8022 14596 8230
rect 14556 8016 14608 8022
rect 14556 7958 14608 7964
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13464 5846 13492 7482
rect 14568 7342 14596 7958
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14660 6322 14688 8774
rect 16592 8634 16620 8910
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 14756 8188 15052 8208
rect 14812 8186 14836 8188
rect 14892 8186 14916 8188
rect 14972 8186 14996 8188
rect 14834 8134 14836 8186
rect 14898 8134 14910 8186
rect 14972 8134 14974 8186
rect 14812 8132 14836 8134
rect 14892 8132 14916 8134
rect 14972 8132 14996 8134
rect 14756 8112 15052 8132
rect 15304 7954 15332 8366
rect 16592 8022 16620 8570
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15304 7410 15332 7890
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 14756 7100 15052 7120
rect 14812 7098 14836 7100
rect 14892 7098 14916 7100
rect 14972 7098 14996 7100
rect 14834 7046 14836 7098
rect 14898 7046 14910 7098
rect 14972 7046 14974 7098
rect 14812 7044 14836 7046
rect 14892 7044 14916 7046
rect 14972 7044 14996 7046
rect 14756 7024 15052 7044
rect 17420 6866 17448 10474
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17788 10130 17816 10406
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 18064 9042 18092 11018
rect 18206 10908 18502 10928
rect 18262 10906 18286 10908
rect 18342 10906 18366 10908
rect 18422 10906 18446 10908
rect 18284 10854 18286 10906
rect 18348 10854 18360 10906
rect 18422 10854 18424 10906
rect 18262 10852 18286 10854
rect 18342 10852 18366 10854
rect 18422 10852 18446 10854
rect 18206 10832 18502 10852
rect 18616 10674 18644 11086
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18708 10062 18736 10950
rect 18892 10674 18920 12582
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 20088 11218 20116 12242
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 20180 10538 20208 11018
rect 20456 10810 20484 13330
rect 20640 13025 20668 13806
rect 20626 13016 20682 13025
rect 20626 12951 20682 12960
rect 20628 12708 20680 12714
rect 20628 12650 20680 12656
rect 20640 12442 20668 12650
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20444 10804 20496 10810
rect 20444 10746 20496 10752
rect 20168 10532 20220 10538
rect 20168 10474 20220 10480
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18206 9820 18502 9840
rect 18262 9818 18286 9820
rect 18342 9818 18366 9820
rect 18422 9818 18446 9820
rect 18284 9766 18286 9818
rect 18348 9766 18360 9818
rect 18422 9766 18424 9818
rect 18262 9764 18286 9766
rect 18342 9764 18366 9766
rect 18422 9764 18446 9766
rect 18206 9744 18502 9764
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 18052 9036 18104 9042
rect 18052 8978 18104 8984
rect 18064 8514 18092 8978
rect 18206 8732 18502 8752
rect 18262 8730 18286 8732
rect 18342 8730 18366 8732
rect 18422 8730 18446 8732
rect 18284 8678 18286 8730
rect 18348 8678 18360 8730
rect 18422 8678 18424 8730
rect 18262 8676 18286 8678
rect 18342 8676 18366 8678
rect 18422 8676 18446 8678
rect 18206 8656 18502 8676
rect 18616 8634 18644 9114
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18064 8486 18184 8514
rect 18156 8430 18184 8486
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 18064 8022 18092 8366
rect 18616 8090 18644 8570
rect 18708 8430 18736 8910
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18052 8016 18104 8022
rect 18052 7958 18104 7964
rect 18206 7644 18502 7664
rect 18262 7642 18286 7644
rect 18342 7642 18366 7644
rect 18422 7642 18446 7644
rect 18284 7590 18286 7642
rect 18348 7590 18360 7642
rect 18422 7590 18424 7642
rect 18262 7588 18286 7590
rect 18342 7588 18366 7590
rect 18422 7588 18446 7590
rect 18206 7568 18502 7588
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 13452 5840 13504 5846
rect 13452 5782 13504 5788
rect 14660 5778 14688 6258
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 14756 6012 15052 6032
rect 14812 6010 14836 6012
rect 14892 6010 14916 6012
rect 14972 6010 14996 6012
rect 14834 5958 14836 6010
rect 14898 5958 14910 6010
rect 14972 5958 14974 6010
rect 14812 5956 14836 5958
rect 14892 5956 14916 5958
rect 14972 5956 14996 5958
rect 14756 5936 15052 5956
rect 14832 5840 14884 5846
rect 14832 5782 14884 5788
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14844 5166 14872 5782
rect 15120 5370 15148 6190
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15212 5846 15240 6054
rect 15948 5914 15976 6802
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 16224 6322 16252 6734
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 17512 6254 17540 6734
rect 17500 6248 17552 6254
rect 17500 6190 17552 6196
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 15200 5840 15252 5846
rect 15200 5782 15252 5788
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15212 5302 15240 5646
rect 15200 5296 15252 5302
rect 15200 5238 15252 5244
rect 15304 5166 15332 5714
rect 17328 5370 17356 5714
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17512 5166 17540 6190
rect 17696 5846 17724 6190
rect 17684 5840 17736 5846
rect 17684 5782 17736 5788
rect 17788 5234 17816 6938
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17880 6254 17908 6802
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18206 6556 18502 6576
rect 18262 6554 18286 6556
rect 18342 6554 18366 6556
rect 18422 6554 18446 6556
rect 18284 6502 18286 6554
rect 18348 6502 18360 6554
rect 18422 6502 18424 6554
rect 18262 6500 18286 6502
rect 18342 6500 18366 6502
rect 18422 6500 18446 6502
rect 18206 6480 18502 6500
rect 18708 6254 18736 6734
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 17880 5778 17908 6190
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 17500 5160 17552 5166
rect 17500 5102 17552 5108
rect 14756 4924 15052 4944
rect 14812 4922 14836 4924
rect 14892 4922 14916 4924
rect 14972 4922 14996 4924
rect 14834 4870 14836 4922
rect 14898 4870 14910 4922
rect 14972 4870 14974 4922
rect 14812 4868 14836 4870
rect 14892 4868 14916 4870
rect 14972 4868 14996 4870
rect 14756 4848 15052 4868
rect 15304 4214 15332 5102
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 15292 4208 15344 4214
rect 15292 4150 15344 4156
rect 15568 4004 15620 4010
rect 15568 3946 15620 3952
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13924 3126 13952 3538
rect 14660 3194 14688 3878
rect 14756 3836 15052 3856
rect 14812 3834 14836 3836
rect 14892 3834 14916 3836
rect 14972 3834 14996 3836
rect 14834 3782 14836 3834
rect 14898 3782 14910 3834
rect 14972 3782 14974 3834
rect 14812 3780 14836 3782
rect 14892 3780 14916 3782
rect 14972 3780 14996 3782
rect 14756 3760 15052 3780
rect 15396 3670 15424 3878
rect 15580 3738 15608 3946
rect 15568 3732 15620 3738
rect 15568 3674 15620 3680
rect 15384 3664 15436 3670
rect 15384 3606 15436 3612
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15580 3194 15608 3470
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 13912 3120 13964 3126
rect 14660 3074 14688 3130
rect 13912 3062 13964 3068
rect 13372 2910 13492 2938
rect 13464 2854 13492 2910
rect 12900 2848 12952 2854
rect 12900 2790 12952 2796
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 12912 2650 12940 2790
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13832 2582 13860 2790
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 13924 2514 13952 3062
rect 14568 3046 14688 3074
rect 16040 3058 16068 3334
rect 17328 3058 17356 4422
rect 16028 3052 16080 3058
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14292 2582 14320 2926
rect 14280 2576 14332 2582
rect 14280 2518 14332 2524
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 13832 800 13860 2382
rect 14568 2310 14596 3046
rect 16028 2994 16080 3000
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 14660 2650 14688 2926
rect 14756 2748 15052 2768
rect 14812 2746 14836 2748
rect 14892 2746 14916 2748
rect 14972 2746 14996 2748
rect 14834 2694 14836 2746
rect 14898 2694 14910 2746
rect 14972 2694 14974 2746
rect 14812 2692 14836 2694
rect 14892 2692 14916 2694
rect 14972 2692 14996 2694
rect 14756 2672 15052 2692
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 15660 2508 15712 2514
rect 15660 2450 15712 2456
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 15672 800 15700 2450
rect 16132 2446 16160 2994
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 17052 800 17080 2450
rect 17512 2310 17540 5102
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17696 4826 17724 4966
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 17788 4486 17816 4966
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17880 2582 17908 5714
rect 18206 5468 18502 5488
rect 18262 5466 18286 5468
rect 18342 5466 18366 5468
rect 18422 5466 18446 5468
rect 18284 5414 18286 5466
rect 18348 5414 18360 5466
rect 18422 5414 18424 5466
rect 18262 5412 18286 5414
rect 18342 5412 18366 5414
rect 18422 5412 18446 5414
rect 18206 5392 18502 5412
rect 18616 4622 18644 6054
rect 18708 5914 18736 6190
rect 18696 5908 18748 5914
rect 18696 5850 18748 5856
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18206 4380 18502 4400
rect 18262 4378 18286 4380
rect 18342 4378 18366 4380
rect 18422 4378 18446 4380
rect 18284 4326 18286 4378
rect 18348 4326 18360 4378
rect 18422 4326 18424 4378
rect 18262 4324 18286 4326
rect 18342 4324 18366 4326
rect 18422 4324 18446 4326
rect 18206 4304 18502 4324
rect 18052 4004 18104 4010
rect 18052 3946 18104 3952
rect 18064 2922 18092 3946
rect 18206 3292 18502 3312
rect 18262 3290 18286 3292
rect 18342 3290 18366 3292
rect 18422 3290 18446 3292
rect 18284 3238 18286 3290
rect 18348 3238 18360 3290
rect 18422 3238 18424 3290
rect 18262 3236 18286 3238
rect 18342 3236 18366 3238
rect 18422 3236 18446 3238
rect 18206 3216 18502 3236
rect 18052 2916 18104 2922
rect 18052 2858 18104 2864
rect 18800 2650 18828 10406
rect 19156 8900 19208 8906
rect 19156 8842 19208 8848
rect 19168 8634 19196 8842
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18892 5710 18920 6190
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18892 5370 18920 5646
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 20732 4826 20760 16646
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20824 5778 20852 16526
rect 20916 12306 20944 17682
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 21008 11354 21036 18022
rect 21192 16590 21220 22374
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 21086 15736 21142 15745
rect 21086 15671 21142 15680
rect 21100 14958 21128 15671
rect 21088 14952 21140 14958
rect 21088 14894 21140 14900
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 20904 11280 20956 11286
rect 20904 11222 20956 11228
rect 20916 10266 20944 11222
rect 21086 10296 21142 10305
rect 20904 10260 20956 10266
rect 21086 10231 21142 10240
rect 20904 10202 20956 10208
rect 21100 10130 21128 10231
rect 21088 10124 21140 10130
rect 21088 10066 21140 10072
rect 21088 8424 21140 8430
rect 21088 8366 21140 8372
rect 20904 8288 20956 8294
rect 21100 8265 21128 8366
rect 20904 8230 20956 8236
rect 21086 8256 21142 8265
rect 20916 7886 20944 8230
rect 21086 8191 21142 8200
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 20904 6724 20956 6730
rect 20904 6666 20956 6672
rect 20916 5914 20944 6666
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 20812 5772 20864 5778
rect 20812 5714 20864 5720
rect 21088 5772 21140 5778
rect 21088 5714 21140 5720
rect 21100 5545 21128 5714
rect 21086 5536 21142 5545
rect 21086 5471 21142 5480
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19444 4282 19472 4626
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19628 4146 19656 4762
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 19616 4140 19668 4146
rect 19616 4082 19668 4088
rect 19628 2990 19656 4082
rect 20180 3942 20208 4218
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 19616 2984 19668 2990
rect 19616 2926 19668 2932
rect 18788 2644 18840 2650
rect 18788 2586 18840 2592
rect 20180 2582 20208 3878
rect 21088 3596 21140 3602
rect 21088 3538 21140 3544
rect 20812 3460 20864 3466
rect 20812 3402 20864 3408
rect 20824 3194 20852 3402
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 21100 2825 21128 3538
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 21086 2816 21142 2825
rect 21086 2751 21142 2760
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 20168 2576 20220 2582
rect 20168 2518 20220 2524
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 18206 2204 18502 2224
rect 18262 2202 18286 2204
rect 18342 2202 18366 2204
rect 18422 2202 18446 2204
rect 18284 2150 18286 2202
rect 18348 2150 18360 2202
rect 18422 2150 18424 2202
rect 18262 2148 18286 2150
rect 18342 2148 18366 2150
rect 18422 2148 18446 2150
rect 18206 2128 18502 2148
rect 18892 800 18920 2450
rect 20720 2372 20772 2378
rect 20720 2314 20772 2320
rect 20732 800 20760 2314
rect 22112 800 22140 2926
rect 478 0 534 800
rect 1858 0 1914 800
rect 3698 0 3754 800
rect 5538 0 5594 800
rect 6918 0 6974 800
rect 8758 0 8814 800
rect 10598 0 10654 800
rect 11978 0 12034 800
rect 13818 0 13874 800
rect 15658 0 15714 800
rect 17038 0 17094 800
rect 18878 0 18934 800
rect 20718 0 20774 800
rect 22098 0 22154 800
<< via2 >>
rect 1490 23160 1546 23216
rect 4406 22874 4462 22876
rect 4486 22874 4542 22876
rect 4566 22874 4622 22876
rect 4646 22874 4702 22876
rect 4406 22822 4432 22874
rect 4432 22822 4462 22874
rect 4486 22822 4496 22874
rect 4496 22822 4542 22874
rect 4566 22822 4612 22874
rect 4612 22822 4622 22874
rect 4646 22822 4676 22874
rect 4676 22822 4702 22874
rect 4406 22820 4462 22822
rect 4486 22820 4542 22822
rect 4566 22820 4622 22822
rect 4646 22820 4702 22822
rect 1398 20440 1454 20496
rect 1398 17740 1454 17776
rect 1398 17720 1400 17740
rect 1400 17720 1452 17740
rect 1452 17720 1454 17740
rect 1398 15680 1454 15736
rect 1490 12980 1546 13016
rect 1490 12960 1492 12980
rect 1492 12960 1544 12980
rect 1544 12960 1546 12980
rect 4406 21786 4462 21788
rect 4486 21786 4542 21788
rect 4566 21786 4622 21788
rect 4646 21786 4702 21788
rect 4406 21734 4432 21786
rect 4432 21734 4462 21786
rect 4486 21734 4496 21786
rect 4496 21734 4542 21786
rect 4566 21734 4612 21786
rect 4612 21734 4622 21786
rect 4646 21734 4676 21786
rect 4676 21734 4702 21786
rect 4406 21732 4462 21734
rect 4486 21732 4542 21734
rect 4566 21732 4622 21734
rect 4646 21732 4702 21734
rect 4406 20698 4462 20700
rect 4486 20698 4542 20700
rect 4566 20698 4622 20700
rect 4646 20698 4702 20700
rect 4406 20646 4432 20698
rect 4432 20646 4462 20698
rect 4486 20646 4496 20698
rect 4496 20646 4542 20698
rect 4566 20646 4612 20698
rect 4612 20646 4622 20698
rect 4646 20646 4676 20698
rect 4676 20646 4702 20698
rect 4406 20644 4462 20646
rect 4486 20644 4542 20646
rect 4566 20644 4622 20646
rect 4646 20644 4702 20646
rect 4406 19610 4462 19612
rect 4486 19610 4542 19612
rect 4566 19610 4622 19612
rect 4646 19610 4702 19612
rect 4406 19558 4432 19610
rect 4432 19558 4462 19610
rect 4486 19558 4496 19610
rect 4496 19558 4542 19610
rect 4566 19558 4612 19610
rect 4612 19558 4622 19610
rect 4646 19558 4676 19610
rect 4676 19558 4702 19610
rect 4406 19556 4462 19558
rect 4486 19556 4542 19558
rect 4566 19556 4622 19558
rect 4646 19556 4702 19558
rect 4406 18522 4462 18524
rect 4486 18522 4542 18524
rect 4566 18522 4622 18524
rect 4646 18522 4702 18524
rect 4406 18470 4432 18522
rect 4432 18470 4462 18522
rect 4486 18470 4496 18522
rect 4496 18470 4542 18522
rect 4566 18470 4612 18522
rect 4612 18470 4622 18522
rect 4646 18470 4676 18522
rect 4676 18470 4702 18522
rect 4406 18468 4462 18470
rect 4486 18468 4542 18470
rect 4566 18468 4622 18470
rect 4646 18468 4702 18470
rect 4406 17434 4462 17436
rect 4486 17434 4542 17436
rect 4566 17434 4622 17436
rect 4646 17434 4702 17436
rect 4406 17382 4432 17434
rect 4432 17382 4462 17434
rect 4486 17382 4496 17434
rect 4496 17382 4542 17434
rect 4566 17382 4612 17434
rect 4612 17382 4622 17434
rect 4646 17382 4676 17434
rect 4676 17382 4702 17434
rect 4406 17380 4462 17382
rect 4486 17380 4542 17382
rect 4566 17380 4622 17382
rect 4646 17380 4702 17382
rect 4406 16346 4462 16348
rect 4486 16346 4542 16348
rect 4566 16346 4622 16348
rect 4646 16346 4702 16348
rect 4406 16294 4432 16346
rect 4432 16294 4462 16346
rect 4486 16294 4496 16346
rect 4496 16294 4542 16346
rect 4566 16294 4612 16346
rect 4612 16294 4622 16346
rect 4646 16294 4676 16346
rect 4676 16294 4702 16346
rect 4406 16292 4462 16294
rect 4486 16292 4542 16294
rect 4566 16292 4622 16294
rect 4646 16292 4702 16294
rect 1490 10240 1546 10296
rect 1398 8200 1454 8256
rect 4406 15258 4462 15260
rect 4486 15258 4542 15260
rect 4566 15258 4622 15260
rect 4646 15258 4702 15260
rect 4406 15206 4432 15258
rect 4432 15206 4462 15258
rect 4486 15206 4496 15258
rect 4496 15206 4542 15258
rect 4566 15206 4612 15258
rect 4612 15206 4622 15258
rect 4646 15206 4676 15258
rect 4676 15206 4702 15258
rect 4406 15204 4462 15206
rect 4486 15204 4542 15206
rect 4566 15204 4622 15206
rect 4646 15204 4702 15206
rect 4406 14170 4462 14172
rect 4486 14170 4542 14172
rect 4566 14170 4622 14172
rect 4646 14170 4702 14172
rect 4406 14118 4432 14170
rect 4432 14118 4462 14170
rect 4486 14118 4496 14170
rect 4496 14118 4542 14170
rect 4566 14118 4612 14170
rect 4612 14118 4622 14170
rect 4646 14118 4676 14170
rect 4676 14118 4702 14170
rect 4406 14116 4462 14118
rect 4486 14116 4542 14118
rect 4566 14116 4622 14118
rect 4646 14116 4702 14118
rect 4406 13082 4462 13084
rect 4486 13082 4542 13084
rect 4566 13082 4622 13084
rect 4646 13082 4702 13084
rect 4406 13030 4432 13082
rect 4432 13030 4462 13082
rect 4486 13030 4496 13082
rect 4496 13030 4542 13082
rect 4566 13030 4612 13082
rect 4612 13030 4622 13082
rect 4646 13030 4676 13082
rect 4676 13030 4702 13082
rect 4406 13028 4462 13030
rect 4486 13028 4542 13030
rect 4566 13028 4622 13030
rect 4646 13028 4702 13030
rect 1490 5516 1492 5536
rect 1492 5516 1544 5536
rect 1544 5516 1546 5536
rect 1490 5480 1546 5516
rect 4406 11994 4462 11996
rect 4486 11994 4542 11996
rect 4566 11994 4622 11996
rect 4646 11994 4702 11996
rect 4406 11942 4432 11994
rect 4432 11942 4462 11994
rect 4486 11942 4496 11994
rect 4496 11942 4542 11994
rect 4566 11942 4612 11994
rect 4612 11942 4622 11994
rect 4646 11942 4676 11994
rect 4676 11942 4702 11994
rect 4406 11940 4462 11942
rect 4486 11940 4542 11942
rect 4566 11940 4622 11942
rect 4646 11940 4702 11942
rect 1398 2760 1454 2816
rect 4406 10906 4462 10908
rect 4486 10906 4542 10908
rect 4566 10906 4622 10908
rect 4646 10906 4702 10908
rect 4406 10854 4432 10906
rect 4432 10854 4462 10906
rect 4486 10854 4496 10906
rect 4496 10854 4542 10906
rect 4566 10854 4612 10906
rect 4612 10854 4622 10906
rect 4646 10854 4676 10906
rect 4676 10854 4702 10906
rect 4406 10852 4462 10854
rect 4486 10852 4542 10854
rect 4566 10852 4622 10854
rect 4646 10852 4702 10854
rect 4406 9818 4462 9820
rect 4486 9818 4542 9820
rect 4566 9818 4622 9820
rect 4646 9818 4702 9820
rect 4406 9766 4432 9818
rect 4432 9766 4462 9818
rect 4486 9766 4496 9818
rect 4496 9766 4542 9818
rect 4566 9766 4612 9818
rect 4612 9766 4622 9818
rect 4646 9766 4676 9818
rect 4676 9766 4702 9818
rect 4406 9764 4462 9766
rect 4486 9764 4542 9766
rect 4566 9764 4622 9766
rect 4646 9764 4702 9766
rect 4406 8730 4462 8732
rect 4486 8730 4542 8732
rect 4566 8730 4622 8732
rect 4646 8730 4702 8732
rect 4406 8678 4432 8730
rect 4432 8678 4462 8730
rect 4486 8678 4496 8730
rect 4496 8678 4542 8730
rect 4566 8678 4612 8730
rect 4612 8678 4622 8730
rect 4646 8678 4676 8730
rect 4676 8678 4702 8730
rect 4406 8676 4462 8678
rect 4486 8676 4542 8678
rect 4566 8676 4622 8678
rect 4646 8676 4702 8678
rect 4406 7642 4462 7644
rect 4486 7642 4542 7644
rect 4566 7642 4622 7644
rect 4646 7642 4702 7644
rect 4406 7590 4432 7642
rect 4432 7590 4462 7642
rect 4486 7590 4496 7642
rect 4496 7590 4542 7642
rect 4566 7590 4612 7642
rect 4612 7590 4622 7642
rect 4646 7590 4676 7642
rect 4676 7590 4702 7642
rect 4406 7588 4462 7590
rect 4486 7588 4542 7590
rect 4566 7588 4622 7590
rect 4646 7588 4702 7590
rect 4406 6554 4462 6556
rect 4486 6554 4542 6556
rect 4566 6554 4622 6556
rect 4646 6554 4702 6556
rect 4406 6502 4432 6554
rect 4432 6502 4462 6554
rect 4486 6502 4496 6554
rect 4496 6502 4542 6554
rect 4566 6502 4612 6554
rect 4612 6502 4622 6554
rect 4646 6502 4676 6554
rect 4676 6502 4702 6554
rect 4406 6500 4462 6502
rect 4486 6500 4542 6502
rect 4566 6500 4622 6502
rect 4646 6500 4702 6502
rect 4406 5466 4462 5468
rect 4486 5466 4542 5468
rect 4566 5466 4622 5468
rect 4646 5466 4702 5468
rect 4406 5414 4432 5466
rect 4432 5414 4462 5466
rect 4486 5414 4496 5466
rect 4496 5414 4542 5466
rect 4566 5414 4612 5466
rect 4612 5414 4622 5466
rect 4646 5414 4676 5466
rect 4676 5414 4702 5466
rect 4406 5412 4462 5414
rect 4486 5412 4542 5414
rect 4566 5412 4622 5414
rect 4646 5412 4702 5414
rect 4406 4378 4462 4380
rect 4486 4378 4542 4380
rect 4566 4378 4622 4380
rect 4646 4378 4702 4380
rect 4406 4326 4432 4378
rect 4432 4326 4462 4378
rect 4486 4326 4496 4378
rect 4496 4326 4542 4378
rect 4566 4326 4612 4378
rect 4612 4326 4622 4378
rect 4646 4326 4676 4378
rect 4676 4326 4702 4378
rect 4406 4324 4462 4326
rect 4486 4324 4542 4326
rect 4566 4324 4622 4326
rect 4646 4324 4702 4326
rect 4406 3290 4462 3292
rect 4486 3290 4542 3292
rect 4566 3290 4622 3292
rect 4646 3290 4702 3292
rect 4406 3238 4432 3290
rect 4432 3238 4462 3290
rect 4486 3238 4496 3290
rect 4496 3238 4542 3290
rect 4566 3238 4612 3290
rect 4612 3238 4622 3290
rect 4646 3238 4676 3290
rect 4676 3238 4702 3290
rect 4406 3236 4462 3238
rect 4486 3236 4542 3238
rect 4566 3236 4622 3238
rect 4646 3236 4702 3238
rect 11306 22874 11362 22876
rect 11386 22874 11442 22876
rect 11466 22874 11522 22876
rect 11546 22874 11602 22876
rect 11306 22822 11332 22874
rect 11332 22822 11362 22874
rect 11386 22822 11396 22874
rect 11396 22822 11442 22874
rect 11466 22822 11512 22874
rect 11512 22822 11522 22874
rect 11546 22822 11576 22874
rect 11576 22822 11602 22874
rect 11306 22820 11362 22822
rect 11386 22820 11442 22822
rect 11466 22820 11522 22822
rect 11546 22820 11602 22822
rect 7856 22330 7912 22332
rect 7936 22330 7992 22332
rect 8016 22330 8072 22332
rect 8096 22330 8152 22332
rect 7856 22278 7882 22330
rect 7882 22278 7912 22330
rect 7936 22278 7946 22330
rect 7946 22278 7992 22330
rect 8016 22278 8062 22330
rect 8062 22278 8072 22330
rect 8096 22278 8126 22330
rect 8126 22278 8152 22330
rect 7856 22276 7912 22278
rect 7936 22276 7992 22278
rect 8016 22276 8072 22278
rect 8096 22276 8152 22278
rect 7856 21242 7912 21244
rect 7936 21242 7992 21244
rect 8016 21242 8072 21244
rect 8096 21242 8152 21244
rect 7856 21190 7882 21242
rect 7882 21190 7912 21242
rect 7936 21190 7946 21242
rect 7946 21190 7992 21242
rect 8016 21190 8062 21242
rect 8062 21190 8072 21242
rect 8096 21190 8126 21242
rect 8126 21190 8152 21242
rect 7856 21188 7912 21190
rect 7936 21188 7992 21190
rect 8016 21188 8072 21190
rect 8096 21188 8152 21190
rect 7856 20154 7912 20156
rect 7936 20154 7992 20156
rect 8016 20154 8072 20156
rect 8096 20154 8152 20156
rect 7856 20102 7882 20154
rect 7882 20102 7912 20154
rect 7936 20102 7946 20154
rect 7946 20102 7992 20154
rect 8016 20102 8062 20154
rect 8062 20102 8072 20154
rect 8096 20102 8126 20154
rect 8126 20102 8152 20154
rect 7856 20100 7912 20102
rect 7936 20100 7992 20102
rect 8016 20100 8072 20102
rect 8096 20100 8152 20102
rect 7194 12552 7250 12608
rect 7856 19066 7912 19068
rect 7936 19066 7992 19068
rect 8016 19066 8072 19068
rect 8096 19066 8152 19068
rect 7856 19014 7882 19066
rect 7882 19014 7912 19066
rect 7936 19014 7946 19066
rect 7946 19014 7992 19066
rect 8016 19014 8062 19066
rect 8062 19014 8072 19066
rect 8096 19014 8126 19066
rect 8126 19014 8152 19066
rect 7856 19012 7912 19014
rect 7936 19012 7992 19014
rect 8016 19012 8072 19014
rect 8096 19012 8152 19014
rect 7856 17978 7912 17980
rect 7936 17978 7992 17980
rect 8016 17978 8072 17980
rect 8096 17978 8152 17980
rect 7856 17926 7882 17978
rect 7882 17926 7912 17978
rect 7936 17926 7946 17978
rect 7946 17926 7992 17978
rect 8016 17926 8062 17978
rect 8062 17926 8072 17978
rect 8096 17926 8126 17978
rect 8126 17926 8152 17978
rect 7856 17924 7912 17926
rect 7936 17924 7992 17926
rect 8016 17924 8072 17926
rect 8096 17924 8152 17926
rect 7856 16890 7912 16892
rect 7936 16890 7992 16892
rect 8016 16890 8072 16892
rect 8096 16890 8152 16892
rect 7856 16838 7882 16890
rect 7882 16838 7912 16890
rect 7936 16838 7946 16890
rect 7946 16838 7992 16890
rect 8016 16838 8062 16890
rect 8062 16838 8072 16890
rect 8096 16838 8126 16890
rect 8126 16838 8152 16890
rect 7856 16836 7912 16838
rect 7936 16836 7992 16838
rect 8016 16836 8072 16838
rect 8096 16836 8152 16838
rect 7856 15802 7912 15804
rect 7936 15802 7992 15804
rect 8016 15802 8072 15804
rect 8096 15802 8152 15804
rect 7856 15750 7882 15802
rect 7882 15750 7912 15802
rect 7936 15750 7946 15802
rect 7946 15750 7992 15802
rect 8016 15750 8062 15802
rect 8062 15750 8072 15802
rect 8096 15750 8126 15802
rect 8126 15750 8152 15802
rect 7856 15748 7912 15750
rect 7936 15748 7992 15750
rect 8016 15748 8072 15750
rect 8096 15748 8152 15750
rect 7856 14714 7912 14716
rect 7936 14714 7992 14716
rect 8016 14714 8072 14716
rect 8096 14714 8152 14716
rect 7856 14662 7882 14714
rect 7882 14662 7912 14714
rect 7936 14662 7946 14714
rect 7946 14662 7992 14714
rect 8016 14662 8062 14714
rect 8062 14662 8072 14714
rect 8096 14662 8126 14714
rect 8126 14662 8152 14714
rect 7856 14660 7912 14662
rect 7936 14660 7992 14662
rect 8016 14660 8072 14662
rect 8096 14660 8152 14662
rect 7856 13626 7912 13628
rect 7936 13626 7992 13628
rect 8016 13626 8072 13628
rect 8096 13626 8152 13628
rect 7856 13574 7882 13626
rect 7882 13574 7912 13626
rect 7936 13574 7946 13626
rect 7946 13574 7992 13626
rect 8016 13574 8062 13626
rect 8062 13574 8072 13626
rect 8096 13574 8126 13626
rect 8126 13574 8152 13626
rect 7856 13572 7912 13574
rect 7936 13572 7992 13574
rect 8016 13572 8072 13574
rect 8096 13572 8152 13574
rect 7562 12552 7618 12608
rect 7856 12538 7912 12540
rect 7936 12538 7992 12540
rect 8016 12538 8072 12540
rect 8096 12538 8152 12540
rect 7856 12486 7882 12538
rect 7882 12486 7912 12538
rect 7936 12486 7946 12538
rect 7946 12486 7992 12538
rect 8016 12486 8062 12538
rect 8062 12486 8072 12538
rect 8096 12486 8126 12538
rect 8126 12486 8152 12538
rect 7856 12484 7912 12486
rect 7936 12484 7992 12486
rect 8016 12484 8072 12486
rect 8096 12484 8152 12486
rect 7856 11450 7912 11452
rect 7936 11450 7992 11452
rect 8016 11450 8072 11452
rect 8096 11450 8152 11452
rect 7856 11398 7882 11450
rect 7882 11398 7912 11450
rect 7936 11398 7946 11450
rect 7946 11398 7992 11450
rect 8016 11398 8062 11450
rect 8062 11398 8072 11450
rect 8096 11398 8126 11450
rect 8126 11398 8152 11450
rect 7856 11396 7912 11398
rect 7936 11396 7992 11398
rect 8016 11396 8072 11398
rect 8096 11396 8152 11398
rect 7856 10362 7912 10364
rect 7936 10362 7992 10364
rect 8016 10362 8072 10364
rect 8096 10362 8152 10364
rect 7856 10310 7882 10362
rect 7882 10310 7912 10362
rect 7936 10310 7946 10362
rect 7946 10310 7992 10362
rect 8016 10310 8062 10362
rect 8062 10310 8072 10362
rect 8096 10310 8126 10362
rect 8126 10310 8152 10362
rect 7856 10308 7912 10310
rect 7936 10308 7992 10310
rect 8016 10308 8072 10310
rect 8096 10308 8152 10310
rect 7856 9274 7912 9276
rect 7936 9274 7992 9276
rect 8016 9274 8072 9276
rect 8096 9274 8152 9276
rect 7856 9222 7882 9274
rect 7882 9222 7912 9274
rect 7936 9222 7946 9274
rect 7946 9222 7992 9274
rect 8016 9222 8062 9274
rect 8062 9222 8072 9274
rect 8096 9222 8126 9274
rect 8126 9222 8152 9274
rect 7856 9220 7912 9222
rect 7936 9220 7992 9222
rect 8016 9220 8072 9222
rect 8096 9220 8152 9222
rect 7856 8186 7912 8188
rect 7936 8186 7992 8188
rect 8016 8186 8072 8188
rect 8096 8186 8152 8188
rect 7856 8134 7882 8186
rect 7882 8134 7912 8186
rect 7936 8134 7946 8186
rect 7946 8134 7992 8186
rect 8016 8134 8062 8186
rect 8062 8134 8072 8186
rect 8096 8134 8126 8186
rect 8126 8134 8152 8186
rect 7856 8132 7912 8134
rect 7936 8132 7992 8134
rect 8016 8132 8072 8134
rect 8096 8132 8152 8134
rect 7856 7098 7912 7100
rect 7936 7098 7992 7100
rect 8016 7098 8072 7100
rect 8096 7098 8152 7100
rect 7856 7046 7882 7098
rect 7882 7046 7912 7098
rect 7936 7046 7946 7098
rect 7946 7046 7992 7098
rect 8016 7046 8062 7098
rect 8062 7046 8072 7098
rect 8096 7046 8126 7098
rect 8126 7046 8152 7098
rect 7856 7044 7912 7046
rect 7936 7044 7992 7046
rect 8016 7044 8072 7046
rect 8096 7044 8152 7046
rect 7856 6010 7912 6012
rect 7936 6010 7992 6012
rect 8016 6010 8072 6012
rect 8096 6010 8152 6012
rect 7856 5958 7882 6010
rect 7882 5958 7912 6010
rect 7936 5958 7946 6010
rect 7946 5958 7992 6010
rect 8016 5958 8062 6010
rect 8062 5958 8072 6010
rect 8096 5958 8126 6010
rect 8126 5958 8152 6010
rect 7856 5956 7912 5958
rect 7936 5956 7992 5958
rect 8016 5956 8072 5958
rect 8096 5956 8152 5958
rect 7856 4922 7912 4924
rect 7936 4922 7992 4924
rect 8016 4922 8072 4924
rect 8096 4922 8152 4924
rect 7856 4870 7882 4922
rect 7882 4870 7912 4922
rect 7936 4870 7946 4922
rect 7946 4870 7992 4922
rect 8016 4870 8062 4922
rect 8062 4870 8072 4922
rect 8096 4870 8126 4922
rect 8126 4870 8152 4922
rect 7856 4868 7912 4870
rect 7936 4868 7992 4870
rect 8016 4868 8072 4870
rect 8096 4868 8152 4870
rect 7856 3834 7912 3836
rect 7936 3834 7992 3836
rect 8016 3834 8072 3836
rect 8096 3834 8152 3836
rect 7856 3782 7882 3834
rect 7882 3782 7912 3834
rect 7936 3782 7946 3834
rect 7946 3782 7992 3834
rect 8016 3782 8062 3834
rect 8062 3782 8072 3834
rect 8096 3782 8126 3834
rect 8126 3782 8152 3834
rect 7856 3780 7912 3782
rect 7936 3780 7992 3782
rect 8016 3780 8072 3782
rect 8096 3780 8152 3782
rect 7856 2746 7912 2748
rect 7936 2746 7992 2748
rect 8016 2746 8072 2748
rect 8096 2746 8152 2748
rect 7856 2694 7882 2746
rect 7882 2694 7912 2746
rect 7936 2694 7946 2746
rect 7946 2694 7992 2746
rect 8016 2694 8062 2746
rect 8062 2694 8072 2746
rect 8096 2694 8126 2746
rect 8126 2694 8152 2746
rect 7856 2692 7912 2694
rect 7936 2692 7992 2694
rect 8016 2692 8072 2694
rect 8096 2692 8152 2694
rect 18206 22874 18262 22876
rect 18286 22874 18342 22876
rect 18366 22874 18422 22876
rect 18446 22874 18502 22876
rect 18206 22822 18232 22874
rect 18232 22822 18262 22874
rect 18286 22822 18296 22874
rect 18296 22822 18342 22874
rect 18366 22822 18412 22874
rect 18412 22822 18422 22874
rect 18446 22822 18476 22874
rect 18476 22822 18502 22874
rect 18206 22820 18262 22822
rect 18286 22820 18342 22822
rect 18366 22820 18422 22822
rect 18446 22820 18502 22822
rect 21086 23160 21142 23216
rect 11306 21786 11362 21788
rect 11386 21786 11442 21788
rect 11466 21786 11522 21788
rect 11546 21786 11602 21788
rect 11306 21734 11332 21786
rect 11332 21734 11362 21786
rect 11386 21734 11396 21786
rect 11396 21734 11442 21786
rect 11466 21734 11512 21786
rect 11512 21734 11522 21786
rect 11546 21734 11576 21786
rect 11576 21734 11602 21786
rect 11306 21732 11362 21734
rect 11386 21732 11442 21734
rect 11466 21732 11522 21734
rect 11546 21732 11602 21734
rect 11306 20698 11362 20700
rect 11386 20698 11442 20700
rect 11466 20698 11522 20700
rect 11546 20698 11602 20700
rect 11306 20646 11332 20698
rect 11332 20646 11362 20698
rect 11386 20646 11396 20698
rect 11396 20646 11442 20698
rect 11466 20646 11512 20698
rect 11512 20646 11522 20698
rect 11546 20646 11576 20698
rect 11576 20646 11602 20698
rect 11306 20644 11362 20646
rect 11386 20644 11442 20646
rect 11466 20644 11522 20646
rect 11546 20644 11602 20646
rect 11306 19610 11362 19612
rect 11386 19610 11442 19612
rect 11466 19610 11522 19612
rect 11546 19610 11602 19612
rect 11306 19558 11332 19610
rect 11332 19558 11362 19610
rect 11386 19558 11396 19610
rect 11396 19558 11442 19610
rect 11466 19558 11512 19610
rect 11512 19558 11522 19610
rect 11546 19558 11576 19610
rect 11576 19558 11602 19610
rect 11306 19556 11362 19558
rect 11386 19556 11442 19558
rect 11466 19556 11522 19558
rect 11546 19556 11602 19558
rect 11306 18522 11362 18524
rect 11386 18522 11442 18524
rect 11466 18522 11522 18524
rect 11546 18522 11602 18524
rect 11306 18470 11332 18522
rect 11332 18470 11362 18522
rect 11386 18470 11396 18522
rect 11396 18470 11442 18522
rect 11466 18470 11512 18522
rect 11512 18470 11522 18522
rect 11546 18470 11576 18522
rect 11576 18470 11602 18522
rect 11306 18468 11362 18470
rect 11386 18468 11442 18470
rect 11466 18468 11522 18470
rect 11546 18468 11602 18470
rect 11306 17434 11362 17436
rect 11386 17434 11442 17436
rect 11466 17434 11522 17436
rect 11546 17434 11602 17436
rect 11306 17382 11332 17434
rect 11332 17382 11362 17434
rect 11386 17382 11396 17434
rect 11396 17382 11442 17434
rect 11466 17382 11512 17434
rect 11512 17382 11522 17434
rect 11546 17382 11576 17434
rect 11576 17382 11602 17434
rect 11306 17380 11362 17382
rect 11386 17380 11442 17382
rect 11466 17380 11522 17382
rect 11546 17380 11602 17382
rect 11306 16346 11362 16348
rect 11386 16346 11442 16348
rect 11466 16346 11522 16348
rect 11546 16346 11602 16348
rect 11306 16294 11332 16346
rect 11332 16294 11362 16346
rect 11386 16294 11396 16346
rect 11396 16294 11442 16346
rect 11466 16294 11512 16346
rect 11512 16294 11522 16346
rect 11546 16294 11576 16346
rect 11576 16294 11602 16346
rect 11306 16292 11362 16294
rect 11386 16292 11442 16294
rect 11466 16292 11522 16294
rect 11546 16292 11602 16294
rect 11306 15258 11362 15260
rect 11386 15258 11442 15260
rect 11466 15258 11522 15260
rect 11546 15258 11602 15260
rect 11306 15206 11332 15258
rect 11332 15206 11362 15258
rect 11386 15206 11396 15258
rect 11396 15206 11442 15258
rect 11466 15206 11512 15258
rect 11512 15206 11522 15258
rect 11546 15206 11576 15258
rect 11576 15206 11602 15258
rect 11306 15204 11362 15206
rect 11386 15204 11442 15206
rect 11466 15204 11522 15206
rect 11546 15204 11602 15206
rect 11306 14170 11362 14172
rect 11386 14170 11442 14172
rect 11466 14170 11522 14172
rect 11546 14170 11602 14172
rect 11306 14118 11332 14170
rect 11332 14118 11362 14170
rect 11386 14118 11396 14170
rect 11396 14118 11442 14170
rect 11466 14118 11512 14170
rect 11512 14118 11522 14170
rect 11546 14118 11576 14170
rect 11576 14118 11602 14170
rect 11306 14116 11362 14118
rect 11386 14116 11442 14118
rect 11466 14116 11522 14118
rect 11546 14116 11602 14118
rect 11306 13082 11362 13084
rect 11386 13082 11442 13084
rect 11466 13082 11522 13084
rect 11546 13082 11602 13084
rect 11306 13030 11332 13082
rect 11332 13030 11362 13082
rect 11386 13030 11396 13082
rect 11396 13030 11442 13082
rect 11466 13030 11512 13082
rect 11512 13030 11522 13082
rect 11546 13030 11576 13082
rect 11576 13030 11602 13082
rect 11306 13028 11362 13030
rect 11386 13028 11442 13030
rect 11466 13028 11522 13030
rect 11546 13028 11602 13030
rect 11306 11994 11362 11996
rect 11386 11994 11442 11996
rect 11466 11994 11522 11996
rect 11546 11994 11602 11996
rect 11306 11942 11332 11994
rect 11332 11942 11362 11994
rect 11386 11942 11396 11994
rect 11396 11942 11442 11994
rect 11466 11942 11512 11994
rect 11512 11942 11522 11994
rect 11546 11942 11576 11994
rect 11576 11942 11602 11994
rect 11306 11940 11362 11942
rect 11386 11940 11442 11942
rect 11466 11940 11522 11942
rect 11546 11940 11602 11942
rect 11306 10906 11362 10908
rect 11386 10906 11442 10908
rect 11466 10906 11522 10908
rect 11546 10906 11602 10908
rect 11306 10854 11332 10906
rect 11332 10854 11362 10906
rect 11386 10854 11396 10906
rect 11396 10854 11442 10906
rect 11466 10854 11512 10906
rect 11512 10854 11522 10906
rect 11546 10854 11576 10906
rect 11576 10854 11602 10906
rect 11306 10852 11362 10854
rect 11386 10852 11442 10854
rect 11466 10852 11522 10854
rect 11546 10852 11602 10854
rect 11306 9818 11362 9820
rect 11386 9818 11442 9820
rect 11466 9818 11522 9820
rect 11546 9818 11602 9820
rect 11306 9766 11332 9818
rect 11332 9766 11362 9818
rect 11386 9766 11396 9818
rect 11396 9766 11442 9818
rect 11466 9766 11512 9818
rect 11512 9766 11522 9818
rect 11546 9766 11576 9818
rect 11576 9766 11602 9818
rect 11306 9764 11362 9766
rect 11386 9764 11442 9766
rect 11466 9764 11522 9766
rect 11546 9764 11602 9766
rect 11306 8730 11362 8732
rect 11386 8730 11442 8732
rect 11466 8730 11522 8732
rect 11546 8730 11602 8732
rect 11306 8678 11332 8730
rect 11332 8678 11362 8730
rect 11386 8678 11396 8730
rect 11396 8678 11442 8730
rect 11466 8678 11512 8730
rect 11512 8678 11522 8730
rect 11546 8678 11576 8730
rect 11576 8678 11602 8730
rect 11306 8676 11362 8678
rect 11386 8676 11442 8678
rect 11466 8676 11522 8678
rect 11546 8676 11602 8678
rect 11306 7642 11362 7644
rect 11386 7642 11442 7644
rect 11466 7642 11522 7644
rect 11546 7642 11602 7644
rect 11306 7590 11332 7642
rect 11332 7590 11362 7642
rect 11386 7590 11396 7642
rect 11396 7590 11442 7642
rect 11466 7590 11512 7642
rect 11512 7590 11522 7642
rect 11546 7590 11576 7642
rect 11576 7590 11602 7642
rect 11306 7588 11362 7590
rect 11386 7588 11442 7590
rect 11466 7588 11522 7590
rect 11546 7588 11602 7590
rect 11306 6554 11362 6556
rect 11386 6554 11442 6556
rect 11466 6554 11522 6556
rect 11546 6554 11602 6556
rect 11306 6502 11332 6554
rect 11332 6502 11362 6554
rect 11386 6502 11396 6554
rect 11396 6502 11442 6554
rect 11466 6502 11512 6554
rect 11512 6502 11522 6554
rect 11546 6502 11576 6554
rect 11576 6502 11602 6554
rect 11306 6500 11362 6502
rect 11386 6500 11442 6502
rect 11466 6500 11522 6502
rect 11546 6500 11602 6502
rect 11306 5466 11362 5468
rect 11386 5466 11442 5468
rect 11466 5466 11522 5468
rect 11546 5466 11602 5468
rect 11306 5414 11332 5466
rect 11332 5414 11362 5466
rect 11386 5414 11396 5466
rect 11396 5414 11442 5466
rect 11466 5414 11512 5466
rect 11512 5414 11522 5466
rect 11546 5414 11576 5466
rect 11576 5414 11602 5466
rect 11306 5412 11362 5414
rect 11386 5412 11442 5414
rect 11466 5412 11522 5414
rect 11546 5412 11602 5414
rect 11306 4378 11362 4380
rect 11386 4378 11442 4380
rect 11466 4378 11522 4380
rect 11546 4378 11602 4380
rect 11306 4326 11332 4378
rect 11332 4326 11362 4378
rect 11386 4326 11396 4378
rect 11396 4326 11442 4378
rect 11466 4326 11512 4378
rect 11512 4326 11522 4378
rect 11546 4326 11576 4378
rect 11576 4326 11602 4378
rect 11306 4324 11362 4326
rect 11386 4324 11442 4326
rect 11466 4324 11522 4326
rect 11546 4324 11602 4326
rect 11306 3290 11362 3292
rect 11386 3290 11442 3292
rect 11466 3290 11522 3292
rect 11546 3290 11602 3292
rect 11306 3238 11332 3290
rect 11332 3238 11362 3290
rect 11386 3238 11396 3290
rect 11396 3238 11442 3290
rect 11466 3238 11512 3290
rect 11512 3238 11522 3290
rect 11546 3238 11576 3290
rect 11576 3238 11602 3290
rect 11306 3236 11362 3238
rect 11386 3236 11442 3238
rect 11466 3236 11522 3238
rect 11546 3236 11602 3238
rect 4406 2202 4462 2204
rect 4486 2202 4542 2204
rect 4566 2202 4622 2204
rect 4646 2202 4702 2204
rect 4406 2150 4432 2202
rect 4432 2150 4462 2202
rect 4486 2150 4496 2202
rect 4496 2150 4542 2202
rect 4566 2150 4612 2202
rect 4612 2150 4622 2202
rect 4646 2150 4676 2202
rect 4676 2150 4702 2202
rect 4406 2148 4462 2150
rect 4486 2148 4542 2150
rect 4566 2148 4622 2150
rect 4646 2148 4702 2150
rect 11306 2202 11362 2204
rect 11386 2202 11442 2204
rect 11466 2202 11522 2204
rect 11546 2202 11602 2204
rect 11306 2150 11332 2202
rect 11332 2150 11362 2202
rect 11386 2150 11396 2202
rect 11396 2150 11442 2202
rect 11466 2150 11512 2202
rect 11512 2150 11522 2202
rect 11546 2150 11576 2202
rect 11576 2150 11602 2202
rect 11306 2148 11362 2150
rect 11386 2148 11442 2150
rect 11466 2148 11522 2150
rect 11546 2148 11602 2150
rect 14756 22330 14812 22332
rect 14836 22330 14892 22332
rect 14916 22330 14972 22332
rect 14996 22330 15052 22332
rect 14756 22278 14782 22330
rect 14782 22278 14812 22330
rect 14836 22278 14846 22330
rect 14846 22278 14892 22330
rect 14916 22278 14962 22330
rect 14962 22278 14972 22330
rect 14996 22278 15026 22330
rect 15026 22278 15052 22330
rect 14756 22276 14812 22278
rect 14836 22276 14892 22278
rect 14916 22276 14972 22278
rect 14996 22276 15052 22278
rect 14756 21242 14812 21244
rect 14836 21242 14892 21244
rect 14916 21242 14972 21244
rect 14996 21242 15052 21244
rect 14756 21190 14782 21242
rect 14782 21190 14812 21242
rect 14836 21190 14846 21242
rect 14846 21190 14892 21242
rect 14916 21190 14962 21242
rect 14962 21190 14972 21242
rect 14996 21190 15026 21242
rect 15026 21190 15052 21242
rect 14756 21188 14812 21190
rect 14836 21188 14892 21190
rect 14916 21188 14972 21190
rect 14996 21188 15052 21190
rect 14756 20154 14812 20156
rect 14836 20154 14892 20156
rect 14916 20154 14972 20156
rect 14996 20154 15052 20156
rect 14756 20102 14782 20154
rect 14782 20102 14812 20154
rect 14836 20102 14846 20154
rect 14846 20102 14892 20154
rect 14916 20102 14962 20154
rect 14962 20102 14972 20154
rect 14996 20102 15026 20154
rect 15026 20102 15052 20154
rect 14756 20100 14812 20102
rect 14836 20100 14892 20102
rect 14916 20100 14972 20102
rect 14996 20100 15052 20102
rect 14756 19066 14812 19068
rect 14836 19066 14892 19068
rect 14916 19066 14972 19068
rect 14996 19066 15052 19068
rect 14756 19014 14782 19066
rect 14782 19014 14812 19066
rect 14836 19014 14846 19066
rect 14846 19014 14892 19066
rect 14916 19014 14962 19066
rect 14962 19014 14972 19066
rect 14996 19014 15026 19066
rect 15026 19014 15052 19066
rect 14756 19012 14812 19014
rect 14836 19012 14892 19014
rect 14916 19012 14972 19014
rect 14996 19012 15052 19014
rect 14756 17978 14812 17980
rect 14836 17978 14892 17980
rect 14916 17978 14972 17980
rect 14996 17978 15052 17980
rect 14756 17926 14782 17978
rect 14782 17926 14812 17978
rect 14836 17926 14846 17978
rect 14846 17926 14892 17978
rect 14916 17926 14962 17978
rect 14962 17926 14972 17978
rect 14996 17926 15026 17978
rect 15026 17926 15052 17978
rect 14756 17924 14812 17926
rect 14836 17924 14892 17926
rect 14916 17924 14972 17926
rect 14996 17924 15052 17926
rect 14756 16890 14812 16892
rect 14836 16890 14892 16892
rect 14916 16890 14972 16892
rect 14996 16890 15052 16892
rect 14756 16838 14782 16890
rect 14782 16838 14812 16890
rect 14836 16838 14846 16890
rect 14846 16838 14892 16890
rect 14916 16838 14962 16890
rect 14962 16838 14972 16890
rect 14996 16838 15026 16890
rect 15026 16838 15052 16890
rect 14756 16836 14812 16838
rect 14836 16836 14892 16838
rect 14916 16836 14972 16838
rect 14996 16836 15052 16838
rect 14756 15802 14812 15804
rect 14836 15802 14892 15804
rect 14916 15802 14972 15804
rect 14996 15802 15052 15804
rect 14756 15750 14782 15802
rect 14782 15750 14812 15802
rect 14836 15750 14846 15802
rect 14846 15750 14892 15802
rect 14916 15750 14962 15802
rect 14962 15750 14972 15802
rect 14996 15750 15026 15802
rect 15026 15750 15052 15802
rect 14756 15748 14812 15750
rect 14836 15748 14892 15750
rect 14916 15748 14972 15750
rect 14996 15748 15052 15750
rect 14756 14714 14812 14716
rect 14836 14714 14892 14716
rect 14916 14714 14972 14716
rect 14996 14714 15052 14716
rect 14756 14662 14782 14714
rect 14782 14662 14812 14714
rect 14836 14662 14846 14714
rect 14846 14662 14892 14714
rect 14916 14662 14962 14714
rect 14962 14662 14972 14714
rect 14996 14662 15026 14714
rect 15026 14662 15052 14714
rect 14756 14660 14812 14662
rect 14836 14660 14892 14662
rect 14916 14660 14972 14662
rect 14996 14660 15052 14662
rect 14756 13626 14812 13628
rect 14836 13626 14892 13628
rect 14916 13626 14972 13628
rect 14996 13626 15052 13628
rect 14756 13574 14782 13626
rect 14782 13574 14812 13626
rect 14836 13574 14846 13626
rect 14846 13574 14892 13626
rect 14916 13574 14962 13626
rect 14962 13574 14972 13626
rect 14996 13574 15026 13626
rect 15026 13574 15052 13626
rect 14756 13572 14812 13574
rect 14836 13572 14892 13574
rect 14916 13572 14972 13574
rect 14996 13572 15052 13574
rect 14756 12538 14812 12540
rect 14836 12538 14892 12540
rect 14916 12538 14972 12540
rect 14996 12538 15052 12540
rect 14756 12486 14782 12538
rect 14782 12486 14812 12538
rect 14836 12486 14846 12538
rect 14846 12486 14892 12538
rect 14916 12486 14962 12538
rect 14962 12486 14972 12538
rect 14996 12486 15026 12538
rect 15026 12486 15052 12538
rect 14756 12484 14812 12486
rect 14836 12484 14892 12486
rect 14916 12484 14972 12486
rect 14996 12484 15052 12486
rect 14756 11450 14812 11452
rect 14836 11450 14892 11452
rect 14916 11450 14972 11452
rect 14996 11450 15052 11452
rect 14756 11398 14782 11450
rect 14782 11398 14812 11450
rect 14836 11398 14846 11450
rect 14846 11398 14892 11450
rect 14916 11398 14962 11450
rect 14962 11398 14972 11450
rect 14996 11398 15026 11450
rect 15026 11398 15052 11450
rect 14756 11396 14812 11398
rect 14836 11396 14892 11398
rect 14916 11396 14972 11398
rect 14996 11396 15052 11398
rect 14756 10362 14812 10364
rect 14836 10362 14892 10364
rect 14916 10362 14972 10364
rect 14996 10362 15052 10364
rect 14756 10310 14782 10362
rect 14782 10310 14812 10362
rect 14836 10310 14846 10362
rect 14846 10310 14892 10362
rect 14916 10310 14962 10362
rect 14962 10310 14972 10362
rect 14996 10310 15026 10362
rect 15026 10310 15052 10362
rect 14756 10308 14812 10310
rect 14836 10308 14892 10310
rect 14916 10308 14972 10310
rect 14996 10308 15052 10310
rect 14756 9274 14812 9276
rect 14836 9274 14892 9276
rect 14916 9274 14972 9276
rect 14996 9274 15052 9276
rect 14756 9222 14782 9274
rect 14782 9222 14812 9274
rect 14836 9222 14846 9274
rect 14846 9222 14892 9274
rect 14916 9222 14962 9274
rect 14962 9222 14972 9274
rect 14996 9222 15026 9274
rect 15026 9222 15052 9274
rect 14756 9220 14812 9222
rect 14836 9220 14892 9222
rect 14916 9220 14972 9222
rect 14996 9220 15052 9222
rect 18206 21786 18262 21788
rect 18286 21786 18342 21788
rect 18366 21786 18422 21788
rect 18446 21786 18502 21788
rect 18206 21734 18232 21786
rect 18232 21734 18262 21786
rect 18286 21734 18296 21786
rect 18296 21734 18342 21786
rect 18366 21734 18412 21786
rect 18412 21734 18422 21786
rect 18446 21734 18476 21786
rect 18476 21734 18502 21786
rect 18206 21732 18262 21734
rect 18286 21732 18342 21734
rect 18366 21732 18422 21734
rect 18446 21732 18502 21734
rect 18206 20698 18262 20700
rect 18286 20698 18342 20700
rect 18366 20698 18422 20700
rect 18446 20698 18502 20700
rect 18206 20646 18232 20698
rect 18232 20646 18262 20698
rect 18286 20646 18296 20698
rect 18296 20646 18342 20698
rect 18366 20646 18412 20698
rect 18412 20646 18422 20698
rect 18446 20646 18476 20698
rect 18476 20646 18502 20698
rect 18206 20644 18262 20646
rect 18286 20644 18342 20646
rect 18366 20644 18422 20646
rect 18446 20644 18502 20646
rect 18206 19610 18262 19612
rect 18286 19610 18342 19612
rect 18366 19610 18422 19612
rect 18446 19610 18502 19612
rect 18206 19558 18232 19610
rect 18232 19558 18262 19610
rect 18286 19558 18296 19610
rect 18296 19558 18342 19610
rect 18366 19558 18412 19610
rect 18412 19558 18422 19610
rect 18446 19558 18476 19610
rect 18476 19558 18502 19610
rect 18206 19556 18262 19558
rect 18286 19556 18342 19558
rect 18366 19556 18422 19558
rect 18446 19556 18502 19558
rect 20626 20440 20682 20496
rect 18206 18522 18262 18524
rect 18286 18522 18342 18524
rect 18366 18522 18422 18524
rect 18446 18522 18502 18524
rect 18206 18470 18232 18522
rect 18232 18470 18262 18522
rect 18286 18470 18296 18522
rect 18296 18470 18342 18522
rect 18366 18470 18412 18522
rect 18412 18470 18422 18522
rect 18446 18470 18476 18522
rect 18476 18470 18502 18522
rect 18206 18468 18262 18470
rect 18286 18468 18342 18470
rect 18366 18468 18422 18470
rect 18446 18468 18502 18470
rect 18206 17434 18262 17436
rect 18286 17434 18342 17436
rect 18366 17434 18422 17436
rect 18446 17434 18502 17436
rect 18206 17382 18232 17434
rect 18232 17382 18262 17434
rect 18286 17382 18296 17434
rect 18296 17382 18342 17434
rect 18366 17382 18412 17434
rect 18412 17382 18422 17434
rect 18446 17382 18476 17434
rect 18476 17382 18502 17434
rect 18206 17380 18262 17382
rect 18286 17380 18342 17382
rect 18366 17380 18422 17382
rect 18446 17380 18502 17382
rect 18206 16346 18262 16348
rect 18286 16346 18342 16348
rect 18366 16346 18422 16348
rect 18446 16346 18502 16348
rect 18206 16294 18232 16346
rect 18232 16294 18262 16346
rect 18286 16294 18296 16346
rect 18296 16294 18342 16346
rect 18366 16294 18412 16346
rect 18412 16294 18422 16346
rect 18446 16294 18476 16346
rect 18476 16294 18502 16346
rect 18206 16292 18262 16294
rect 18286 16292 18342 16294
rect 18366 16292 18422 16294
rect 18446 16292 18502 16294
rect 18206 15258 18262 15260
rect 18286 15258 18342 15260
rect 18366 15258 18422 15260
rect 18446 15258 18502 15260
rect 18206 15206 18232 15258
rect 18232 15206 18262 15258
rect 18286 15206 18296 15258
rect 18296 15206 18342 15258
rect 18366 15206 18412 15258
rect 18412 15206 18422 15258
rect 18446 15206 18476 15258
rect 18476 15206 18502 15258
rect 18206 15204 18262 15206
rect 18286 15204 18342 15206
rect 18366 15204 18422 15206
rect 18446 15204 18502 15206
rect 18206 14170 18262 14172
rect 18286 14170 18342 14172
rect 18366 14170 18422 14172
rect 18446 14170 18502 14172
rect 18206 14118 18232 14170
rect 18232 14118 18262 14170
rect 18286 14118 18296 14170
rect 18296 14118 18342 14170
rect 18366 14118 18412 14170
rect 18412 14118 18422 14170
rect 18446 14118 18476 14170
rect 18476 14118 18502 14170
rect 18206 14116 18262 14118
rect 18286 14116 18342 14118
rect 18366 14116 18422 14118
rect 18446 14116 18502 14118
rect 18206 13082 18262 13084
rect 18286 13082 18342 13084
rect 18366 13082 18422 13084
rect 18446 13082 18502 13084
rect 18206 13030 18232 13082
rect 18232 13030 18262 13082
rect 18286 13030 18296 13082
rect 18296 13030 18342 13082
rect 18366 13030 18412 13082
rect 18412 13030 18422 13082
rect 18446 13030 18476 13082
rect 18476 13030 18502 13082
rect 18206 13028 18262 13030
rect 18286 13028 18342 13030
rect 18366 13028 18422 13030
rect 18446 13028 18502 13030
rect 20626 17720 20682 17776
rect 18206 11994 18262 11996
rect 18286 11994 18342 11996
rect 18366 11994 18422 11996
rect 18446 11994 18502 11996
rect 18206 11942 18232 11994
rect 18232 11942 18262 11994
rect 18286 11942 18296 11994
rect 18296 11942 18342 11994
rect 18366 11942 18412 11994
rect 18412 11942 18422 11994
rect 18446 11942 18476 11994
rect 18476 11942 18502 11994
rect 18206 11940 18262 11942
rect 18286 11940 18342 11942
rect 18366 11940 18422 11942
rect 18446 11940 18502 11942
rect 14756 8186 14812 8188
rect 14836 8186 14892 8188
rect 14916 8186 14972 8188
rect 14996 8186 15052 8188
rect 14756 8134 14782 8186
rect 14782 8134 14812 8186
rect 14836 8134 14846 8186
rect 14846 8134 14892 8186
rect 14916 8134 14962 8186
rect 14962 8134 14972 8186
rect 14996 8134 15026 8186
rect 15026 8134 15052 8186
rect 14756 8132 14812 8134
rect 14836 8132 14892 8134
rect 14916 8132 14972 8134
rect 14996 8132 15052 8134
rect 14756 7098 14812 7100
rect 14836 7098 14892 7100
rect 14916 7098 14972 7100
rect 14996 7098 15052 7100
rect 14756 7046 14782 7098
rect 14782 7046 14812 7098
rect 14836 7046 14846 7098
rect 14846 7046 14892 7098
rect 14916 7046 14962 7098
rect 14962 7046 14972 7098
rect 14996 7046 15026 7098
rect 15026 7046 15052 7098
rect 14756 7044 14812 7046
rect 14836 7044 14892 7046
rect 14916 7044 14972 7046
rect 14996 7044 15052 7046
rect 18206 10906 18262 10908
rect 18286 10906 18342 10908
rect 18366 10906 18422 10908
rect 18446 10906 18502 10908
rect 18206 10854 18232 10906
rect 18232 10854 18262 10906
rect 18286 10854 18296 10906
rect 18296 10854 18342 10906
rect 18366 10854 18412 10906
rect 18412 10854 18422 10906
rect 18446 10854 18476 10906
rect 18476 10854 18502 10906
rect 18206 10852 18262 10854
rect 18286 10852 18342 10854
rect 18366 10852 18422 10854
rect 18446 10852 18502 10854
rect 20626 12960 20682 13016
rect 18206 9818 18262 9820
rect 18286 9818 18342 9820
rect 18366 9818 18422 9820
rect 18446 9818 18502 9820
rect 18206 9766 18232 9818
rect 18232 9766 18262 9818
rect 18286 9766 18296 9818
rect 18296 9766 18342 9818
rect 18366 9766 18412 9818
rect 18412 9766 18422 9818
rect 18446 9766 18476 9818
rect 18476 9766 18502 9818
rect 18206 9764 18262 9766
rect 18286 9764 18342 9766
rect 18366 9764 18422 9766
rect 18446 9764 18502 9766
rect 18206 8730 18262 8732
rect 18286 8730 18342 8732
rect 18366 8730 18422 8732
rect 18446 8730 18502 8732
rect 18206 8678 18232 8730
rect 18232 8678 18262 8730
rect 18286 8678 18296 8730
rect 18296 8678 18342 8730
rect 18366 8678 18412 8730
rect 18412 8678 18422 8730
rect 18446 8678 18476 8730
rect 18476 8678 18502 8730
rect 18206 8676 18262 8678
rect 18286 8676 18342 8678
rect 18366 8676 18422 8678
rect 18446 8676 18502 8678
rect 18206 7642 18262 7644
rect 18286 7642 18342 7644
rect 18366 7642 18422 7644
rect 18446 7642 18502 7644
rect 18206 7590 18232 7642
rect 18232 7590 18262 7642
rect 18286 7590 18296 7642
rect 18296 7590 18342 7642
rect 18366 7590 18412 7642
rect 18412 7590 18422 7642
rect 18446 7590 18476 7642
rect 18476 7590 18502 7642
rect 18206 7588 18262 7590
rect 18286 7588 18342 7590
rect 18366 7588 18422 7590
rect 18446 7588 18502 7590
rect 14756 6010 14812 6012
rect 14836 6010 14892 6012
rect 14916 6010 14972 6012
rect 14996 6010 15052 6012
rect 14756 5958 14782 6010
rect 14782 5958 14812 6010
rect 14836 5958 14846 6010
rect 14846 5958 14892 6010
rect 14916 5958 14962 6010
rect 14962 5958 14972 6010
rect 14996 5958 15026 6010
rect 15026 5958 15052 6010
rect 14756 5956 14812 5958
rect 14836 5956 14892 5958
rect 14916 5956 14972 5958
rect 14996 5956 15052 5958
rect 18206 6554 18262 6556
rect 18286 6554 18342 6556
rect 18366 6554 18422 6556
rect 18446 6554 18502 6556
rect 18206 6502 18232 6554
rect 18232 6502 18262 6554
rect 18286 6502 18296 6554
rect 18296 6502 18342 6554
rect 18366 6502 18412 6554
rect 18412 6502 18422 6554
rect 18446 6502 18476 6554
rect 18476 6502 18502 6554
rect 18206 6500 18262 6502
rect 18286 6500 18342 6502
rect 18366 6500 18422 6502
rect 18446 6500 18502 6502
rect 14756 4922 14812 4924
rect 14836 4922 14892 4924
rect 14916 4922 14972 4924
rect 14996 4922 15052 4924
rect 14756 4870 14782 4922
rect 14782 4870 14812 4922
rect 14836 4870 14846 4922
rect 14846 4870 14892 4922
rect 14916 4870 14962 4922
rect 14962 4870 14972 4922
rect 14996 4870 15026 4922
rect 15026 4870 15052 4922
rect 14756 4868 14812 4870
rect 14836 4868 14892 4870
rect 14916 4868 14972 4870
rect 14996 4868 15052 4870
rect 14756 3834 14812 3836
rect 14836 3834 14892 3836
rect 14916 3834 14972 3836
rect 14996 3834 15052 3836
rect 14756 3782 14782 3834
rect 14782 3782 14812 3834
rect 14836 3782 14846 3834
rect 14846 3782 14892 3834
rect 14916 3782 14962 3834
rect 14962 3782 14972 3834
rect 14996 3782 15026 3834
rect 15026 3782 15052 3834
rect 14756 3780 14812 3782
rect 14836 3780 14892 3782
rect 14916 3780 14972 3782
rect 14996 3780 15052 3782
rect 14756 2746 14812 2748
rect 14836 2746 14892 2748
rect 14916 2746 14972 2748
rect 14996 2746 15052 2748
rect 14756 2694 14782 2746
rect 14782 2694 14812 2746
rect 14836 2694 14846 2746
rect 14846 2694 14892 2746
rect 14916 2694 14962 2746
rect 14962 2694 14972 2746
rect 14996 2694 15026 2746
rect 15026 2694 15052 2746
rect 14756 2692 14812 2694
rect 14836 2692 14892 2694
rect 14916 2692 14972 2694
rect 14996 2692 15052 2694
rect 18206 5466 18262 5468
rect 18286 5466 18342 5468
rect 18366 5466 18422 5468
rect 18446 5466 18502 5468
rect 18206 5414 18232 5466
rect 18232 5414 18262 5466
rect 18286 5414 18296 5466
rect 18296 5414 18342 5466
rect 18366 5414 18412 5466
rect 18412 5414 18422 5466
rect 18446 5414 18476 5466
rect 18476 5414 18502 5466
rect 18206 5412 18262 5414
rect 18286 5412 18342 5414
rect 18366 5412 18422 5414
rect 18446 5412 18502 5414
rect 18206 4378 18262 4380
rect 18286 4378 18342 4380
rect 18366 4378 18422 4380
rect 18446 4378 18502 4380
rect 18206 4326 18232 4378
rect 18232 4326 18262 4378
rect 18286 4326 18296 4378
rect 18296 4326 18342 4378
rect 18366 4326 18412 4378
rect 18412 4326 18422 4378
rect 18446 4326 18476 4378
rect 18476 4326 18502 4378
rect 18206 4324 18262 4326
rect 18286 4324 18342 4326
rect 18366 4324 18422 4326
rect 18446 4324 18502 4326
rect 18206 3290 18262 3292
rect 18286 3290 18342 3292
rect 18366 3290 18422 3292
rect 18446 3290 18502 3292
rect 18206 3238 18232 3290
rect 18232 3238 18262 3290
rect 18286 3238 18296 3290
rect 18296 3238 18342 3290
rect 18366 3238 18412 3290
rect 18412 3238 18422 3290
rect 18446 3238 18476 3290
rect 18476 3238 18502 3290
rect 18206 3236 18262 3238
rect 18286 3236 18342 3238
rect 18366 3236 18422 3238
rect 18446 3236 18502 3238
rect 21086 15680 21142 15736
rect 21086 10240 21142 10296
rect 21086 8200 21142 8256
rect 21086 5480 21142 5536
rect 21086 2760 21142 2816
rect 18206 2202 18262 2204
rect 18286 2202 18342 2204
rect 18366 2202 18422 2204
rect 18446 2202 18502 2204
rect 18206 2150 18232 2202
rect 18232 2150 18262 2202
rect 18286 2150 18296 2202
rect 18296 2150 18342 2202
rect 18366 2150 18412 2202
rect 18412 2150 18422 2202
rect 18446 2150 18476 2202
rect 18476 2150 18502 2202
rect 18206 2148 18262 2150
rect 18286 2148 18342 2150
rect 18366 2148 18422 2150
rect 18446 2148 18502 2150
<< metal3 >>
rect 0 23218 800 23248
rect 1485 23218 1551 23221
rect 0 23216 1551 23218
rect 0 23160 1490 23216
rect 1546 23160 1551 23216
rect 0 23158 1551 23160
rect 0 23128 800 23158
rect 1485 23155 1551 23158
rect 21081 23218 21147 23221
rect 22179 23218 22979 23248
rect 21081 23216 22979 23218
rect 21081 23160 21086 23216
rect 21142 23160 22979 23216
rect 21081 23158 22979 23160
rect 21081 23155 21147 23158
rect 22179 23128 22979 23158
rect 4394 22880 4714 22881
rect 4394 22816 4402 22880
rect 4466 22816 4482 22880
rect 4546 22816 4562 22880
rect 4626 22816 4642 22880
rect 4706 22816 4714 22880
rect 4394 22815 4714 22816
rect 11294 22880 11614 22881
rect 11294 22816 11302 22880
rect 11366 22816 11382 22880
rect 11446 22816 11462 22880
rect 11526 22816 11542 22880
rect 11606 22816 11614 22880
rect 11294 22815 11614 22816
rect 18194 22880 18514 22881
rect 18194 22816 18202 22880
rect 18266 22816 18282 22880
rect 18346 22816 18362 22880
rect 18426 22816 18442 22880
rect 18506 22816 18514 22880
rect 18194 22815 18514 22816
rect 7844 22336 8164 22337
rect 7844 22272 7852 22336
rect 7916 22272 7932 22336
rect 7996 22272 8012 22336
rect 8076 22272 8092 22336
rect 8156 22272 8164 22336
rect 7844 22271 8164 22272
rect 14744 22336 15064 22337
rect 14744 22272 14752 22336
rect 14816 22272 14832 22336
rect 14896 22272 14912 22336
rect 14976 22272 14992 22336
rect 15056 22272 15064 22336
rect 14744 22271 15064 22272
rect 4394 21792 4714 21793
rect 4394 21728 4402 21792
rect 4466 21728 4482 21792
rect 4546 21728 4562 21792
rect 4626 21728 4642 21792
rect 4706 21728 4714 21792
rect 4394 21727 4714 21728
rect 11294 21792 11614 21793
rect 11294 21728 11302 21792
rect 11366 21728 11382 21792
rect 11446 21728 11462 21792
rect 11526 21728 11542 21792
rect 11606 21728 11614 21792
rect 11294 21727 11614 21728
rect 18194 21792 18514 21793
rect 18194 21728 18202 21792
rect 18266 21728 18282 21792
rect 18346 21728 18362 21792
rect 18426 21728 18442 21792
rect 18506 21728 18514 21792
rect 18194 21727 18514 21728
rect 7844 21248 8164 21249
rect 7844 21184 7852 21248
rect 7916 21184 7932 21248
rect 7996 21184 8012 21248
rect 8076 21184 8092 21248
rect 8156 21184 8164 21248
rect 7844 21183 8164 21184
rect 14744 21248 15064 21249
rect 14744 21184 14752 21248
rect 14816 21184 14832 21248
rect 14896 21184 14912 21248
rect 14976 21184 14992 21248
rect 15056 21184 15064 21248
rect 14744 21183 15064 21184
rect 4394 20704 4714 20705
rect 4394 20640 4402 20704
rect 4466 20640 4482 20704
rect 4546 20640 4562 20704
rect 4626 20640 4642 20704
rect 4706 20640 4714 20704
rect 4394 20639 4714 20640
rect 11294 20704 11614 20705
rect 11294 20640 11302 20704
rect 11366 20640 11382 20704
rect 11446 20640 11462 20704
rect 11526 20640 11542 20704
rect 11606 20640 11614 20704
rect 11294 20639 11614 20640
rect 18194 20704 18514 20705
rect 18194 20640 18202 20704
rect 18266 20640 18282 20704
rect 18346 20640 18362 20704
rect 18426 20640 18442 20704
rect 18506 20640 18514 20704
rect 18194 20639 18514 20640
rect 0 20498 800 20528
rect 1393 20498 1459 20501
rect 0 20496 1459 20498
rect 0 20440 1398 20496
rect 1454 20440 1459 20496
rect 0 20438 1459 20440
rect 0 20408 800 20438
rect 1393 20435 1459 20438
rect 20621 20498 20687 20501
rect 22179 20498 22979 20528
rect 20621 20496 22979 20498
rect 20621 20440 20626 20496
rect 20682 20440 22979 20496
rect 20621 20438 22979 20440
rect 20621 20435 20687 20438
rect 22179 20408 22979 20438
rect 7844 20160 8164 20161
rect 7844 20096 7852 20160
rect 7916 20096 7932 20160
rect 7996 20096 8012 20160
rect 8076 20096 8092 20160
rect 8156 20096 8164 20160
rect 7844 20095 8164 20096
rect 14744 20160 15064 20161
rect 14744 20096 14752 20160
rect 14816 20096 14832 20160
rect 14896 20096 14912 20160
rect 14976 20096 14992 20160
rect 15056 20096 15064 20160
rect 14744 20095 15064 20096
rect 4394 19616 4714 19617
rect 4394 19552 4402 19616
rect 4466 19552 4482 19616
rect 4546 19552 4562 19616
rect 4626 19552 4642 19616
rect 4706 19552 4714 19616
rect 4394 19551 4714 19552
rect 11294 19616 11614 19617
rect 11294 19552 11302 19616
rect 11366 19552 11382 19616
rect 11446 19552 11462 19616
rect 11526 19552 11542 19616
rect 11606 19552 11614 19616
rect 11294 19551 11614 19552
rect 18194 19616 18514 19617
rect 18194 19552 18202 19616
rect 18266 19552 18282 19616
rect 18346 19552 18362 19616
rect 18426 19552 18442 19616
rect 18506 19552 18514 19616
rect 18194 19551 18514 19552
rect 7844 19072 8164 19073
rect 7844 19008 7852 19072
rect 7916 19008 7932 19072
rect 7996 19008 8012 19072
rect 8076 19008 8092 19072
rect 8156 19008 8164 19072
rect 7844 19007 8164 19008
rect 14744 19072 15064 19073
rect 14744 19008 14752 19072
rect 14816 19008 14832 19072
rect 14896 19008 14912 19072
rect 14976 19008 14992 19072
rect 15056 19008 15064 19072
rect 14744 19007 15064 19008
rect 4394 18528 4714 18529
rect 4394 18464 4402 18528
rect 4466 18464 4482 18528
rect 4546 18464 4562 18528
rect 4626 18464 4642 18528
rect 4706 18464 4714 18528
rect 4394 18463 4714 18464
rect 11294 18528 11614 18529
rect 11294 18464 11302 18528
rect 11366 18464 11382 18528
rect 11446 18464 11462 18528
rect 11526 18464 11542 18528
rect 11606 18464 11614 18528
rect 11294 18463 11614 18464
rect 18194 18528 18514 18529
rect 18194 18464 18202 18528
rect 18266 18464 18282 18528
rect 18346 18464 18362 18528
rect 18426 18464 18442 18528
rect 18506 18464 18514 18528
rect 18194 18463 18514 18464
rect 7844 17984 8164 17985
rect 7844 17920 7852 17984
rect 7916 17920 7932 17984
rect 7996 17920 8012 17984
rect 8076 17920 8092 17984
rect 8156 17920 8164 17984
rect 7844 17919 8164 17920
rect 14744 17984 15064 17985
rect 14744 17920 14752 17984
rect 14816 17920 14832 17984
rect 14896 17920 14912 17984
rect 14976 17920 14992 17984
rect 15056 17920 15064 17984
rect 14744 17919 15064 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 20621 17778 20687 17781
rect 22179 17778 22979 17808
rect 20621 17776 22979 17778
rect 20621 17720 20626 17776
rect 20682 17720 22979 17776
rect 20621 17718 22979 17720
rect 20621 17715 20687 17718
rect 22179 17688 22979 17718
rect 4394 17440 4714 17441
rect 4394 17376 4402 17440
rect 4466 17376 4482 17440
rect 4546 17376 4562 17440
rect 4626 17376 4642 17440
rect 4706 17376 4714 17440
rect 4394 17375 4714 17376
rect 11294 17440 11614 17441
rect 11294 17376 11302 17440
rect 11366 17376 11382 17440
rect 11446 17376 11462 17440
rect 11526 17376 11542 17440
rect 11606 17376 11614 17440
rect 11294 17375 11614 17376
rect 18194 17440 18514 17441
rect 18194 17376 18202 17440
rect 18266 17376 18282 17440
rect 18346 17376 18362 17440
rect 18426 17376 18442 17440
rect 18506 17376 18514 17440
rect 18194 17375 18514 17376
rect 7844 16896 8164 16897
rect 7844 16832 7852 16896
rect 7916 16832 7932 16896
rect 7996 16832 8012 16896
rect 8076 16832 8092 16896
rect 8156 16832 8164 16896
rect 7844 16831 8164 16832
rect 14744 16896 15064 16897
rect 14744 16832 14752 16896
rect 14816 16832 14832 16896
rect 14896 16832 14912 16896
rect 14976 16832 14992 16896
rect 15056 16832 15064 16896
rect 14744 16831 15064 16832
rect 4394 16352 4714 16353
rect 4394 16288 4402 16352
rect 4466 16288 4482 16352
rect 4546 16288 4562 16352
rect 4626 16288 4642 16352
rect 4706 16288 4714 16352
rect 4394 16287 4714 16288
rect 11294 16352 11614 16353
rect 11294 16288 11302 16352
rect 11366 16288 11382 16352
rect 11446 16288 11462 16352
rect 11526 16288 11542 16352
rect 11606 16288 11614 16352
rect 11294 16287 11614 16288
rect 18194 16352 18514 16353
rect 18194 16288 18202 16352
rect 18266 16288 18282 16352
rect 18346 16288 18362 16352
rect 18426 16288 18442 16352
rect 18506 16288 18514 16352
rect 18194 16287 18514 16288
rect 7844 15808 8164 15809
rect 0 15738 800 15768
rect 7844 15744 7852 15808
rect 7916 15744 7932 15808
rect 7996 15744 8012 15808
rect 8076 15744 8092 15808
rect 8156 15744 8164 15808
rect 7844 15743 8164 15744
rect 14744 15808 15064 15809
rect 14744 15744 14752 15808
rect 14816 15744 14832 15808
rect 14896 15744 14912 15808
rect 14976 15744 14992 15808
rect 15056 15744 15064 15808
rect 14744 15743 15064 15744
rect 1393 15738 1459 15741
rect 0 15736 1459 15738
rect 0 15680 1398 15736
rect 1454 15680 1459 15736
rect 0 15678 1459 15680
rect 0 15648 800 15678
rect 1393 15675 1459 15678
rect 21081 15738 21147 15741
rect 22179 15738 22979 15768
rect 21081 15736 22979 15738
rect 21081 15680 21086 15736
rect 21142 15680 22979 15736
rect 21081 15678 22979 15680
rect 21081 15675 21147 15678
rect 22179 15648 22979 15678
rect 4394 15264 4714 15265
rect 4394 15200 4402 15264
rect 4466 15200 4482 15264
rect 4546 15200 4562 15264
rect 4626 15200 4642 15264
rect 4706 15200 4714 15264
rect 4394 15199 4714 15200
rect 11294 15264 11614 15265
rect 11294 15200 11302 15264
rect 11366 15200 11382 15264
rect 11446 15200 11462 15264
rect 11526 15200 11542 15264
rect 11606 15200 11614 15264
rect 11294 15199 11614 15200
rect 18194 15264 18514 15265
rect 18194 15200 18202 15264
rect 18266 15200 18282 15264
rect 18346 15200 18362 15264
rect 18426 15200 18442 15264
rect 18506 15200 18514 15264
rect 18194 15199 18514 15200
rect 7844 14720 8164 14721
rect 7844 14656 7852 14720
rect 7916 14656 7932 14720
rect 7996 14656 8012 14720
rect 8076 14656 8092 14720
rect 8156 14656 8164 14720
rect 7844 14655 8164 14656
rect 14744 14720 15064 14721
rect 14744 14656 14752 14720
rect 14816 14656 14832 14720
rect 14896 14656 14912 14720
rect 14976 14656 14992 14720
rect 15056 14656 15064 14720
rect 14744 14655 15064 14656
rect 4394 14176 4714 14177
rect 4394 14112 4402 14176
rect 4466 14112 4482 14176
rect 4546 14112 4562 14176
rect 4626 14112 4642 14176
rect 4706 14112 4714 14176
rect 4394 14111 4714 14112
rect 11294 14176 11614 14177
rect 11294 14112 11302 14176
rect 11366 14112 11382 14176
rect 11446 14112 11462 14176
rect 11526 14112 11542 14176
rect 11606 14112 11614 14176
rect 11294 14111 11614 14112
rect 18194 14176 18514 14177
rect 18194 14112 18202 14176
rect 18266 14112 18282 14176
rect 18346 14112 18362 14176
rect 18426 14112 18442 14176
rect 18506 14112 18514 14176
rect 18194 14111 18514 14112
rect 7844 13632 8164 13633
rect 7844 13568 7852 13632
rect 7916 13568 7932 13632
rect 7996 13568 8012 13632
rect 8076 13568 8092 13632
rect 8156 13568 8164 13632
rect 7844 13567 8164 13568
rect 14744 13632 15064 13633
rect 14744 13568 14752 13632
rect 14816 13568 14832 13632
rect 14896 13568 14912 13632
rect 14976 13568 14992 13632
rect 15056 13568 15064 13632
rect 14744 13567 15064 13568
rect 4394 13088 4714 13089
rect 0 13018 800 13048
rect 4394 13024 4402 13088
rect 4466 13024 4482 13088
rect 4546 13024 4562 13088
rect 4626 13024 4642 13088
rect 4706 13024 4714 13088
rect 4394 13023 4714 13024
rect 11294 13088 11614 13089
rect 11294 13024 11302 13088
rect 11366 13024 11382 13088
rect 11446 13024 11462 13088
rect 11526 13024 11542 13088
rect 11606 13024 11614 13088
rect 11294 13023 11614 13024
rect 18194 13088 18514 13089
rect 18194 13024 18202 13088
rect 18266 13024 18282 13088
rect 18346 13024 18362 13088
rect 18426 13024 18442 13088
rect 18506 13024 18514 13088
rect 18194 13023 18514 13024
rect 1485 13018 1551 13021
rect 0 13016 1551 13018
rect 0 12960 1490 13016
rect 1546 12960 1551 13016
rect 0 12958 1551 12960
rect 0 12928 800 12958
rect 1485 12955 1551 12958
rect 20621 13018 20687 13021
rect 22179 13018 22979 13048
rect 20621 13016 22979 13018
rect 20621 12960 20626 13016
rect 20682 12960 22979 13016
rect 20621 12958 22979 12960
rect 20621 12955 20687 12958
rect 22179 12928 22979 12958
rect 7189 12610 7255 12613
rect 7557 12610 7623 12613
rect 7189 12608 7623 12610
rect 7189 12552 7194 12608
rect 7250 12552 7562 12608
rect 7618 12552 7623 12608
rect 7189 12550 7623 12552
rect 7189 12547 7255 12550
rect 7557 12547 7623 12550
rect 7844 12544 8164 12545
rect 7844 12480 7852 12544
rect 7916 12480 7932 12544
rect 7996 12480 8012 12544
rect 8076 12480 8092 12544
rect 8156 12480 8164 12544
rect 7844 12479 8164 12480
rect 14744 12544 15064 12545
rect 14744 12480 14752 12544
rect 14816 12480 14832 12544
rect 14896 12480 14912 12544
rect 14976 12480 14992 12544
rect 15056 12480 15064 12544
rect 14744 12479 15064 12480
rect 4394 12000 4714 12001
rect 4394 11936 4402 12000
rect 4466 11936 4482 12000
rect 4546 11936 4562 12000
rect 4626 11936 4642 12000
rect 4706 11936 4714 12000
rect 4394 11935 4714 11936
rect 11294 12000 11614 12001
rect 11294 11936 11302 12000
rect 11366 11936 11382 12000
rect 11446 11936 11462 12000
rect 11526 11936 11542 12000
rect 11606 11936 11614 12000
rect 11294 11935 11614 11936
rect 18194 12000 18514 12001
rect 18194 11936 18202 12000
rect 18266 11936 18282 12000
rect 18346 11936 18362 12000
rect 18426 11936 18442 12000
rect 18506 11936 18514 12000
rect 18194 11935 18514 11936
rect 7844 11456 8164 11457
rect 7844 11392 7852 11456
rect 7916 11392 7932 11456
rect 7996 11392 8012 11456
rect 8076 11392 8092 11456
rect 8156 11392 8164 11456
rect 7844 11391 8164 11392
rect 14744 11456 15064 11457
rect 14744 11392 14752 11456
rect 14816 11392 14832 11456
rect 14896 11392 14912 11456
rect 14976 11392 14992 11456
rect 15056 11392 15064 11456
rect 14744 11391 15064 11392
rect 4394 10912 4714 10913
rect 4394 10848 4402 10912
rect 4466 10848 4482 10912
rect 4546 10848 4562 10912
rect 4626 10848 4642 10912
rect 4706 10848 4714 10912
rect 4394 10847 4714 10848
rect 11294 10912 11614 10913
rect 11294 10848 11302 10912
rect 11366 10848 11382 10912
rect 11446 10848 11462 10912
rect 11526 10848 11542 10912
rect 11606 10848 11614 10912
rect 11294 10847 11614 10848
rect 18194 10912 18514 10913
rect 18194 10848 18202 10912
rect 18266 10848 18282 10912
rect 18346 10848 18362 10912
rect 18426 10848 18442 10912
rect 18506 10848 18514 10912
rect 18194 10847 18514 10848
rect 7844 10368 8164 10369
rect 0 10298 800 10328
rect 7844 10304 7852 10368
rect 7916 10304 7932 10368
rect 7996 10304 8012 10368
rect 8076 10304 8092 10368
rect 8156 10304 8164 10368
rect 7844 10303 8164 10304
rect 14744 10368 15064 10369
rect 14744 10304 14752 10368
rect 14816 10304 14832 10368
rect 14896 10304 14912 10368
rect 14976 10304 14992 10368
rect 15056 10304 15064 10368
rect 14744 10303 15064 10304
rect 1485 10298 1551 10301
rect 0 10296 1551 10298
rect 0 10240 1490 10296
rect 1546 10240 1551 10296
rect 0 10238 1551 10240
rect 0 10208 800 10238
rect 1485 10235 1551 10238
rect 21081 10298 21147 10301
rect 22179 10298 22979 10328
rect 21081 10296 22979 10298
rect 21081 10240 21086 10296
rect 21142 10240 22979 10296
rect 21081 10238 22979 10240
rect 21081 10235 21147 10238
rect 22179 10208 22979 10238
rect 4394 9824 4714 9825
rect 4394 9760 4402 9824
rect 4466 9760 4482 9824
rect 4546 9760 4562 9824
rect 4626 9760 4642 9824
rect 4706 9760 4714 9824
rect 4394 9759 4714 9760
rect 11294 9824 11614 9825
rect 11294 9760 11302 9824
rect 11366 9760 11382 9824
rect 11446 9760 11462 9824
rect 11526 9760 11542 9824
rect 11606 9760 11614 9824
rect 11294 9759 11614 9760
rect 18194 9824 18514 9825
rect 18194 9760 18202 9824
rect 18266 9760 18282 9824
rect 18346 9760 18362 9824
rect 18426 9760 18442 9824
rect 18506 9760 18514 9824
rect 18194 9759 18514 9760
rect 7844 9280 8164 9281
rect 7844 9216 7852 9280
rect 7916 9216 7932 9280
rect 7996 9216 8012 9280
rect 8076 9216 8092 9280
rect 8156 9216 8164 9280
rect 7844 9215 8164 9216
rect 14744 9280 15064 9281
rect 14744 9216 14752 9280
rect 14816 9216 14832 9280
rect 14896 9216 14912 9280
rect 14976 9216 14992 9280
rect 15056 9216 15064 9280
rect 14744 9215 15064 9216
rect 4394 8736 4714 8737
rect 4394 8672 4402 8736
rect 4466 8672 4482 8736
rect 4546 8672 4562 8736
rect 4626 8672 4642 8736
rect 4706 8672 4714 8736
rect 4394 8671 4714 8672
rect 11294 8736 11614 8737
rect 11294 8672 11302 8736
rect 11366 8672 11382 8736
rect 11446 8672 11462 8736
rect 11526 8672 11542 8736
rect 11606 8672 11614 8736
rect 11294 8671 11614 8672
rect 18194 8736 18514 8737
rect 18194 8672 18202 8736
rect 18266 8672 18282 8736
rect 18346 8672 18362 8736
rect 18426 8672 18442 8736
rect 18506 8672 18514 8736
rect 18194 8671 18514 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 21081 8258 21147 8261
rect 22179 8258 22979 8288
rect 21081 8256 22979 8258
rect 21081 8200 21086 8256
rect 21142 8200 22979 8256
rect 21081 8198 22979 8200
rect 21081 8195 21147 8198
rect 7844 8192 8164 8193
rect 7844 8128 7852 8192
rect 7916 8128 7932 8192
rect 7996 8128 8012 8192
rect 8076 8128 8092 8192
rect 8156 8128 8164 8192
rect 7844 8127 8164 8128
rect 14744 8192 15064 8193
rect 14744 8128 14752 8192
rect 14816 8128 14832 8192
rect 14896 8128 14912 8192
rect 14976 8128 14992 8192
rect 15056 8128 15064 8192
rect 22179 8168 22979 8198
rect 14744 8127 15064 8128
rect 4394 7648 4714 7649
rect 4394 7584 4402 7648
rect 4466 7584 4482 7648
rect 4546 7584 4562 7648
rect 4626 7584 4642 7648
rect 4706 7584 4714 7648
rect 4394 7583 4714 7584
rect 11294 7648 11614 7649
rect 11294 7584 11302 7648
rect 11366 7584 11382 7648
rect 11446 7584 11462 7648
rect 11526 7584 11542 7648
rect 11606 7584 11614 7648
rect 11294 7583 11614 7584
rect 18194 7648 18514 7649
rect 18194 7584 18202 7648
rect 18266 7584 18282 7648
rect 18346 7584 18362 7648
rect 18426 7584 18442 7648
rect 18506 7584 18514 7648
rect 18194 7583 18514 7584
rect 7844 7104 8164 7105
rect 7844 7040 7852 7104
rect 7916 7040 7932 7104
rect 7996 7040 8012 7104
rect 8076 7040 8092 7104
rect 8156 7040 8164 7104
rect 7844 7039 8164 7040
rect 14744 7104 15064 7105
rect 14744 7040 14752 7104
rect 14816 7040 14832 7104
rect 14896 7040 14912 7104
rect 14976 7040 14992 7104
rect 15056 7040 15064 7104
rect 14744 7039 15064 7040
rect 4394 6560 4714 6561
rect 4394 6496 4402 6560
rect 4466 6496 4482 6560
rect 4546 6496 4562 6560
rect 4626 6496 4642 6560
rect 4706 6496 4714 6560
rect 4394 6495 4714 6496
rect 11294 6560 11614 6561
rect 11294 6496 11302 6560
rect 11366 6496 11382 6560
rect 11446 6496 11462 6560
rect 11526 6496 11542 6560
rect 11606 6496 11614 6560
rect 11294 6495 11614 6496
rect 18194 6560 18514 6561
rect 18194 6496 18202 6560
rect 18266 6496 18282 6560
rect 18346 6496 18362 6560
rect 18426 6496 18442 6560
rect 18506 6496 18514 6560
rect 18194 6495 18514 6496
rect 7844 6016 8164 6017
rect 7844 5952 7852 6016
rect 7916 5952 7932 6016
rect 7996 5952 8012 6016
rect 8076 5952 8092 6016
rect 8156 5952 8164 6016
rect 7844 5951 8164 5952
rect 14744 6016 15064 6017
rect 14744 5952 14752 6016
rect 14816 5952 14832 6016
rect 14896 5952 14912 6016
rect 14976 5952 14992 6016
rect 15056 5952 15064 6016
rect 14744 5951 15064 5952
rect 0 5538 800 5568
rect 1485 5538 1551 5541
rect 0 5536 1551 5538
rect 0 5480 1490 5536
rect 1546 5480 1551 5536
rect 0 5478 1551 5480
rect 0 5448 800 5478
rect 1485 5475 1551 5478
rect 21081 5538 21147 5541
rect 22179 5538 22979 5568
rect 21081 5536 22979 5538
rect 21081 5480 21086 5536
rect 21142 5480 22979 5536
rect 21081 5478 22979 5480
rect 21081 5475 21147 5478
rect 4394 5472 4714 5473
rect 4394 5408 4402 5472
rect 4466 5408 4482 5472
rect 4546 5408 4562 5472
rect 4626 5408 4642 5472
rect 4706 5408 4714 5472
rect 4394 5407 4714 5408
rect 11294 5472 11614 5473
rect 11294 5408 11302 5472
rect 11366 5408 11382 5472
rect 11446 5408 11462 5472
rect 11526 5408 11542 5472
rect 11606 5408 11614 5472
rect 11294 5407 11614 5408
rect 18194 5472 18514 5473
rect 18194 5408 18202 5472
rect 18266 5408 18282 5472
rect 18346 5408 18362 5472
rect 18426 5408 18442 5472
rect 18506 5408 18514 5472
rect 22179 5448 22979 5478
rect 18194 5407 18514 5408
rect 7844 4928 8164 4929
rect 7844 4864 7852 4928
rect 7916 4864 7932 4928
rect 7996 4864 8012 4928
rect 8076 4864 8092 4928
rect 8156 4864 8164 4928
rect 7844 4863 8164 4864
rect 14744 4928 15064 4929
rect 14744 4864 14752 4928
rect 14816 4864 14832 4928
rect 14896 4864 14912 4928
rect 14976 4864 14992 4928
rect 15056 4864 15064 4928
rect 14744 4863 15064 4864
rect 4394 4384 4714 4385
rect 4394 4320 4402 4384
rect 4466 4320 4482 4384
rect 4546 4320 4562 4384
rect 4626 4320 4642 4384
rect 4706 4320 4714 4384
rect 4394 4319 4714 4320
rect 11294 4384 11614 4385
rect 11294 4320 11302 4384
rect 11366 4320 11382 4384
rect 11446 4320 11462 4384
rect 11526 4320 11542 4384
rect 11606 4320 11614 4384
rect 11294 4319 11614 4320
rect 18194 4384 18514 4385
rect 18194 4320 18202 4384
rect 18266 4320 18282 4384
rect 18346 4320 18362 4384
rect 18426 4320 18442 4384
rect 18506 4320 18514 4384
rect 18194 4319 18514 4320
rect 7844 3840 8164 3841
rect 7844 3776 7852 3840
rect 7916 3776 7932 3840
rect 7996 3776 8012 3840
rect 8076 3776 8092 3840
rect 8156 3776 8164 3840
rect 7844 3775 8164 3776
rect 14744 3840 15064 3841
rect 14744 3776 14752 3840
rect 14816 3776 14832 3840
rect 14896 3776 14912 3840
rect 14976 3776 14992 3840
rect 15056 3776 15064 3840
rect 14744 3775 15064 3776
rect 4394 3296 4714 3297
rect 4394 3232 4402 3296
rect 4466 3232 4482 3296
rect 4546 3232 4562 3296
rect 4626 3232 4642 3296
rect 4706 3232 4714 3296
rect 4394 3231 4714 3232
rect 11294 3296 11614 3297
rect 11294 3232 11302 3296
rect 11366 3232 11382 3296
rect 11446 3232 11462 3296
rect 11526 3232 11542 3296
rect 11606 3232 11614 3296
rect 11294 3231 11614 3232
rect 18194 3296 18514 3297
rect 18194 3232 18202 3296
rect 18266 3232 18282 3296
rect 18346 3232 18362 3296
rect 18426 3232 18442 3296
rect 18506 3232 18514 3296
rect 18194 3231 18514 3232
rect 0 2818 800 2848
rect 1393 2818 1459 2821
rect 0 2816 1459 2818
rect 0 2760 1398 2816
rect 1454 2760 1459 2816
rect 0 2758 1459 2760
rect 0 2728 800 2758
rect 1393 2755 1459 2758
rect 21081 2818 21147 2821
rect 22179 2818 22979 2848
rect 21081 2816 22979 2818
rect 21081 2760 21086 2816
rect 21142 2760 22979 2816
rect 21081 2758 22979 2760
rect 21081 2755 21147 2758
rect 7844 2752 8164 2753
rect 7844 2688 7852 2752
rect 7916 2688 7932 2752
rect 7996 2688 8012 2752
rect 8076 2688 8092 2752
rect 8156 2688 8164 2752
rect 7844 2687 8164 2688
rect 14744 2752 15064 2753
rect 14744 2688 14752 2752
rect 14816 2688 14832 2752
rect 14896 2688 14912 2752
rect 14976 2688 14992 2752
rect 15056 2688 15064 2752
rect 22179 2728 22979 2758
rect 14744 2687 15064 2688
rect 4394 2208 4714 2209
rect 4394 2144 4402 2208
rect 4466 2144 4482 2208
rect 4546 2144 4562 2208
rect 4626 2144 4642 2208
rect 4706 2144 4714 2208
rect 4394 2143 4714 2144
rect 11294 2208 11614 2209
rect 11294 2144 11302 2208
rect 11366 2144 11382 2208
rect 11446 2144 11462 2208
rect 11526 2144 11542 2208
rect 11606 2144 11614 2208
rect 11294 2143 11614 2144
rect 18194 2208 18514 2209
rect 18194 2144 18202 2208
rect 18266 2144 18282 2208
rect 18346 2144 18362 2208
rect 18426 2144 18442 2208
rect 18506 2144 18514 2208
rect 18194 2143 18514 2144
<< via3 >>
rect 4402 22876 4466 22880
rect 4402 22820 4406 22876
rect 4406 22820 4462 22876
rect 4462 22820 4466 22876
rect 4402 22816 4466 22820
rect 4482 22876 4546 22880
rect 4482 22820 4486 22876
rect 4486 22820 4542 22876
rect 4542 22820 4546 22876
rect 4482 22816 4546 22820
rect 4562 22876 4626 22880
rect 4562 22820 4566 22876
rect 4566 22820 4622 22876
rect 4622 22820 4626 22876
rect 4562 22816 4626 22820
rect 4642 22876 4706 22880
rect 4642 22820 4646 22876
rect 4646 22820 4702 22876
rect 4702 22820 4706 22876
rect 4642 22816 4706 22820
rect 11302 22876 11366 22880
rect 11302 22820 11306 22876
rect 11306 22820 11362 22876
rect 11362 22820 11366 22876
rect 11302 22816 11366 22820
rect 11382 22876 11446 22880
rect 11382 22820 11386 22876
rect 11386 22820 11442 22876
rect 11442 22820 11446 22876
rect 11382 22816 11446 22820
rect 11462 22876 11526 22880
rect 11462 22820 11466 22876
rect 11466 22820 11522 22876
rect 11522 22820 11526 22876
rect 11462 22816 11526 22820
rect 11542 22876 11606 22880
rect 11542 22820 11546 22876
rect 11546 22820 11602 22876
rect 11602 22820 11606 22876
rect 11542 22816 11606 22820
rect 18202 22876 18266 22880
rect 18202 22820 18206 22876
rect 18206 22820 18262 22876
rect 18262 22820 18266 22876
rect 18202 22816 18266 22820
rect 18282 22876 18346 22880
rect 18282 22820 18286 22876
rect 18286 22820 18342 22876
rect 18342 22820 18346 22876
rect 18282 22816 18346 22820
rect 18362 22876 18426 22880
rect 18362 22820 18366 22876
rect 18366 22820 18422 22876
rect 18422 22820 18426 22876
rect 18362 22816 18426 22820
rect 18442 22876 18506 22880
rect 18442 22820 18446 22876
rect 18446 22820 18502 22876
rect 18502 22820 18506 22876
rect 18442 22816 18506 22820
rect 7852 22332 7916 22336
rect 7852 22276 7856 22332
rect 7856 22276 7912 22332
rect 7912 22276 7916 22332
rect 7852 22272 7916 22276
rect 7932 22332 7996 22336
rect 7932 22276 7936 22332
rect 7936 22276 7992 22332
rect 7992 22276 7996 22332
rect 7932 22272 7996 22276
rect 8012 22332 8076 22336
rect 8012 22276 8016 22332
rect 8016 22276 8072 22332
rect 8072 22276 8076 22332
rect 8012 22272 8076 22276
rect 8092 22332 8156 22336
rect 8092 22276 8096 22332
rect 8096 22276 8152 22332
rect 8152 22276 8156 22332
rect 8092 22272 8156 22276
rect 14752 22332 14816 22336
rect 14752 22276 14756 22332
rect 14756 22276 14812 22332
rect 14812 22276 14816 22332
rect 14752 22272 14816 22276
rect 14832 22332 14896 22336
rect 14832 22276 14836 22332
rect 14836 22276 14892 22332
rect 14892 22276 14896 22332
rect 14832 22272 14896 22276
rect 14912 22332 14976 22336
rect 14912 22276 14916 22332
rect 14916 22276 14972 22332
rect 14972 22276 14976 22332
rect 14912 22272 14976 22276
rect 14992 22332 15056 22336
rect 14992 22276 14996 22332
rect 14996 22276 15052 22332
rect 15052 22276 15056 22332
rect 14992 22272 15056 22276
rect 4402 21788 4466 21792
rect 4402 21732 4406 21788
rect 4406 21732 4462 21788
rect 4462 21732 4466 21788
rect 4402 21728 4466 21732
rect 4482 21788 4546 21792
rect 4482 21732 4486 21788
rect 4486 21732 4542 21788
rect 4542 21732 4546 21788
rect 4482 21728 4546 21732
rect 4562 21788 4626 21792
rect 4562 21732 4566 21788
rect 4566 21732 4622 21788
rect 4622 21732 4626 21788
rect 4562 21728 4626 21732
rect 4642 21788 4706 21792
rect 4642 21732 4646 21788
rect 4646 21732 4702 21788
rect 4702 21732 4706 21788
rect 4642 21728 4706 21732
rect 11302 21788 11366 21792
rect 11302 21732 11306 21788
rect 11306 21732 11362 21788
rect 11362 21732 11366 21788
rect 11302 21728 11366 21732
rect 11382 21788 11446 21792
rect 11382 21732 11386 21788
rect 11386 21732 11442 21788
rect 11442 21732 11446 21788
rect 11382 21728 11446 21732
rect 11462 21788 11526 21792
rect 11462 21732 11466 21788
rect 11466 21732 11522 21788
rect 11522 21732 11526 21788
rect 11462 21728 11526 21732
rect 11542 21788 11606 21792
rect 11542 21732 11546 21788
rect 11546 21732 11602 21788
rect 11602 21732 11606 21788
rect 11542 21728 11606 21732
rect 18202 21788 18266 21792
rect 18202 21732 18206 21788
rect 18206 21732 18262 21788
rect 18262 21732 18266 21788
rect 18202 21728 18266 21732
rect 18282 21788 18346 21792
rect 18282 21732 18286 21788
rect 18286 21732 18342 21788
rect 18342 21732 18346 21788
rect 18282 21728 18346 21732
rect 18362 21788 18426 21792
rect 18362 21732 18366 21788
rect 18366 21732 18422 21788
rect 18422 21732 18426 21788
rect 18362 21728 18426 21732
rect 18442 21788 18506 21792
rect 18442 21732 18446 21788
rect 18446 21732 18502 21788
rect 18502 21732 18506 21788
rect 18442 21728 18506 21732
rect 7852 21244 7916 21248
rect 7852 21188 7856 21244
rect 7856 21188 7912 21244
rect 7912 21188 7916 21244
rect 7852 21184 7916 21188
rect 7932 21244 7996 21248
rect 7932 21188 7936 21244
rect 7936 21188 7992 21244
rect 7992 21188 7996 21244
rect 7932 21184 7996 21188
rect 8012 21244 8076 21248
rect 8012 21188 8016 21244
rect 8016 21188 8072 21244
rect 8072 21188 8076 21244
rect 8012 21184 8076 21188
rect 8092 21244 8156 21248
rect 8092 21188 8096 21244
rect 8096 21188 8152 21244
rect 8152 21188 8156 21244
rect 8092 21184 8156 21188
rect 14752 21244 14816 21248
rect 14752 21188 14756 21244
rect 14756 21188 14812 21244
rect 14812 21188 14816 21244
rect 14752 21184 14816 21188
rect 14832 21244 14896 21248
rect 14832 21188 14836 21244
rect 14836 21188 14892 21244
rect 14892 21188 14896 21244
rect 14832 21184 14896 21188
rect 14912 21244 14976 21248
rect 14912 21188 14916 21244
rect 14916 21188 14972 21244
rect 14972 21188 14976 21244
rect 14912 21184 14976 21188
rect 14992 21244 15056 21248
rect 14992 21188 14996 21244
rect 14996 21188 15052 21244
rect 15052 21188 15056 21244
rect 14992 21184 15056 21188
rect 4402 20700 4466 20704
rect 4402 20644 4406 20700
rect 4406 20644 4462 20700
rect 4462 20644 4466 20700
rect 4402 20640 4466 20644
rect 4482 20700 4546 20704
rect 4482 20644 4486 20700
rect 4486 20644 4542 20700
rect 4542 20644 4546 20700
rect 4482 20640 4546 20644
rect 4562 20700 4626 20704
rect 4562 20644 4566 20700
rect 4566 20644 4622 20700
rect 4622 20644 4626 20700
rect 4562 20640 4626 20644
rect 4642 20700 4706 20704
rect 4642 20644 4646 20700
rect 4646 20644 4702 20700
rect 4702 20644 4706 20700
rect 4642 20640 4706 20644
rect 11302 20700 11366 20704
rect 11302 20644 11306 20700
rect 11306 20644 11362 20700
rect 11362 20644 11366 20700
rect 11302 20640 11366 20644
rect 11382 20700 11446 20704
rect 11382 20644 11386 20700
rect 11386 20644 11442 20700
rect 11442 20644 11446 20700
rect 11382 20640 11446 20644
rect 11462 20700 11526 20704
rect 11462 20644 11466 20700
rect 11466 20644 11522 20700
rect 11522 20644 11526 20700
rect 11462 20640 11526 20644
rect 11542 20700 11606 20704
rect 11542 20644 11546 20700
rect 11546 20644 11602 20700
rect 11602 20644 11606 20700
rect 11542 20640 11606 20644
rect 18202 20700 18266 20704
rect 18202 20644 18206 20700
rect 18206 20644 18262 20700
rect 18262 20644 18266 20700
rect 18202 20640 18266 20644
rect 18282 20700 18346 20704
rect 18282 20644 18286 20700
rect 18286 20644 18342 20700
rect 18342 20644 18346 20700
rect 18282 20640 18346 20644
rect 18362 20700 18426 20704
rect 18362 20644 18366 20700
rect 18366 20644 18422 20700
rect 18422 20644 18426 20700
rect 18362 20640 18426 20644
rect 18442 20700 18506 20704
rect 18442 20644 18446 20700
rect 18446 20644 18502 20700
rect 18502 20644 18506 20700
rect 18442 20640 18506 20644
rect 7852 20156 7916 20160
rect 7852 20100 7856 20156
rect 7856 20100 7912 20156
rect 7912 20100 7916 20156
rect 7852 20096 7916 20100
rect 7932 20156 7996 20160
rect 7932 20100 7936 20156
rect 7936 20100 7992 20156
rect 7992 20100 7996 20156
rect 7932 20096 7996 20100
rect 8012 20156 8076 20160
rect 8012 20100 8016 20156
rect 8016 20100 8072 20156
rect 8072 20100 8076 20156
rect 8012 20096 8076 20100
rect 8092 20156 8156 20160
rect 8092 20100 8096 20156
rect 8096 20100 8152 20156
rect 8152 20100 8156 20156
rect 8092 20096 8156 20100
rect 14752 20156 14816 20160
rect 14752 20100 14756 20156
rect 14756 20100 14812 20156
rect 14812 20100 14816 20156
rect 14752 20096 14816 20100
rect 14832 20156 14896 20160
rect 14832 20100 14836 20156
rect 14836 20100 14892 20156
rect 14892 20100 14896 20156
rect 14832 20096 14896 20100
rect 14912 20156 14976 20160
rect 14912 20100 14916 20156
rect 14916 20100 14972 20156
rect 14972 20100 14976 20156
rect 14912 20096 14976 20100
rect 14992 20156 15056 20160
rect 14992 20100 14996 20156
rect 14996 20100 15052 20156
rect 15052 20100 15056 20156
rect 14992 20096 15056 20100
rect 4402 19612 4466 19616
rect 4402 19556 4406 19612
rect 4406 19556 4462 19612
rect 4462 19556 4466 19612
rect 4402 19552 4466 19556
rect 4482 19612 4546 19616
rect 4482 19556 4486 19612
rect 4486 19556 4542 19612
rect 4542 19556 4546 19612
rect 4482 19552 4546 19556
rect 4562 19612 4626 19616
rect 4562 19556 4566 19612
rect 4566 19556 4622 19612
rect 4622 19556 4626 19612
rect 4562 19552 4626 19556
rect 4642 19612 4706 19616
rect 4642 19556 4646 19612
rect 4646 19556 4702 19612
rect 4702 19556 4706 19612
rect 4642 19552 4706 19556
rect 11302 19612 11366 19616
rect 11302 19556 11306 19612
rect 11306 19556 11362 19612
rect 11362 19556 11366 19612
rect 11302 19552 11366 19556
rect 11382 19612 11446 19616
rect 11382 19556 11386 19612
rect 11386 19556 11442 19612
rect 11442 19556 11446 19612
rect 11382 19552 11446 19556
rect 11462 19612 11526 19616
rect 11462 19556 11466 19612
rect 11466 19556 11522 19612
rect 11522 19556 11526 19612
rect 11462 19552 11526 19556
rect 11542 19612 11606 19616
rect 11542 19556 11546 19612
rect 11546 19556 11602 19612
rect 11602 19556 11606 19612
rect 11542 19552 11606 19556
rect 18202 19612 18266 19616
rect 18202 19556 18206 19612
rect 18206 19556 18262 19612
rect 18262 19556 18266 19612
rect 18202 19552 18266 19556
rect 18282 19612 18346 19616
rect 18282 19556 18286 19612
rect 18286 19556 18342 19612
rect 18342 19556 18346 19612
rect 18282 19552 18346 19556
rect 18362 19612 18426 19616
rect 18362 19556 18366 19612
rect 18366 19556 18422 19612
rect 18422 19556 18426 19612
rect 18362 19552 18426 19556
rect 18442 19612 18506 19616
rect 18442 19556 18446 19612
rect 18446 19556 18502 19612
rect 18502 19556 18506 19612
rect 18442 19552 18506 19556
rect 7852 19068 7916 19072
rect 7852 19012 7856 19068
rect 7856 19012 7912 19068
rect 7912 19012 7916 19068
rect 7852 19008 7916 19012
rect 7932 19068 7996 19072
rect 7932 19012 7936 19068
rect 7936 19012 7992 19068
rect 7992 19012 7996 19068
rect 7932 19008 7996 19012
rect 8012 19068 8076 19072
rect 8012 19012 8016 19068
rect 8016 19012 8072 19068
rect 8072 19012 8076 19068
rect 8012 19008 8076 19012
rect 8092 19068 8156 19072
rect 8092 19012 8096 19068
rect 8096 19012 8152 19068
rect 8152 19012 8156 19068
rect 8092 19008 8156 19012
rect 14752 19068 14816 19072
rect 14752 19012 14756 19068
rect 14756 19012 14812 19068
rect 14812 19012 14816 19068
rect 14752 19008 14816 19012
rect 14832 19068 14896 19072
rect 14832 19012 14836 19068
rect 14836 19012 14892 19068
rect 14892 19012 14896 19068
rect 14832 19008 14896 19012
rect 14912 19068 14976 19072
rect 14912 19012 14916 19068
rect 14916 19012 14972 19068
rect 14972 19012 14976 19068
rect 14912 19008 14976 19012
rect 14992 19068 15056 19072
rect 14992 19012 14996 19068
rect 14996 19012 15052 19068
rect 15052 19012 15056 19068
rect 14992 19008 15056 19012
rect 4402 18524 4466 18528
rect 4402 18468 4406 18524
rect 4406 18468 4462 18524
rect 4462 18468 4466 18524
rect 4402 18464 4466 18468
rect 4482 18524 4546 18528
rect 4482 18468 4486 18524
rect 4486 18468 4542 18524
rect 4542 18468 4546 18524
rect 4482 18464 4546 18468
rect 4562 18524 4626 18528
rect 4562 18468 4566 18524
rect 4566 18468 4622 18524
rect 4622 18468 4626 18524
rect 4562 18464 4626 18468
rect 4642 18524 4706 18528
rect 4642 18468 4646 18524
rect 4646 18468 4702 18524
rect 4702 18468 4706 18524
rect 4642 18464 4706 18468
rect 11302 18524 11366 18528
rect 11302 18468 11306 18524
rect 11306 18468 11362 18524
rect 11362 18468 11366 18524
rect 11302 18464 11366 18468
rect 11382 18524 11446 18528
rect 11382 18468 11386 18524
rect 11386 18468 11442 18524
rect 11442 18468 11446 18524
rect 11382 18464 11446 18468
rect 11462 18524 11526 18528
rect 11462 18468 11466 18524
rect 11466 18468 11522 18524
rect 11522 18468 11526 18524
rect 11462 18464 11526 18468
rect 11542 18524 11606 18528
rect 11542 18468 11546 18524
rect 11546 18468 11602 18524
rect 11602 18468 11606 18524
rect 11542 18464 11606 18468
rect 18202 18524 18266 18528
rect 18202 18468 18206 18524
rect 18206 18468 18262 18524
rect 18262 18468 18266 18524
rect 18202 18464 18266 18468
rect 18282 18524 18346 18528
rect 18282 18468 18286 18524
rect 18286 18468 18342 18524
rect 18342 18468 18346 18524
rect 18282 18464 18346 18468
rect 18362 18524 18426 18528
rect 18362 18468 18366 18524
rect 18366 18468 18422 18524
rect 18422 18468 18426 18524
rect 18362 18464 18426 18468
rect 18442 18524 18506 18528
rect 18442 18468 18446 18524
rect 18446 18468 18502 18524
rect 18502 18468 18506 18524
rect 18442 18464 18506 18468
rect 7852 17980 7916 17984
rect 7852 17924 7856 17980
rect 7856 17924 7912 17980
rect 7912 17924 7916 17980
rect 7852 17920 7916 17924
rect 7932 17980 7996 17984
rect 7932 17924 7936 17980
rect 7936 17924 7992 17980
rect 7992 17924 7996 17980
rect 7932 17920 7996 17924
rect 8012 17980 8076 17984
rect 8012 17924 8016 17980
rect 8016 17924 8072 17980
rect 8072 17924 8076 17980
rect 8012 17920 8076 17924
rect 8092 17980 8156 17984
rect 8092 17924 8096 17980
rect 8096 17924 8152 17980
rect 8152 17924 8156 17980
rect 8092 17920 8156 17924
rect 14752 17980 14816 17984
rect 14752 17924 14756 17980
rect 14756 17924 14812 17980
rect 14812 17924 14816 17980
rect 14752 17920 14816 17924
rect 14832 17980 14896 17984
rect 14832 17924 14836 17980
rect 14836 17924 14892 17980
rect 14892 17924 14896 17980
rect 14832 17920 14896 17924
rect 14912 17980 14976 17984
rect 14912 17924 14916 17980
rect 14916 17924 14972 17980
rect 14972 17924 14976 17980
rect 14912 17920 14976 17924
rect 14992 17980 15056 17984
rect 14992 17924 14996 17980
rect 14996 17924 15052 17980
rect 15052 17924 15056 17980
rect 14992 17920 15056 17924
rect 4402 17436 4466 17440
rect 4402 17380 4406 17436
rect 4406 17380 4462 17436
rect 4462 17380 4466 17436
rect 4402 17376 4466 17380
rect 4482 17436 4546 17440
rect 4482 17380 4486 17436
rect 4486 17380 4542 17436
rect 4542 17380 4546 17436
rect 4482 17376 4546 17380
rect 4562 17436 4626 17440
rect 4562 17380 4566 17436
rect 4566 17380 4622 17436
rect 4622 17380 4626 17436
rect 4562 17376 4626 17380
rect 4642 17436 4706 17440
rect 4642 17380 4646 17436
rect 4646 17380 4702 17436
rect 4702 17380 4706 17436
rect 4642 17376 4706 17380
rect 11302 17436 11366 17440
rect 11302 17380 11306 17436
rect 11306 17380 11362 17436
rect 11362 17380 11366 17436
rect 11302 17376 11366 17380
rect 11382 17436 11446 17440
rect 11382 17380 11386 17436
rect 11386 17380 11442 17436
rect 11442 17380 11446 17436
rect 11382 17376 11446 17380
rect 11462 17436 11526 17440
rect 11462 17380 11466 17436
rect 11466 17380 11522 17436
rect 11522 17380 11526 17436
rect 11462 17376 11526 17380
rect 11542 17436 11606 17440
rect 11542 17380 11546 17436
rect 11546 17380 11602 17436
rect 11602 17380 11606 17436
rect 11542 17376 11606 17380
rect 18202 17436 18266 17440
rect 18202 17380 18206 17436
rect 18206 17380 18262 17436
rect 18262 17380 18266 17436
rect 18202 17376 18266 17380
rect 18282 17436 18346 17440
rect 18282 17380 18286 17436
rect 18286 17380 18342 17436
rect 18342 17380 18346 17436
rect 18282 17376 18346 17380
rect 18362 17436 18426 17440
rect 18362 17380 18366 17436
rect 18366 17380 18422 17436
rect 18422 17380 18426 17436
rect 18362 17376 18426 17380
rect 18442 17436 18506 17440
rect 18442 17380 18446 17436
rect 18446 17380 18502 17436
rect 18502 17380 18506 17436
rect 18442 17376 18506 17380
rect 7852 16892 7916 16896
rect 7852 16836 7856 16892
rect 7856 16836 7912 16892
rect 7912 16836 7916 16892
rect 7852 16832 7916 16836
rect 7932 16892 7996 16896
rect 7932 16836 7936 16892
rect 7936 16836 7992 16892
rect 7992 16836 7996 16892
rect 7932 16832 7996 16836
rect 8012 16892 8076 16896
rect 8012 16836 8016 16892
rect 8016 16836 8072 16892
rect 8072 16836 8076 16892
rect 8012 16832 8076 16836
rect 8092 16892 8156 16896
rect 8092 16836 8096 16892
rect 8096 16836 8152 16892
rect 8152 16836 8156 16892
rect 8092 16832 8156 16836
rect 14752 16892 14816 16896
rect 14752 16836 14756 16892
rect 14756 16836 14812 16892
rect 14812 16836 14816 16892
rect 14752 16832 14816 16836
rect 14832 16892 14896 16896
rect 14832 16836 14836 16892
rect 14836 16836 14892 16892
rect 14892 16836 14896 16892
rect 14832 16832 14896 16836
rect 14912 16892 14976 16896
rect 14912 16836 14916 16892
rect 14916 16836 14972 16892
rect 14972 16836 14976 16892
rect 14912 16832 14976 16836
rect 14992 16892 15056 16896
rect 14992 16836 14996 16892
rect 14996 16836 15052 16892
rect 15052 16836 15056 16892
rect 14992 16832 15056 16836
rect 4402 16348 4466 16352
rect 4402 16292 4406 16348
rect 4406 16292 4462 16348
rect 4462 16292 4466 16348
rect 4402 16288 4466 16292
rect 4482 16348 4546 16352
rect 4482 16292 4486 16348
rect 4486 16292 4542 16348
rect 4542 16292 4546 16348
rect 4482 16288 4546 16292
rect 4562 16348 4626 16352
rect 4562 16292 4566 16348
rect 4566 16292 4622 16348
rect 4622 16292 4626 16348
rect 4562 16288 4626 16292
rect 4642 16348 4706 16352
rect 4642 16292 4646 16348
rect 4646 16292 4702 16348
rect 4702 16292 4706 16348
rect 4642 16288 4706 16292
rect 11302 16348 11366 16352
rect 11302 16292 11306 16348
rect 11306 16292 11362 16348
rect 11362 16292 11366 16348
rect 11302 16288 11366 16292
rect 11382 16348 11446 16352
rect 11382 16292 11386 16348
rect 11386 16292 11442 16348
rect 11442 16292 11446 16348
rect 11382 16288 11446 16292
rect 11462 16348 11526 16352
rect 11462 16292 11466 16348
rect 11466 16292 11522 16348
rect 11522 16292 11526 16348
rect 11462 16288 11526 16292
rect 11542 16348 11606 16352
rect 11542 16292 11546 16348
rect 11546 16292 11602 16348
rect 11602 16292 11606 16348
rect 11542 16288 11606 16292
rect 18202 16348 18266 16352
rect 18202 16292 18206 16348
rect 18206 16292 18262 16348
rect 18262 16292 18266 16348
rect 18202 16288 18266 16292
rect 18282 16348 18346 16352
rect 18282 16292 18286 16348
rect 18286 16292 18342 16348
rect 18342 16292 18346 16348
rect 18282 16288 18346 16292
rect 18362 16348 18426 16352
rect 18362 16292 18366 16348
rect 18366 16292 18422 16348
rect 18422 16292 18426 16348
rect 18362 16288 18426 16292
rect 18442 16348 18506 16352
rect 18442 16292 18446 16348
rect 18446 16292 18502 16348
rect 18502 16292 18506 16348
rect 18442 16288 18506 16292
rect 7852 15804 7916 15808
rect 7852 15748 7856 15804
rect 7856 15748 7912 15804
rect 7912 15748 7916 15804
rect 7852 15744 7916 15748
rect 7932 15804 7996 15808
rect 7932 15748 7936 15804
rect 7936 15748 7992 15804
rect 7992 15748 7996 15804
rect 7932 15744 7996 15748
rect 8012 15804 8076 15808
rect 8012 15748 8016 15804
rect 8016 15748 8072 15804
rect 8072 15748 8076 15804
rect 8012 15744 8076 15748
rect 8092 15804 8156 15808
rect 8092 15748 8096 15804
rect 8096 15748 8152 15804
rect 8152 15748 8156 15804
rect 8092 15744 8156 15748
rect 14752 15804 14816 15808
rect 14752 15748 14756 15804
rect 14756 15748 14812 15804
rect 14812 15748 14816 15804
rect 14752 15744 14816 15748
rect 14832 15804 14896 15808
rect 14832 15748 14836 15804
rect 14836 15748 14892 15804
rect 14892 15748 14896 15804
rect 14832 15744 14896 15748
rect 14912 15804 14976 15808
rect 14912 15748 14916 15804
rect 14916 15748 14972 15804
rect 14972 15748 14976 15804
rect 14912 15744 14976 15748
rect 14992 15804 15056 15808
rect 14992 15748 14996 15804
rect 14996 15748 15052 15804
rect 15052 15748 15056 15804
rect 14992 15744 15056 15748
rect 4402 15260 4466 15264
rect 4402 15204 4406 15260
rect 4406 15204 4462 15260
rect 4462 15204 4466 15260
rect 4402 15200 4466 15204
rect 4482 15260 4546 15264
rect 4482 15204 4486 15260
rect 4486 15204 4542 15260
rect 4542 15204 4546 15260
rect 4482 15200 4546 15204
rect 4562 15260 4626 15264
rect 4562 15204 4566 15260
rect 4566 15204 4622 15260
rect 4622 15204 4626 15260
rect 4562 15200 4626 15204
rect 4642 15260 4706 15264
rect 4642 15204 4646 15260
rect 4646 15204 4702 15260
rect 4702 15204 4706 15260
rect 4642 15200 4706 15204
rect 11302 15260 11366 15264
rect 11302 15204 11306 15260
rect 11306 15204 11362 15260
rect 11362 15204 11366 15260
rect 11302 15200 11366 15204
rect 11382 15260 11446 15264
rect 11382 15204 11386 15260
rect 11386 15204 11442 15260
rect 11442 15204 11446 15260
rect 11382 15200 11446 15204
rect 11462 15260 11526 15264
rect 11462 15204 11466 15260
rect 11466 15204 11522 15260
rect 11522 15204 11526 15260
rect 11462 15200 11526 15204
rect 11542 15260 11606 15264
rect 11542 15204 11546 15260
rect 11546 15204 11602 15260
rect 11602 15204 11606 15260
rect 11542 15200 11606 15204
rect 18202 15260 18266 15264
rect 18202 15204 18206 15260
rect 18206 15204 18262 15260
rect 18262 15204 18266 15260
rect 18202 15200 18266 15204
rect 18282 15260 18346 15264
rect 18282 15204 18286 15260
rect 18286 15204 18342 15260
rect 18342 15204 18346 15260
rect 18282 15200 18346 15204
rect 18362 15260 18426 15264
rect 18362 15204 18366 15260
rect 18366 15204 18422 15260
rect 18422 15204 18426 15260
rect 18362 15200 18426 15204
rect 18442 15260 18506 15264
rect 18442 15204 18446 15260
rect 18446 15204 18502 15260
rect 18502 15204 18506 15260
rect 18442 15200 18506 15204
rect 7852 14716 7916 14720
rect 7852 14660 7856 14716
rect 7856 14660 7912 14716
rect 7912 14660 7916 14716
rect 7852 14656 7916 14660
rect 7932 14716 7996 14720
rect 7932 14660 7936 14716
rect 7936 14660 7992 14716
rect 7992 14660 7996 14716
rect 7932 14656 7996 14660
rect 8012 14716 8076 14720
rect 8012 14660 8016 14716
rect 8016 14660 8072 14716
rect 8072 14660 8076 14716
rect 8012 14656 8076 14660
rect 8092 14716 8156 14720
rect 8092 14660 8096 14716
rect 8096 14660 8152 14716
rect 8152 14660 8156 14716
rect 8092 14656 8156 14660
rect 14752 14716 14816 14720
rect 14752 14660 14756 14716
rect 14756 14660 14812 14716
rect 14812 14660 14816 14716
rect 14752 14656 14816 14660
rect 14832 14716 14896 14720
rect 14832 14660 14836 14716
rect 14836 14660 14892 14716
rect 14892 14660 14896 14716
rect 14832 14656 14896 14660
rect 14912 14716 14976 14720
rect 14912 14660 14916 14716
rect 14916 14660 14972 14716
rect 14972 14660 14976 14716
rect 14912 14656 14976 14660
rect 14992 14716 15056 14720
rect 14992 14660 14996 14716
rect 14996 14660 15052 14716
rect 15052 14660 15056 14716
rect 14992 14656 15056 14660
rect 4402 14172 4466 14176
rect 4402 14116 4406 14172
rect 4406 14116 4462 14172
rect 4462 14116 4466 14172
rect 4402 14112 4466 14116
rect 4482 14172 4546 14176
rect 4482 14116 4486 14172
rect 4486 14116 4542 14172
rect 4542 14116 4546 14172
rect 4482 14112 4546 14116
rect 4562 14172 4626 14176
rect 4562 14116 4566 14172
rect 4566 14116 4622 14172
rect 4622 14116 4626 14172
rect 4562 14112 4626 14116
rect 4642 14172 4706 14176
rect 4642 14116 4646 14172
rect 4646 14116 4702 14172
rect 4702 14116 4706 14172
rect 4642 14112 4706 14116
rect 11302 14172 11366 14176
rect 11302 14116 11306 14172
rect 11306 14116 11362 14172
rect 11362 14116 11366 14172
rect 11302 14112 11366 14116
rect 11382 14172 11446 14176
rect 11382 14116 11386 14172
rect 11386 14116 11442 14172
rect 11442 14116 11446 14172
rect 11382 14112 11446 14116
rect 11462 14172 11526 14176
rect 11462 14116 11466 14172
rect 11466 14116 11522 14172
rect 11522 14116 11526 14172
rect 11462 14112 11526 14116
rect 11542 14172 11606 14176
rect 11542 14116 11546 14172
rect 11546 14116 11602 14172
rect 11602 14116 11606 14172
rect 11542 14112 11606 14116
rect 18202 14172 18266 14176
rect 18202 14116 18206 14172
rect 18206 14116 18262 14172
rect 18262 14116 18266 14172
rect 18202 14112 18266 14116
rect 18282 14172 18346 14176
rect 18282 14116 18286 14172
rect 18286 14116 18342 14172
rect 18342 14116 18346 14172
rect 18282 14112 18346 14116
rect 18362 14172 18426 14176
rect 18362 14116 18366 14172
rect 18366 14116 18422 14172
rect 18422 14116 18426 14172
rect 18362 14112 18426 14116
rect 18442 14172 18506 14176
rect 18442 14116 18446 14172
rect 18446 14116 18502 14172
rect 18502 14116 18506 14172
rect 18442 14112 18506 14116
rect 7852 13628 7916 13632
rect 7852 13572 7856 13628
rect 7856 13572 7912 13628
rect 7912 13572 7916 13628
rect 7852 13568 7916 13572
rect 7932 13628 7996 13632
rect 7932 13572 7936 13628
rect 7936 13572 7992 13628
rect 7992 13572 7996 13628
rect 7932 13568 7996 13572
rect 8012 13628 8076 13632
rect 8012 13572 8016 13628
rect 8016 13572 8072 13628
rect 8072 13572 8076 13628
rect 8012 13568 8076 13572
rect 8092 13628 8156 13632
rect 8092 13572 8096 13628
rect 8096 13572 8152 13628
rect 8152 13572 8156 13628
rect 8092 13568 8156 13572
rect 14752 13628 14816 13632
rect 14752 13572 14756 13628
rect 14756 13572 14812 13628
rect 14812 13572 14816 13628
rect 14752 13568 14816 13572
rect 14832 13628 14896 13632
rect 14832 13572 14836 13628
rect 14836 13572 14892 13628
rect 14892 13572 14896 13628
rect 14832 13568 14896 13572
rect 14912 13628 14976 13632
rect 14912 13572 14916 13628
rect 14916 13572 14972 13628
rect 14972 13572 14976 13628
rect 14912 13568 14976 13572
rect 14992 13628 15056 13632
rect 14992 13572 14996 13628
rect 14996 13572 15052 13628
rect 15052 13572 15056 13628
rect 14992 13568 15056 13572
rect 4402 13084 4466 13088
rect 4402 13028 4406 13084
rect 4406 13028 4462 13084
rect 4462 13028 4466 13084
rect 4402 13024 4466 13028
rect 4482 13084 4546 13088
rect 4482 13028 4486 13084
rect 4486 13028 4542 13084
rect 4542 13028 4546 13084
rect 4482 13024 4546 13028
rect 4562 13084 4626 13088
rect 4562 13028 4566 13084
rect 4566 13028 4622 13084
rect 4622 13028 4626 13084
rect 4562 13024 4626 13028
rect 4642 13084 4706 13088
rect 4642 13028 4646 13084
rect 4646 13028 4702 13084
rect 4702 13028 4706 13084
rect 4642 13024 4706 13028
rect 11302 13084 11366 13088
rect 11302 13028 11306 13084
rect 11306 13028 11362 13084
rect 11362 13028 11366 13084
rect 11302 13024 11366 13028
rect 11382 13084 11446 13088
rect 11382 13028 11386 13084
rect 11386 13028 11442 13084
rect 11442 13028 11446 13084
rect 11382 13024 11446 13028
rect 11462 13084 11526 13088
rect 11462 13028 11466 13084
rect 11466 13028 11522 13084
rect 11522 13028 11526 13084
rect 11462 13024 11526 13028
rect 11542 13084 11606 13088
rect 11542 13028 11546 13084
rect 11546 13028 11602 13084
rect 11602 13028 11606 13084
rect 11542 13024 11606 13028
rect 18202 13084 18266 13088
rect 18202 13028 18206 13084
rect 18206 13028 18262 13084
rect 18262 13028 18266 13084
rect 18202 13024 18266 13028
rect 18282 13084 18346 13088
rect 18282 13028 18286 13084
rect 18286 13028 18342 13084
rect 18342 13028 18346 13084
rect 18282 13024 18346 13028
rect 18362 13084 18426 13088
rect 18362 13028 18366 13084
rect 18366 13028 18422 13084
rect 18422 13028 18426 13084
rect 18362 13024 18426 13028
rect 18442 13084 18506 13088
rect 18442 13028 18446 13084
rect 18446 13028 18502 13084
rect 18502 13028 18506 13084
rect 18442 13024 18506 13028
rect 7852 12540 7916 12544
rect 7852 12484 7856 12540
rect 7856 12484 7912 12540
rect 7912 12484 7916 12540
rect 7852 12480 7916 12484
rect 7932 12540 7996 12544
rect 7932 12484 7936 12540
rect 7936 12484 7992 12540
rect 7992 12484 7996 12540
rect 7932 12480 7996 12484
rect 8012 12540 8076 12544
rect 8012 12484 8016 12540
rect 8016 12484 8072 12540
rect 8072 12484 8076 12540
rect 8012 12480 8076 12484
rect 8092 12540 8156 12544
rect 8092 12484 8096 12540
rect 8096 12484 8152 12540
rect 8152 12484 8156 12540
rect 8092 12480 8156 12484
rect 14752 12540 14816 12544
rect 14752 12484 14756 12540
rect 14756 12484 14812 12540
rect 14812 12484 14816 12540
rect 14752 12480 14816 12484
rect 14832 12540 14896 12544
rect 14832 12484 14836 12540
rect 14836 12484 14892 12540
rect 14892 12484 14896 12540
rect 14832 12480 14896 12484
rect 14912 12540 14976 12544
rect 14912 12484 14916 12540
rect 14916 12484 14972 12540
rect 14972 12484 14976 12540
rect 14912 12480 14976 12484
rect 14992 12540 15056 12544
rect 14992 12484 14996 12540
rect 14996 12484 15052 12540
rect 15052 12484 15056 12540
rect 14992 12480 15056 12484
rect 4402 11996 4466 12000
rect 4402 11940 4406 11996
rect 4406 11940 4462 11996
rect 4462 11940 4466 11996
rect 4402 11936 4466 11940
rect 4482 11996 4546 12000
rect 4482 11940 4486 11996
rect 4486 11940 4542 11996
rect 4542 11940 4546 11996
rect 4482 11936 4546 11940
rect 4562 11996 4626 12000
rect 4562 11940 4566 11996
rect 4566 11940 4622 11996
rect 4622 11940 4626 11996
rect 4562 11936 4626 11940
rect 4642 11996 4706 12000
rect 4642 11940 4646 11996
rect 4646 11940 4702 11996
rect 4702 11940 4706 11996
rect 4642 11936 4706 11940
rect 11302 11996 11366 12000
rect 11302 11940 11306 11996
rect 11306 11940 11362 11996
rect 11362 11940 11366 11996
rect 11302 11936 11366 11940
rect 11382 11996 11446 12000
rect 11382 11940 11386 11996
rect 11386 11940 11442 11996
rect 11442 11940 11446 11996
rect 11382 11936 11446 11940
rect 11462 11996 11526 12000
rect 11462 11940 11466 11996
rect 11466 11940 11522 11996
rect 11522 11940 11526 11996
rect 11462 11936 11526 11940
rect 11542 11996 11606 12000
rect 11542 11940 11546 11996
rect 11546 11940 11602 11996
rect 11602 11940 11606 11996
rect 11542 11936 11606 11940
rect 18202 11996 18266 12000
rect 18202 11940 18206 11996
rect 18206 11940 18262 11996
rect 18262 11940 18266 11996
rect 18202 11936 18266 11940
rect 18282 11996 18346 12000
rect 18282 11940 18286 11996
rect 18286 11940 18342 11996
rect 18342 11940 18346 11996
rect 18282 11936 18346 11940
rect 18362 11996 18426 12000
rect 18362 11940 18366 11996
rect 18366 11940 18422 11996
rect 18422 11940 18426 11996
rect 18362 11936 18426 11940
rect 18442 11996 18506 12000
rect 18442 11940 18446 11996
rect 18446 11940 18502 11996
rect 18502 11940 18506 11996
rect 18442 11936 18506 11940
rect 7852 11452 7916 11456
rect 7852 11396 7856 11452
rect 7856 11396 7912 11452
rect 7912 11396 7916 11452
rect 7852 11392 7916 11396
rect 7932 11452 7996 11456
rect 7932 11396 7936 11452
rect 7936 11396 7992 11452
rect 7992 11396 7996 11452
rect 7932 11392 7996 11396
rect 8012 11452 8076 11456
rect 8012 11396 8016 11452
rect 8016 11396 8072 11452
rect 8072 11396 8076 11452
rect 8012 11392 8076 11396
rect 8092 11452 8156 11456
rect 8092 11396 8096 11452
rect 8096 11396 8152 11452
rect 8152 11396 8156 11452
rect 8092 11392 8156 11396
rect 14752 11452 14816 11456
rect 14752 11396 14756 11452
rect 14756 11396 14812 11452
rect 14812 11396 14816 11452
rect 14752 11392 14816 11396
rect 14832 11452 14896 11456
rect 14832 11396 14836 11452
rect 14836 11396 14892 11452
rect 14892 11396 14896 11452
rect 14832 11392 14896 11396
rect 14912 11452 14976 11456
rect 14912 11396 14916 11452
rect 14916 11396 14972 11452
rect 14972 11396 14976 11452
rect 14912 11392 14976 11396
rect 14992 11452 15056 11456
rect 14992 11396 14996 11452
rect 14996 11396 15052 11452
rect 15052 11396 15056 11452
rect 14992 11392 15056 11396
rect 4402 10908 4466 10912
rect 4402 10852 4406 10908
rect 4406 10852 4462 10908
rect 4462 10852 4466 10908
rect 4402 10848 4466 10852
rect 4482 10908 4546 10912
rect 4482 10852 4486 10908
rect 4486 10852 4542 10908
rect 4542 10852 4546 10908
rect 4482 10848 4546 10852
rect 4562 10908 4626 10912
rect 4562 10852 4566 10908
rect 4566 10852 4622 10908
rect 4622 10852 4626 10908
rect 4562 10848 4626 10852
rect 4642 10908 4706 10912
rect 4642 10852 4646 10908
rect 4646 10852 4702 10908
rect 4702 10852 4706 10908
rect 4642 10848 4706 10852
rect 11302 10908 11366 10912
rect 11302 10852 11306 10908
rect 11306 10852 11362 10908
rect 11362 10852 11366 10908
rect 11302 10848 11366 10852
rect 11382 10908 11446 10912
rect 11382 10852 11386 10908
rect 11386 10852 11442 10908
rect 11442 10852 11446 10908
rect 11382 10848 11446 10852
rect 11462 10908 11526 10912
rect 11462 10852 11466 10908
rect 11466 10852 11522 10908
rect 11522 10852 11526 10908
rect 11462 10848 11526 10852
rect 11542 10908 11606 10912
rect 11542 10852 11546 10908
rect 11546 10852 11602 10908
rect 11602 10852 11606 10908
rect 11542 10848 11606 10852
rect 18202 10908 18266 10912
rect 18202 10852 18206 10908
rect 18206 10852 18262 10908
rect 18262 10852 18266 10908
rect 18202 10848 18266 10852
rect 18282 10908 18346 10912
rect 18282 10852 18286 10908
rect 18286 10852 18342 10908
rect 18342 10852 18346 10908
rect 18282 10848 18346 10852
rect 18362 10908 18426 10912
rect 18362 10852 18366 10908
rect 18366 10852 18422 10908
rect 18422 10852 18426 10908
rect 18362 10848 18426 10852
rect 18442 10908 18506 10912
rect 18442 10852 18446 10908
rect 18446 10852 18502 10908
rect 18502 10852 18506 10908
rect 18442 10848 18506 10852
rect 7852 10364 7916 10368
rect 7852 10308 7856 10364
rect 7856 10308 7912 10364
rect 7912 10308 7916 10364
rect 7852 10304 7916 10308
rect 7932 10364 7996 10368
rect 7932 10308 7936 10364
rect 7936 10308 7992 10364
rect 7992 10308 7996 10364
rect 7932 10304 7996 10308
rect 8012 10364 8076 10368
rect 8012 10308 8016 10364
rect 8016 10308 8072 10364
rect 8072 10308 8076 10364
rect 8012 10304 8076 10308
rect 8092 10364 8156 10368
rect 8092 10308 8096 10364
rect 8096 10308 8152 10364
rect 8152 10308 8156 10364
rect 8092 10304 8156 10308
rect 14752 10364 14816 10368
rect 14752 10308 14756 10364
rect 14756 10308 14812 10364
rect 14812 10308 14816 10364
rect 14752 10304 14816 10308
rect 14832 10364 14896 10368
rect 14832 10308 14836 10364
rect 14836 10308 14892 10364
rect 14892 10308 14896 10364
rect 14832 10304 14896 10308
rect 14912 10364 14976 10368
rect 14912 10308 14916 10364
rect 14916 10308 14972 10364
rect 14972 10308 14976 10364
rect 14912 10304 14976 10308
rect 14992 10364 15056 10368
rect 14992 10308 14996 10364
rect 14996 10308 15052 10364
rect 15052 10308 15056 10364
rect 14992 10304 15056 10308
rect 4402 9820 4466 9824
rect 4402 9764 4406 9820
rect 4406 9764 4462 9820
rect 4462 9764 4466 9820
rect 4402 9760 4466 9764
rect 4482 9820 4546 9824
rect 4482 9764 4486 9820
rect 4486 9764 4542 9820
rect 4542 9764 4546 9820
rect 4482 9760 4546 9764
rect 4562 9820 4626 9824
rect 4562 9764 4566 9820
rect 4566 9764 4622 9820
rect 4622 9764 4626 9820
rect 4562 9760 4626 9764
rect 4642 9820 4706 9824
rect 4642 9764 4646 9820
rect 4646 9764 4702 9820
rect 4702 9764 4706 9820
rect 4642 9760 4706 9764
rect 11302 9820 11366 9824
rect 11302 9764 11306 9820
rect 11306 9764 11362 9820
rect 11362 9764 11366 9820
rect 11302 9760 11366 9764
rect 11382 9820 11446 9824
rect 11382 9764 11386 9820
rect 11386 9764 11442 9820
rect 11442 9764 11446 9820
rect 11382 9760 11446 9764
rect 11462 9820 11526 9824
rect 11462 9764 11466 9820
rect 11466 9764 11522 9820
rect 11522 9764 11526 9820
rect 11462 9760 11526 9764
rect 11542 9820 11606 9824
rect 11542 9764 11546 9820
rect 11546 9764 11602 9820
rect 11602 9764 11606 9820
rect 11542 9760 11606 9764
rect 18202 9820 18266 9824
rect 18202 9764 18206 9820
rect 18206 9764 18262 9820
rect 18262 9764 18266 9820
rect 18202 9760 18266 9764
rect 18282 9820 18346 9824
rect 18282 9764 18286 9820
rect 18286 9764 18342 9820
rect 18342 9764 18346 9820
rect 18282 9760 18346 9764
rect 18362 9820 18426 9824
rect 18362 9764 18366 9820
rect 18366 9764 18422 9820
rect 18422 9764 18426 9820
rect 18362 9760 18426 9764
rect 18442 9820 18506 9824
rect 18442 9764 18446 9820
rect 18446 9764 18502 9820
rect 18502 9764 18506 9820
rect 18442 9760 18506 9764
rect 7852 9276 7916 9280
rect 7852 9220 7856 9276
rect 7856 9220 7912 9276
rect 7912 9220 7916 9276
rect 7852 9216 7916 9220
rect 7932 9276 7996 9280
rect 7932 9220 7936 9276
rect 7936 9220 7992 9276
rect 7992 9220 7996 9276
rect 7932 9216 7996 9220
rect 8012 9276 8076 9280
rect 8012 9220 8016 9276
rect 8016 9220 8072 9276
rect 8072 9220 8076 9276
rect 8012 9216 8076 9220
rect 8092 9276 8156 9280
rect 8092 9220 8096 9276
rect 8096 9220 8152 9276
rect 8152 9220 8156 9276
rect 8092 9216 8156 9220
rect 14752 9276 14816 9280
rect 14752 9220 14756 9276
rect 14756 9220 14812 9276
rect 14812 9220 14816 9276
rect 14752 9216 14816 9220
rect 14832 9276 14896 9280
rect 14832 9220 14836 9276
rect 14836 9220 14892 9276
rect 14892 9220 14896 9276
rect 14832 9216 14896 9220
rect 14912 9276 14976 9280
rect 14912 9220 14916 9276
rect 14916 9220 14972 9276
rect 14972 9220 14976 9276
rect 14912 9216 14976 9220
rect 14992 9276 15056 9280
rect 14992 9220 14996 9276
rect 14996 9220 15052 9276
rect 15052 9220 15056 9276
rect 14992 9216 15056 9220
rect 4402 8732 4466 8736
rect 4402 8676 4406 8732
rect 4406 8676 4462 8732
rect 4462 8676 4466 8732
rect 4402 8672 4466 8676
rect 4482 8732 4546 8736
rect 4482 8676 4486 8732
rect 4486 8676 4542 8732
rect 4542 8676 4546 8732
rect 4482 8672 4546 8676
rect 4562 8732 4626 8736
rect 4562 8676 4566 8732
rect 4566 8676 4622 8732
rect 4622 8676 4626 8732
rect 4562 8672 4626 8676
rect 4642 8732 4706 8736
rect 4642 8676 4646 8732
rect 4646 8676 4702 8732
rect 4702 8676 4706 8732
rect 4642 8672 4706 8676
rect 11302 8732 11366 8736
rect 11302 8676 11306 8732
rect 11306 8676 11362 8732
rect 11362 8676 11366 8732
rect 11302 8672 11366 8676
rect 11382 8732 11446 8736
rect 11382 8676 11386 8732
rect 11386 8676 11442 8732
rect 11442 8676 11446 8732
rect 11382 8672 11446 8676
rect 11462 8732 11526 8736
rect 11462 8676 11466 8732
rect 11466 8676 11522 8732
rect 11522 8676 11526 8732
rect 11462 8672 11526 8676
rect 11542 8732 11606 8736
rect 11542 8676 11546 8732
rect 11546 8676 11602 8732
rect 11602 8676 11606 8732
rect 11542 8672 11606 8676
rect 18202 8732 18266 8736
rect 18202 8676 18206 8732
rect 18206 8676 18262 8732
rect 18262 8676 18266 8732
rect 18202 8672 18266 8676
rect 18282 8732 18346 8736
rect 18282 8676 18286 8732
rect 18286 8676 18342 8732
rect 18342 8676 18346 8732
rect 18282 8672 18346 8676
rect 18362 8732 18426 8736
rect 18362 8676 18366 8732
rect 18366 8676 18422 8732
rect 18422 8676 18426 8732
rect 18362 8672 18426 8676
rect 18442 8732 18506 8736
rect 18442 8676 18446 8732
rect 18446 8676 18502 8732
rect 18502 8676 18506 8732
rect 18442 8672 18506 8676
rect 7852 8188 7916 8192
rect 7852 8132 7856 8188
rect 7856 8132 7912 8188
rect 7912 8132 7916 8188
rect 7852 8128 7916 8132
rect 7932 8188 7996 8192
rect 7932 8132 7936 8188
rect 7936 8132 7992 8188
rect 7992 8132 7996 8188
rect 7932 8128 7996 8132
rect 8012 8188 8076 8192
rect 8012 8132 8016 8188
rect 8016 8132 8072 8188
rect 8072 8132 8076 8188
rect 8012 8128 8076 8132
rect 8092 8188 8156 8192
rect 8092 8132 8096 8188
rect 8096 8132 8152 8188
rect 8152 8132 8156 8188
rect 8092 8128 8156 8132
rect 14752 8188 14816 8192
rect 14752 8132 14756 8188
rect 14756 8132 14812 8188
rect 14812 8132 14816 8188
rect 14752 8128 14816 8132
rect 14832 8188 14896 8192
rect 14832 8132 14836 8188
rect 14836 8132 14892 8188
rect 14892 8132 14896 8188
rect 14832 8128 14896 8132
rect 14912 8188 14976 8192
rect 14912 8132 14916 8188
rect 14916 8132 14972 8188
rect 14972 8132 14976 8188
rect 14912 8128 14976 8132
rect 14992 8188 15056 8192
rect 14992 8132 14996 8188
rect 14996 8132 15052 8188
rect 15052 8132 15056 8188
rect 14992 8128 15056 8132
rect 4402 7644 4466 7648
rect 4402 7588 4406 7644
rect 4406 7588 4462 7644
rect 4462 7588 4466 7644
rect 4402 7584 4466 7588
rect 4482 7644 4546 7648
rect 4482 7588 4486 7644
rect 4486 7588 4542 7644
rect 4542 7588 4546 7644
rect 4482 7584 4546 7588
rect 4562 7644 4626 7648
rect 4562 7588 4566 7644
rect 4566 7588 4622 7644
rect 4622 7588 4626 7644
rect 4562 7584 4626 7588
rect 4642 7644 4706 7648
rect 4642 7588 4646 7644
rect 4646 7588 4702 7644
rect 4702 7588 4706 7644
rect 4642 7584 4706 7588
rect 11302 7644 11366 7648
rect 11302 7588 11306 7644
rect 11306 7588 11362 7644
rect 11362 7588 11366 7644
rect 11302 7584 11366 7588
rect 11382 7644 11446 7648
rect 11382 7588 11386 7644
rect 11386 7588 11442 7644
rect 11442 7588 11446 7644
rect 11382 7584 11446 7588
rect 11462 7644 11526 7648
rect 11462 7588 11466 7644
rect 11466 7588 11522 7644
rect 11522 7588 11526 7644
rect 11462 7584 11526 7588
rect 11542 7644 11606 7648
rect 11542 7588 11546 7644
rect 11546 7588 11602 7644
rect 11602 7588 11606 7644
rect 11542 7584 11606 7588
rect 18202 7644 18266 7648
rect 18202 7588 18206 7644
rect 18206 7588 18262 7644
rect 18262 7588 18266 7644
rect 18202 7584 18266 7588
rect 18282 7644 18346 7648
rect 18282 7588 18286 7644
rect 18286 7588 18342 7644
rect 18342 7588 18346 7644
rect 18282 7584 18346 7588
rect 18362 7644 18426 7648
rect 18362 7588 18366 7644
rect 18366 7588 18422 7644
rect 18422 7588 18426 7644
rect 18362 7584 18426 7588
rect 18442 7644 18506 7648
rect 18442 7588 18446 7644
rect 18446 7588 18502 7644
rect 18502 7588 18506 7644
rect 18442 7584 18506 7588
rect 7852 7100 7916 7104
rect 7852 7044 7856 7100
rect 7856 7044 7912 7100
rect 7912 7044 7916 7100
rect 7852 7040 7916 7044
rect 7932 7100 7996 7104
rect 7932 7044 7936 7100
rect 7936 7044 7992 7100
rect 7992 7044 7996 7100
rect 7932 7040 7996 7044
rect 8012 7100 8076 7104
rect 8012 7044 8016 7100
rect 8016 7044 8072 7100
rect 8072 7044 8076 7100
rect 8012 7040 8076 7044
rect 8092 7100 8156 7104
rect 8092 7044 8096 7100
rect 8096 7044 8152 7100
rect 8152 7044 8156 7100
rect 8092 7040 8156 7044
rect 14752 7100 14816 7104
rect 14752 7044 14756 7100
rect 14756 7044 14812 7100
rect 14812 7044 14816 7100
rect 14752 7040 14816 7044
rect 14832 7100 14896 7104
rect 14832 7044 14836 7100
rect 14836 7044 14892 7100
rect 14892 7044 14896 7100
rect 14832 7040 14896 7044
rect 14912 7100 14976 7104
rect 14912 7044 14916 7100
rect 14916 7044 14972 7100
rect 14972 7044 14976 7100
rect 14912 7040 14976 7044
rect 14992 7100 15056 7104
rect 14992 7044 14996 7100
rect 14996 7044 15052 7100
rect 15052 7044 15056 7100
rect 14992 7040 15056 7044
rect 4402 6556 4466 6560
rect 4402 6500 4406 6556
rect 4406 6500 4462 6556
rect 4462 6500 4466 6556
rect 4402 6496 4466 6500
rect 4482 6556 4546 6560
rect 4482 6500 4486 6556
rect 4486 6500 4542 6556
rect 4542 6500 4546 6556
rect 4482 6496 4546 6500
rect 4562 6556 4626 6560
rect 4562 6500 4566 6556
rect 4566 6500 4622 6556
rect 4622 6500 4626 6556
rect 4562 6496 4626 6500
rect 4642 6556 4706 6560
rect 4642 6500 4646 6556
rect 4646 6500 4702 6556
rect 4702 6500 4706 6556
rect 4642 6496 4706 6500
rect 11302 6556 11366 6560
rect 11302 6500 11306 6556
rect 11306 6500 11362 6556
rect 11362 6500 11366 6556
rect 11302 6496 11366 6500
rect 11382 6556 11446 6560
rect 11382 6500 11386 6556
rect 11386 6500 11442 6556
rect 11442 6500 11446 6556
rect 11382 6496 11446 6500
rect 11462 6556 11526 6560
rect 11462 6500 11466 6556
rect 11466 6500 11522 6556
rect 11522 6500 11526 6556
rect 11462 6496 11526 6500
rect 11542 6556 11606 6560
rect 11542 6500 11546 6556
rect 11546 6500 11602 6556
rect 11602 6500 11606 6556
rect 11542 6496 11606 6500
rect 18202 6556 18266 6560
rect 18202 6500 18206 6556
rect 18206 6500 18262 6556
rect 18262 6500 18266 6556
rect 18202 6496 18266 6500
rect 18282 6556 18346 6560
rect 18282 6500 18286 6556
rect 18286 6500 18342 6556
rect 18342 6500 18346 6556
rect 18282 6496 18346 6500
rect 18362 6556 18426 6560
rect 18362 6500 18366 6556
rect 18366 6500 18422 6556
rect 18422 6500 18426 6556
rect 18362 6496 18426 6500
rect 18442 6556 18506 6560
rect 18442 6500 18446 6556
rect 18446 6500 18502 6556
rect 18502 6500 18506 6556
rect 18442 6496 18506 6500
rect 7852 6012 7916 6016
rect 7852 5956 7856 6012
rect 7856 5956 7912 6012
rect 7912 5956 7916 6012
rect 7852 5952 7916 5956
rect 7932 6012 7996 6016
rect 7932 5956 7936 6012
rect 7936 5956 7992 6012
rect 7992 5956 7996 6012
rect 7932 5952 7996 5956
rect 8012 6012 8076 6016
rect 8012 5956 8016 6012
rect 8016 5956 8072 6012
rect 8072 5956 8076 6012
rect 8012 5952 8076 5956
rect 8092 6012 8156 6016
rect 8092 5956 8096 6012
rect 8096 5956 8152 6012
rect 8152 5956 8156 6012
rect 8092 5952 8156 5956
rect 14752 6012 14816 6016
rect 14752 5956 14756 6012
rect 14756 5956 14812 6012
rect 14812 5956 14816 6012
rect 14752 5952 14816 5956
rect 14832 6012 14896 6016
rect 14832 5956 14836 6012
rect 14836 5956 14892 6012
rect 14892 5956 14896 6012
rect 14832 5952 14896 5956
rect 14912 6012 14976 6016
rect 14912 5956 14916 6012
rect 14916 5956 14972 6012
rect 14972 5956 14976 6012
rect 14912 5952 14976 5956
rect 14992 6012 15056 6016
rect 14992 5956 14996 6012
rect 14996 5956 15052 6012
rect 15052 5956 15056 6012
rect 14992 5952 15056 5956
rect 4402 5468 4466 5472
rect 4402 5412 4406 5468
rect 4406 5412 4462 5468
rect 4462 5412 4466 5468
rect 4402 5408 4466 5412
rect 4482 5468 4546 5472
rect 4482 5412 4486 5468
rect 4486 5412 4542 5468
rect 4542 5412 4546 5468
rect 4482 5408 4546 5412
rect 4562 5468 4626 5472
rect 4562 5412 4566 5468
rect 4566 5412 4622 5468
rect 4622 5412 4626 5468
rect 4562 5408 4626 5412
rect 4642 5468 4706 5472
rect 4642 5412 4646 5468
rect 4646 5412 4702 5468
rect 4702 5412 4706 5468
rect 4642 5408 4706 5412
rect 11302 5468 11366 5472
rect 11302 5412 11306 5468
rect 11306 5412 11362 5468
rect 11362 5412 11366 5468
rect 11302 5408 11366 5412
rect 11382 5468 11446 5472
rect 11382 5412 11386 5468
rect 11386 5412 11442 5468
rect 11442 5412 11446 5468
rect 11382 5408 11446 5412
rect 11462 5468 11526 5472
rect 11462 5412 11466 5468
rect 11466 5412 11522 5468
rect 11522 5412 11526 5468
rect 11462 5408 11526 5412
rect 11542 5468 11606 5472
rect 11542 5412 11546 5468
rect 11546 5412 11602 5468
rect 11602 5412 11606 5468
rect 11542 5408 11606 5412
rect 18202 5468 18266 5472
rect 18202 5412 18206 5468
rect 18206 5412 18262 5468
rect 18262 5412 18266 5468
rect 18202 5408 18266 5412
rect 18282 5468 18346 5472
rect 18282 5412 18286 5468
rect 18286 5412 18342 5468
rect 18342 5412 18346 5468
rect 18282 5408 18346 5412
rect 18362 5468 18426 5472
rect 18362 5412 18366 5468
rect 18366 5412 18422 5468
rect 18422 5412 18426 5468
rect 18362 5408 18426 5412
rect 18442 5468 18506 5472
rect 18442 5412 18446 5468
rect 18446 5412 18502 5468
rect 18502 5412 18506 5468
rect 18442 5408 18506 5412
rect 7852 4924 7916 4928
rect 7852 4868 7856 4924
rect 7856 4868 7912 4924
rect 7912 4868 7916 4924
rect 7852 4864 7916 4868
rect 7932 4924 7996 4928
rect 7932 4868 7936 4924
rect 7936 4868 7992 4924
rect 7992 4868 7996 4924
rect 7932 4864 7996 4868
rect 8012 4924 8076 4928
rect 8012 4868 8016 4924
rect 8016 4868 8072 4924
rect 8072 4868 8076 4924
rect 8012 4864 8076 4868
rect 8092 4924 8156 4928
rect 8092 4868 8096 4924
rect 8096 4868 8152 4924
rect 8152 4868 8156 4924
rect 8092 4864 8156 4868
rect 14752 4924 14816 4928
rect 14752 4868 14756 4924
rect 14756 4868 14812 4924
rect 14812 4868 14816 4924
rect 14752 4864 14816 4868
rect 14832 4924 14896 4928
rect 14832 4868 14836 4924
rect 14836 4868 14892 4924
rect 14892 4868 14896 4924
rect 14832 4864 14896 4868
rect 14912 4924 14976 4928
rect 14912 4868 14916 4924
rect 14916 4868 14972 4924
rect 14972 4868 14976 4924
rect 14912 4864 14976 4868
rect 14992 4924 15056 4928
rect 14992 4868 14996 4924
rect 14996 4868 15052 4924
rect 15052 4868 15056 4924
rect 14992 4864 15056 4868
rect 4402 4380 4466 4384
rect 4402 4324 4406 4380
rect 4406 4324 4462 4380
rect 4462 4324 4466 4380
rect 4402 4320 4466 4324
rect 4482 4380 4546 4384
rect 4482 4324 4486 4380
rect 4486 4324 4542 4380
rect 4542 4324 4546 4380
rect 4482 4320 4546 4324
rect 4562 4380 4626 4384
rect 4562 4324 4566 4380
rect 4566 4324 4622 4380
rect 4622 4324 4626 4380
rect 4562 4320 4626 4324
rect 4642 4380 4706 4384
rect 4642 4324 4646 4380
rect 4646 4324 4702 4380
rect 4702 4324 4706 4380
rect 4642 4320 4706 4324
rect 11302 4380 11366 4384
rect 11302 4324 11306 4380
rect 11306 4324 11362 4380
rect 11362 4324 11366 4380
rect 11302 4320 11366 4324
rect 11382 4380 11446 4384
rect 11382 4324 11386 4380
rect 11386 4324 11442 4380
rect 11442 4324 11446 4380
rect 11382 4320 11446 4324
rect 11462 4380 11526 4384
rect 11462 4324 11466 4380
rect 11466 4324 11522 4380
rect 11522 4324 11526 4380
rect 11462 4320 11526 4324
rect 11542 4380 11606 4384
rect 11542 4324 11546 4380
rect 11546 4324 11602 4380
rect 11602 4324 11606 4380
rect 11542 4320 11606 4324
rect 18202 4380 18266 4384
rect 18202 4324 18206 4380
rect 18206 4324 18262 4380
rect 18262 4324 18266 4380
rect 18202 4320 18266 4324
rect 18282 4380 18346 4384
rect 18282 4324 18286 4380
rect 18286 4324 18342 4380
rect 18342 4324 18346 4380
rect 18282 4320 18346 4324
rect 18362 4380 18426 4384
rect 18362 4324 18366 4380
rect 18366 4324 18422 4380
rect 18422 4324 18426 4380
rect 18362 4320 18426 4324
rect 18442 4380 18506 4384
rect 18442 4324 18446 4380
rect 18446 4324 18502 4380
rect 18502 4324 18506 4380
rect 18442 4320 18506 4324
rect 7852 3836 7916 3840
rect 7852 3780 7856 3836
rect 7856 3780 7912 3836
rect 7912 3780 7916 3836
rect 7852 3776 7916 3780
rect 7932 3836 7996 3840
rect 7932 3780 7936 3836
rect 7936 3780 7992 3836
rect 7992 3780 7996 3836
rect 7932 3776 7996 3780
rect 8012 3836 8076 3840
rect 8012 3780 8016 3836
rect 8016 3780 8072 3836
rect 8072 3780 8076 3836
rect 8012 3776 8076 3780
rect 8092 3836 8156 3840
rect 8092 3780 8096 3836
rect 8096 3780 8152 3836
rect 8152 3780 8156 3836
rect 8092 3776 8156 3780
rect 14752 3836 14816 3840
rect 14752 3780 14756 3836
rect 14756 3780 14812 3836
rect 14812 3780 14816 3836
rect 14752 3776 14816 3780
rect 14832 3836 14896 3840
rect 14832 3780 14836 3836
rect 14836 3780 14892 3836
rect 14892 3780 14896 3836
rect 14832 3776 14896 3780
rect 14912 3836 14976 3840
rect 14912 3780 14916 3836
rect 14916 3780 14972 3836
rect 14972 3780 14976 3836
rect 14912 3776 14976 3780
rect 14992 3836 15056 3840
rect 14992 3780 14996 3836
rect 14996 3780 15052 3836
rect 15052 3780 15056 3836
rect 14992 3776 15056 3780
rect 4402 3292 4466 3296
rect 4402 3236 4406 3292
rect 4406 3236 4462 3292
rect 4462 3236 4466 3292
rect 4402 3232 4466 3236
rect 4482 3292 4546 3296
rect 4482 3236 4486 3292
rect 4486 3236 4542 3292
rect 4542 3236 4546 3292
rect 4482 3232 4546 3236
rect 4562 3292 4626 3296
rect 4562 3236 4566 3292
rect 4566 3236 4622 3292
rect 4622 3236 4626 3292
rect 4562 3232 4626 3236
rect 4642 3292 4706 3296
rect 4642 3236 4646 3292
rect 4646 3236 4702 3292
rect 4702 3236 4706 3292
rect 4642 3232 4706 3236
rect 11302 3292 11366 3296
rect 11302 3236 11306 3292
rect 11306 3236 11362 3292
rect 11362 3236 11366 3292
rect 11302 3232 11366 3236
rect 11382 3292 11446 3296
rect 11382 3236 11386 3292
rect 11386 3236 11442 3292
rect 11442 3236 11446 3292
rect 11382 3232 11446 3236
rect 11462 3292 11526 3296
rect 11462 3236 11466 3292
rect 11466 3236 11522 3292
rect 11522 3236 11526 3292
rect 11462 3232 11526 3236
rect 11542 3292 11606 3296
rect 11542 3236 11546 3292
rect 11546 3236 11602 3292
rect 11602 3236 11606 3292
rect 11542 3232 11606 3236
rect 18202 3292 18266 3296
rect 18202 3236 18206 3292
rect 18206 3236 18262 3292
rect 18262 3236 18266 3292
rect 18202 3232 18266 3236
rect 18282 3292 18346 3296
rect 18282 3236 18286 3292
rect 18286 3236 18342 3292
rect 18342 3236 18346 3292
rect 18282 3232 18346 3236
rect 18362 3292 18426 3296
rect 18362 3236 18366 3292
rect 18366 3236 18422 3292
rect 18422 3236 18426 3292
rect 18362 3232 18426 3236
rect 18442 3292 18506 3296
rect 18442 3236 18446 3292
rect 18446 3236 18502 3292
rect 18502 3236 18506 3292
rect 18442 3232 18506 3236
rect 7852 2748 7916 2752
rect 7852 2692 7856 2748
rect 7856 2692 7912 2748
rect 7912 2692 7916 2748
rect 7852 2688 7916 2692
rect 7932 2748 7996 2752
rect 7932 2692 7936 2748
rect 7936 2692 7992 2748
rect 7992 2692 7996 2748
rect 7932 2688 7996 2692
rect 8012 2748 8076 2752
rect 8012 2692 8016 2748
rect 8016 2692 8072 2748
rect 8072 2692 8076 2748
rect 8012 2688 8076 2692
rect 8092 2748 8156 2752
rect 8092 2692 8096 2748
rect 8096 2692 8152 2748
rect 8152 2692 8156 2748
rect 8092 2688 8156 2692
rect 14752 2748 14816 2752
rect 14752 2692 14756 2748
rect 14756 2692 14812 2748
rect 14812 2692 14816 2748
rect 14752 2688 14816 2692
rect 14832 2748 14896 2752
rect 14832 2692 14836 2748
rect 14836 2692 14892 2748
rect 14892 2692 14896 2748
rect 14832 2688 14896 2692
rect 14912 2748 14976 2752
rect 14912 2692 14916 2748
rect 14916 2692 14972 2748
rect 14972 2692 14976 2748
rect 14912 2688 14976 2692
rect 14992 2748 15056 2752
rect 14992 2692 14996 2748
rect 14996 2692 15052 2748
rect 15052 2692 15056 2748
rect 14992 2688 15056 2692
rect 4402 2204 4466 2208
rect 4402 2148 4406 2204
rect 4406 2148 4462 2204
rect 4462 2148 4466 2204
rect 4402 2144 4466 2148
rect 4482 2204 4546 2208
rect 4482 2148 4486 2204
rect 4486 2148 4542 2204
rect 4542 2148 4546 2204
rect 4482 2144 4546 2148
rect 4562 2204 4626 2208
rect 4562 2148 4566 2204
rect 4566 2148 4622 2204
rect 4622 2148 4626 2204
rect 4562 2144 4626 2148
rect 4642 2204 4706 2208
rect 4642 2148 4646 2204
rect 4646 2148 4702 2204
rect 4702 2148 4706 2204
rect 4642 2144 4706 2148
rect 11302 2204 11366 2208
rect 11302 2148 11306 2204
rect 11306 2148 11362 2204
rect 11362 2148 11366 2204
rect 11302 2144 11366 2148
rect 11382 2204 11446 2208
rect 11382 2148 11386 2204
rect 11386 2148 11442 2204
rect 11442 2148 11446 2204
rect 11382 2144 11446 2148
rect 11462 2204 11526 2208
rect 11462 2148 11466 2204
rect 11466 2148 11522 2204
rect 11522 2148 11526 2204
rect 11462 2144 11526 2148
rect 11542 2204 11606 2208
rect 11542 2148 11546 2204
rect 11546 2148 11602 2204
rect 11602 2148 11606 2204
rect 11542 2144 11606 2148
rect 18202 2204 18266 2208
rect 18202 2148 18206 2204
rect 18206 2148 18262 2204
rect 18262 2148 18266 2204
rect 18202 2144 18266 2148
rect 18282 2204 18346 2208
rect 18282 2148 18286 2204
rect 18286 2148 18342 2204
rect 18342 2148 18346 2204
rect 18282 2144 18346 2148
rect 18362 2204 18426 2208
rect 18362 2148 18366 2204
rect 18366 2148 18422 2204
rect 18422 2148 18426 2204
rect 18362 2144 18426 2148
rect 18442 2204 18506 2208
rect 18442 2148 18446 2204
rect 18446 2148 18502 2204
rect 18502 2148 18506 2204
rect 18442 2144 18506 2148
<< metal4 >>
rect 4394 22880 4714 22896
rect 4394 22816 4402 22880
rect 4466 22816 4482 22880
rect 4546 22816 4562 22880
rect 4626 22816 4642 22880
rect 4706 22816 4714 22880
rect 4394 21792 4714 22816
rect 4394 21728 4402 21792
rect 4466 21728 4482 21792
rect 4546 21728 4562 21792
rect 4626 21728 4642 21792
rect 4706 21728 4714 21792
rect 4394 20704 4714 21728
rect 4394 20640 4402 20704
rect 4466 20640 4482 20704
rect 4546 20640 4562 20704
rect 4626 20640 4642 20704
rect 4706 20640 4714 20704
rect 4394 19616 4714 20640
rect 4394 19552 4402 19616
rect 4466 19552 4482 19616
rect 4546 19552 4562 19616
rect 4626 19552 4642 19616
rect 4706 19552 4714 19616
rect 4394 19472 4714 19552
rect 4394 19236 4436 19472
rect 4672 19236 4714 19472
rect 4394 18528 4714 19236
rect 4394 18464 4402 18528
rect 4466 18464 4482 18528
rect 4546 18464 4562 18528
rect 4626 18464 4642 18528
rect 4706 18464 4714 18528
rect 4394 17440 4714 18464
rect 4394 17376 4402 17440
rect 4466 17376 4482 17440
rect 4546 17376 4562 17440
rect 4626 17376 4642 17440
rect 4706 17376 4714 17440
rect 4394 16352 4714 17376
rect 4394 16288 4402 16352
rect 4466 16288 4482 16352
rect 4546 16288 4562 16352
rect 4626 16288 4642 16352
rect 4706 16288 4714 16352
rect 4394 15264 4714 16288
rect 4394 15200 4402 15264
rect 4466 15200 4482 15264
rect 4546 15200 4562 15264
rect 4626 15200 4642 15264
rect 4706 15200 4714 15264
rect 4394 14176 4714 15200
rect 4394 14112 4402 14176
rect 4466 14112 4482 14176
rect 4546 14112 4562 14176
rect 4626 14112 4642 14176
rect 4706 14112 4714 14176
rect 4394 13088 4714 14112
rect 4394 13024 4402 13088
rect 4466 13024 4482 13088
rect 4546 13024 4562 13088
rect 4626 13024 4642 13088
rect 4706 13024 4714 13088
rect 4394 12582 4714 13024
rect 4394 12346 4436 12582
rect 4672 12346 4714 12582
rect 4394 12000 4714 12346
rect 4394 11936 4402 12000
rect 4466 11936 4482 12000
rect 4546 11936 4562 12000
rect 4626 11936 4642 12000
rect 4706 11936 4714 12000
rect 4394 10912 4714 11936
rect 4394 10848 4402 10912
rect 4466 10848 4482 10912
rect 4546 10848 4562 10912
rect 4626 10848 4642 10912
rect 4706 10848 4714 10912
rect 4394 9824 4714 10848
rect 4394 9760 4402 9824
rect 4466 9760 4482 9824
rect 4546 9760 4562 9824
rect 4626 9760 4642 9824
rect 4706 9760 4714 9824
rect 4394 8736 4714 9760
rect 4394 8672 4402 8736
rect 4466 8672 4482 8736
rect 4546 8672 4562 8736
rect 4626 8672 4642 8736
rect 4706 8672 4714 8736
rect 4394 7648 4714 8672
rect 4394 7584 4402 7648
rect 4466 7584 4482 7648
rect 4546 7584 4562 7648
rect 4626 7584 4642 7648
rect 4706 7584 4714 7648
rect 4394 6560 4714 7584
rect 4394 6496 4402 6560
rect 4466 6496 4482 6560
rect 4546 6496 4562 6560
rect 4626 6496 4642 6560
rect 4706 6496 4714 6560
rect 4394 5691 4714 6496
rect 4394 5472 4436 5691
rect 4672 5472 4714 5691
rect 4394 5408 4402 5472
rect 4466 5408 4482 5455
rect 4546 5408 4562 5455
rect 4626 5408 4642 5455
rect 4706 5408 4714 5472
rect 4394 4384 4714 5408
rect 4394 4320 4402 4384
rect 4466 4320 4482 4384
rect 4546 4320 4562 4384
rect 4626 4320 4642 4384
rect 4706 4320 4714 4384
rect 4394 3296 4714 4320
rect 4394 3232 4402 3296
rect 4466 3232 4482 3296
rect 4546 3232 4562 3296
rect 4626 3232 4642 3296
rect 4706 3232 4714 3296
rect 4394 2208 4714 3232
rect 4394 2144 4402 2208
rect 4466 2144 4482 2208
rect 4546 2144 4562 2208
rect 4626 2144 4642 2208
rect 4706 2144 4714 2208
rect 4394 2128 4714 2144
rect 7844 22336 8164 22896
rect 7844 22272 7852 22336
rect 7916 22272 7932 22336
rect 7996 22272 8012 22336
rect 8076 22272 8092 22336
rect 8156 22272 8164 22336
rect 7844 21248 8164 22272
rect 7844 21184 7852 21248
rect 7916 21184 7932 21248
rect 7996 21184 8012 21248
rect 8076 21184 8092 21248
rect 8156 21184 8164 21248
rect 7844 20160 8164 21184
rect 7844 20096 7852 20160
rect 7916 20096 7932 20160
rect 7996 20096 8012 20160
rect 8076 20096 8092 20160
rect 8156 20096 8164 20160
rect 7844 19072 8164 20096
rect 7844 19008 7852 19072
rect 7916 19008 7932 19072
rect 7996 19008 8012 19072
rect 8076 19008 8092 19072
rect 8156 19008 8164 19072
rect 7844 17984 8164 19008
rect 7844 17920 7852 17984
rect 7916 17920 7932 17984
rect 7996 17920 8012 17984
rect 8076 17920 8092 17984
rect 8156 17920 8164 17984
rect 7844 16896 8164 17920
rect 7844 16832 7852 16896
rect 7916 16832 7932 16896
rect 7996 16832 8012 16896
rect 8076 16832 8092 16896
rect 8156 16832 8164 16896
rect 7844 16027 8164 16832
rect 7844 15808 7886 16027
rect 8122 15808 8164 16027
rect 7844 15744 7852 15808
rect 7916 15744 7932 15791
rect 7996 15744 8012 15791
rect 8076 15744 8092 15791
rect 8156 15744 8164 15808
rect 7844 14720 8164 15744
rect 7844 14656 7852 14720
rect 7916 14656 7932 14720
rect 7996 14656 8012 14720
rect 8076 14656 8092 14720
rect 8156 14656 8164 14720
rect 7844 13632 8164 14656
rect 7844 13568 7852 13632
rect 7916 13568 7932 13632
rect 7996 13568 8012 13632
rect 8076 13568 8092 13632
rect 8156 13568 8164 13632
rect 7844 12544 8164 13568
rect 7844 12480 7852 12544
rect 7916 12480 7932 12544
rect 7996 12480 8012 12544
rect 8076 12480 8092 12544
rect 8156 12480 8164 12544
rect 7844 11456 8164 12480
rect 7844 11392 7852 11456
rect 7916 11392 7932 11456
rect 7996 11392 8012 11456
rect 8076 11392 8092 11456
rect 8156 11392 8164 11456
rect 7844 10368 8164 11392
rect 7844 10304 7852 10368
rect 7916 10304 7932 10368
rect 7996 10304 8012 10368
rect 8076 10304 8092 10368
rect 8156 10304 8164 10368
rect 7844 9280 8164 10304
rect 7844 9216 7852 9280
rect 7916 9216 7932 9280
rect 7996 9216 8012 9280
rect 8076 9216 8092 9280
rect 8156 9216 8164 9280
rect 7844 9136 8164 9216
rect 7844 8900 7886 9136
rect 8122 8900 8164 9136
rect 7844 8192 8164 8900
rect 7844 8128 7852 8192
rect 7916 8128 7932 8192
rect 7996 8128 8012 8192
rect 8076 8128 8092 8192
rect 8156 8128 8164 8192
rect 7844 7104 8164 8128
rect 7844 7040 7852 7104
rect 7916 7040 7932 7104
rect 7996 7040 8012 7104
rect 8076 7040 8092 7104
rect 8156 7040 8164 7104
rect 7844 6016 8164 7040
rect 7844 5952 7852 6016
rect 7916 5952 7932 6016
rect 7996 5952 8012 6016
rect 8076 5952 8092 6016
rect 8156 5952 8164 6016
rect 7844 4928 8164 5952
rect 7844 4864 7852 4928
rect 7916 4864 7932 4928
rect 7996 4864 8012 4928
rect 8076 4864 8092 4928
rect 8156 4864 8164 4928
rect 7844 3840 8164 4864
rect 7844 3776 7852 3840
rect 7916 3776 7932 3840
rect 7996 3776 8012 3840
rect 8076 3776 8092 3840
rect 8156 3776 8164 3840
rect 7844 2752 8164 3776
rect 7844 2688 7852 2752
rect 7916 2688 7932 2752
rect 7996 2688 8012 2752
rect 8076 2688 8092 2752
rect 8156 2688 8164 2752
rect 7844 2128 8164 2688
rect 11294 22880 11614 22896
rect 11294 22816 11302 22880
rect 11366 22816 11382 22880
rect 11446 22816 11462 22880
rect 11526 22816 11542 22880
rect 11606 22816 11614 22880
rect 11294 21792 11614 22816
rect 11294 21728 11302 21792
rect 11366 21728 11382 21792
rect 11446 21728 11462 21792
rect 11526 21728 11542 21792
rect 11606 21728 11614 21792
rect 11294 20704 11614 21728
rect 11294 20640 11302 20704
rect 11366 20640 11382 20704
rect 11446 20640 11462 20704
rect 11526 20640 11542 20704
rect 11606 20640 11614 20704
rect 11294 19616 11614 20640
rect 11294 19552 11302 19616
rect 11366 19552 11382 19616
rect 11446 19552 11462 19616
rect 11526 19552 11542 19616
rect 11606 19552 11614 19616
rect 11294 19472 11614 19552
rect 11294 19236 11336 19472
rect 11572 19236 11614 19472
rect 11294 18528 11614 19236
rect 11294 18464 11302 18528
rect 11366 18464 11382 18528
rect 11446 18464 11462 18528
rect 11526 18464 11542 18528
rect 11606 18464 11614 18528
rect 11294 17440 11614 18464
rect 11294 17376 11302 17440
rect 11366 17376 11382 17440
rect 11446 17376 11462 17440
rect 11526 17376 11542 17440
rect 11606 17376 11614 17440
rect 11294 16352 11614 17376
rect 11294 16288 11302 16352
rect 11366 16288 11382 16352
rect 11446 16288 11462 16352
rect 11526 16288 11542 16352
rect 11606 16288 11614 16352
rect 11294 15264 11614 16288
rect 11294 15200 11302 15264
rect 11366 15200 11382 15264
rect 11446 15200 11462 15264
rect 11526 15200 11542 15264
rect 11606 15200 11614 15264
rect 11294 14176 11614 15200
rect 11294 14112 11302 14176
rect 11366 14112 11382 14176
rect 11446 14112 11462 14176
rect 11526 14112 11542 14176
rect 11606 14112 11614 14176
rect 11294 13088 11614 14112
rect 11294 13024 11302 13088
rect 11366 13024 11382 13088
rect 11446 13024 11462 13088
rect 11526 13024 11542 13088
rect 11606 13024 11614 13088
rect 11294 12582 11614 13024
rect 11294 12346 11336 12582
rect 11572 12346 11614 12582
rect 11294 12000 11614 12346
rect 11294 11936 11302 12000
rect 11366 11936 11382 12000
rect 11446 11936 11462 12000
rect 11526 11936 11542 12000
rect 11606 11936 11614 12000
rect 11294 10912 11614 11936
rect 11294 10848 11302 10912
rect 11366 10848 11382 10912
rect 11446 10848 11462 10912
rect 11526 10848 11542 10912
rect 11606 10848 11614 10912
rect 11294 9824 11614 10848
rect 11294 9760 11302 9824
rect 11366 9760 11382 9824
rect 11446 9760 11462 9824
rect 11526 9760 11542 9824
rect 11606 9760 11614 9824
rect 11294 8736 11614 9760
rect 11294 8672 11302 8736
rect 11366 8672 11382 8736
rect 11446 8672 11462 8736
rect 11526 8672 11542 8736
rect 11606 8672 11614 8736
rect 11294 7648 11614 8672
rect 11294 7584 11302 7648
rect 11366 7584 11382 7648
rect 11446 7584 11462 7648
rect 11526 7584 11542 7648
rect 11606 7584 11614 7648
rect 11294 6560 11614 7584
rect 11294 6496 11302 6560
rect 11366 6496 11382 6560
rect 11446 6496 11462 6560
rect 11526 6496 11542 6560
rect 11606 6496 11614 6560
rect 11294 5691 11614 6496
rect 11294 5472 11336 5691
rect 11572 5472 11614 5691
rect 11294 5408 11302 5472
rect 11366 5408 11382 5455
rect 11446 5408 11462 5455
rect 11526 5408 11542 5455
rect 11606 5408 11614 5472
rect 11294 4384 11614 5408
rect 11294 4320 11302 4384
rect 11366 4320 11382 4384
rect 11446 4320 11462 4384
rect 11526 4320 11542 4384
rect 11606 4320 11614 4384
rect 11294 3296 11614 4320
rect 11294 3232 11302 3296
rect 11366 3232 11382 3296
rect 11446 3232 11462 3296
rect 11526 3232 11542 3296
rect 11606 3232 11614 3296
rect 11294 2208 11614 3232
rect 11294 2144 11302 2208
rect 11366 2144 11382 2208
rect 11446 2144 11462 2208
rect 11526 2144 11542 2208
rect 11606 2144 11614 2208
rect 11294 2128 11614 2144
rect 14744 22336 15064 22896
rect 14744 22272 14752 22336
rect 14816 22272 14832 22336
rect 14896 22272 14912 22336
rect 14976 22272 14992 22336
rect 15056 22272 15064 22336
rect 14744 21248 15064 22272
rect 14744 21184 14752 21248
rect 14816 21184 14832 21248
rect 14896 21184 14912 21248
rect 14976 21184 14992 21248
rect 15056 21184 15064 21248
rect 14744 20160 15064 21184
rect 14744 20096 14752 20160
rect 14816 20096 14832 20160
rect 14896 20096 14912 20160
rect 14976 20096 14992 20160
rect 15056 20096 15064 20160
rect 14744 19072 15064 20096
rect 14744 19008 14752 19072
rect 14816 19008 14832 19072
rect 14896 19008 14912 19072
rect 14976 19008 14992 19072
rect 15056 19008 15064 19072
rect 14744 17984 15064 19008
rect 14744 17920 14752 17984
rect 14816 17920 14832 17984
rect 14896 17920 14912 17984
rect 14976 17920 14992 17984
rect 15056 17920 15064 17984
rect 14744 16896 15064 17920
rect 14744 16832 14752 16896
rect 14816 16832 14832 16896
rect 14896 16832 14912 16896
rect 14976 16832 14992 16896
rect 15056 16832 15064 16896
rect 14744 16027 15064 16832
rect 14744 15808 14786 16027
rect 15022 15808 15064 16027
rect 14744 15744 14752 15808
rect 14816 15744 14832 15791
rect 14896 15744 14912 15791
rect 14976 15744 14992 15791
rect 15056 15744 15064 15808
rect 14744 14720 15064 15744
rect 14744 14656 14752 14720
rect 14816 14656 14832 14720
rect 14896 14656 14912 14720
rect 14976 14656 14992 14720
rect 15056 14656 15064 14720
rect 14744 13632 15064 14656
rect 14744 13568 14752 13632
rect 14816 13568 14832 13632
rect 14896 13568 14912 13632
rect 14976 13568 14992 13632
rect 15056 13568 15064 13632
rect 14744 12544 15064 13568
rect 14744 12480 14752 12544
rect 14816 12480 14832 12544
rect 14896 12480 14912 12544
rect 14976 12480 14992 12544
rect 15056 12480 15064 12544
rect 14744 11456 15064 12480
rect 14744 11392 14752 11456
rect 14816 11392 14832 11456
rect 14896 11392 14912 11456
rect 14976 11392 14992 11456
rect 15056 11392 15064 11456
rect 14744 10368 15064 11392
rect 14744 10304 14752 10368
rect 14816 10304 14832 10368
rect 14896 10304 14912 10368
rect 14976 10304 14992 10368
rect 15056 10304 15064 10368
rect 14744 9280 15064 10304
rect 14744 9216 14752 9280
rect 14816 9216 14832 9280
rect 14896 9216 14912 9280
rect 14976 9216 14992 9280
rect 15056 9216 15064 9280
rect 14744 9136 15064 9216
rect 14744 8900 14786 9136
rect 15022 8900 15064 9136
rect 14744 8192 15064 8900
rect 14744 8128 14752 8192
rect 14816 8128 14832 8192
rect 14896 8128 14912 8192
rect 14976 8128 14992 8192
rect 15056 8128 15064 8192
rect 14744 7104 15064 8128
rect 14744 7040 14752 7104
rect 14816 7040 14832 7104
rect 14896 7040 14912 7104
rect 14976 7040 14992 7104
rect 15056 7040 15064 7104
rect 14744 6016 15064 7040
rect 14744 5952 14752 6016
rect 14816 5952 14832 6016
rect 14896 5952 14912 6016
rect 14976 5952 14992 6016
rect 15056 5952 15064 6016
rect 14744 4928 15064 5952
rect 14744 4864 14752 4928
rect 14816 4864 14832 4928
rect 14896 4864 14912 4928
rect 14976 4864 14992 4928
rect 15056 4864 15064 4928
rect 14744 3840 15064 4864
rect 14744 3776 14752 3840
rect 14816 3776 14832 3840
rect 14896 3776 14912 3840
rect 14976 3776 14992 3840
rect 15056 3776 15064 3840
rect 14744 2752 15064 3776
rect 14744 2688 14752 2752
rect 14816 2688 14832 2752
rect 14896 2688 14912 2752
rect 14976 2688 14992 2752
rect 15056 2688 15064 2752
rect 14744 2128 15064 2688
rect 18194 22880 18514 22896
rect 18194 22816 18202 22880
rect 18266 22816 18282 22880
rect 18346 22816 18362 22880
rect 18426 22816 18442 22880
rect 18506 22816 18514 22880
rect 18194 21792 18514 22816
rect 18194 21728 18202 21792
rect 18266 21728 18282 21792
rect 18346 21728 18362 21792
rect 18426 21728 18442 21792
rect 18506 21728 18514 21792
rect 18194 20704 18514 21728
rect 18194 20640 18202 20704
rect 18266 20640 18282 20704
rect 18346 20640 18362 20704
rect 18426 20640 18442 20704
rect 18506 20640 18514 20704
rect 18194 19616 18514 20640
rect 18194 19552 18202 19616
rect 18266 19552 18282 19616
rect 18346 19552 18362 19616
rect 18426 19552 18442 19616
rect 18506 19552 18514 19616
rect 18194 19472 18514 19552
rect 18194 19236 18236 19472
rect 18472 19236 18514 19472
rect 18194 18528 18514 19236
rect 18194 18464 18202 18528
rect 18266 18464 18282 18528
rect 18346 18464 18362 18528
rect 18426 18464 18442 18528
rect 18506 18464 18514 18528
rect 18194 17440 18514 18464
rect 18194 17376 18202 17440
rect 18266 17376 18282 17440
rect 18346 17376 18362 17440
rect 18426 17376 18442 17440
rect 18506 17376 18514 17440
rect 18194 16352 18514 17376
rect 18194 16288 18202 16352
rect 18266 16288 18282 16352
rect 18346 16288 18362 16352
rect 18426 16288 18442 16352
rect 18506 16288 18514 16352
rect 18194 15264 18514 16288
rect 18194 15200 18202 15264
rect 18266 15200 18282 15264
rect 18346 15200 18362 15264
rect 18426 15200 18442 15264
rect 18506 15200 18514 15264
rect 18194 14176 18514 15200
rect 18194 14112 18202 14176
rect 18266 14112 18282 14176
rect 18346 14112 18362 14176
rect 18426 14112 18442 14176
rect 18506 14112 18514 14176
rect 18194 13088 18514 14112
rect 18194 13024 18202 13088
rect 18266 13024 18282 13088
rect 18346 13024 18362 13088
rect 18426 13024 18442 13088
rect 18506 13024 18514 13088
rect 18194 12582 18514 13024
rect 18194 12346 18236 12582
rect 18472 12346 18514 12582
rect 18194 12000 18514 12346
rect 18194 11936 18202 12000
rect 18266 11936 18282 12000
rect 18346 11936 18362 12000
rect 18426 11936 18442 12000
rect 18506 11936 18514 12000
rect 18194 10912 18514 11936
rect 18194 10848 18202 10912
rect 18266 10848 18282 10912
rect 18346 10848 18362 10912
rect 18426 10848 18442 10912
rect 18506 10848 18514 10912
rect 18194 9824 18514 10848
rect 18194 9760 18202 9824
rect 18266 9760 18282 9824
rect 18346 9760 18362 9824
rect 18426 9760 18442 9824
rect 18506 9760 18514 9824
rect 18194 8736 18514 9760
rect 18194 8672 18202 8736
rect 18266 8672 18282 8736
rect 18346 8672 18362 8736
rect 18426 8672 18442 8736
rect 18506 8672 18514 8736
rect 18194 7648 18514 8672
rect 18194 7584 18202 7648
rect 18266 7584 18282 7648
rect 18346 7584 18362 7648
rect 18426 7584 18442 7648
rect 18506 7584 18514 7648
rect 18194 6560 18514 7584
rect 18194 6496 18202 6560
rect 18266 6496 18282 6560
rect 18346 6496 18362 6560
rect 18426 6496 18442 6560
rect 18506 6496 18514 6560
rect 18194 5691 18514 6496
rect 18194 5472 18236 5691
rect 18472 5472 18514 5691
rect 18194 5408 18202 5472
rect 18266 5408 18282 5455
rect 18346 5408 18362 5455
rect 18426 5408 18442 5455
rect 18506 5408 18514 5472
rect 18194 4384 18514 5408
rect 18194 4320 18202 4384
rect 18266 4320 18282 4384
rect 18346 4320 18362 4384
rect 18426 4320 18442 4384
rect 18506 4320 18514 4384
rect 18194 3296 18514 4320
rect 18194 3232 18202 3296
rect 18266 3232 18282 3296
rect 18346 3232 18362 3296
rect 18426 3232 18442 3296
rect 18506 3232 18514 3296
rect 18194 2208 18514 3232
rect 18194 2144 18202 2208
rect 18266 2144 18282 2208
rect 18346 2144 18362 2208
rect 18426 2144 18442 2208
rect 18506 2144 18514 2208
rect 18194 2128 18514 2144
<< via4 >>
rect 4436 19236 4672 19472
rect 4436 12346 4672 12582
rect 4436 5472 4672 5691
rect 4436 5455 4466 5472
rect 4466 5455 4482 5472
rect 4482 5455 4546 5472
rect 4546 5455 4562 5472
rect 4562 5455 4626 5472
rect 4626 5455 4642 5472
rect 4642 5455 4672 5472
rect 7886 15808 8122 16027
rect 7886 15791 7916 15808
rect 7916 15791 7932 15808
rect 7932 15791 7996 15808
rect 7996 15791 8012 15808
rect 8012 15791 8076 15808
rect 8076 15791 8092 15808
rect 8092 15791 8122 15808
rect 7886 8900 8122 9136
rect 11336 19236 11572 19472
rect 11336 12346 11572 12582
rect 11336 5472 11572 5691
rect 11336 5455 11366 5472
rect 11366 5455 11382 5472
rect 11382 5455 11446 5472
rect 11446 5455 11462 5472
rect 11462 5455 11526 5472
rect 11526 5455 11542 5472
rect 11542 5455 11572 5472
rect 14786 15808 15022 16027
rect 14786 15791 14816 15808
rect 14816 15791 14832 15808
rect 14832 15791 14896 15808
rect 14896 15791 14912 15808
rect 14912 15791 14976 15808
rect 14976 15791 14992 15808
rect 14992 15791 15022 15808
rect 14786 8900 15022 9136
rect 18236 19236 18472 19472
rect 18236 12346 18472 12582
rect 18236 5472 18472 5691
rect 18236 5455 18266 5472
rect 18266 5455 18282 5472
rect 18282 5455 18346 5472
rect 18346 5455 18362 5472
rect 18362 5455 18426 5472
rect 18426 5455 18442 5472
rect 18442 5455 18472 5472
<< metal5 >>
rect 1104 19472 21804 19515
rect 1104 19236 4436 19472
rect 4672 19236 11336 19472
rect 11572 19236 18236 19472
rect 18472 19236 21804 19472
rect 1104 19194 21804 19236
rect 1104 16027 21804 16069
rect 1104 15791 7886 16027
rect 8122 15791 14786 16027
rect 15022 15791 21804 16027
rect 1104 15749 21804 15791
rect 1104 12582 21804 12624
rect 1104 12346 4436 12582
rect 4672 12346 11336 12582
rect 11572 12346 18236 12582
rect 18472 12346 21804 12582
rect 1104 12304 21804 12346
rect 1104 9136 21804 9179
rect 1104 8900 7886 9136
rect 8122 8900 14786 9136
rect 15022 8900 21804 9136
rect 1104 8858 21804 8900
rect 1104 5691 21804 5733
rect 1104 5455 4436 5691
rect 4672 5455 11336 5691
rect 11572 5455 18236 5691
rect 18472 5455 21804 5691
rect 1104 5413 21804 5455
use sky130_fd_sc_hd__fill_1  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 2208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1619507013
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1618419204
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1618419204
transform 1 0 3312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 2760 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_6
timestamp 1618419204
transform 1 0 1656 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_12
timestamp 1618419204
transform 1 0 2208 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 4508 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1618419204
transform -1 0 5796 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28
timestamp 1618419204
transform 1 0 3680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30
timestamp 1618419204
transform 1 0 3864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 4508 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45
timestamp 1618419204
transform 1 0 5244 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_30
timestamp 1618419204
transform 1 0 3864 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_42
timestamp 1618419204
transform 1 0 4968 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_54
timestamp 1618419204
transform 1 0 6072 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1618419204
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1618419204
transform 1 0 6348 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 5796 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1618419204
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1618419204
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_70
timestamp 1618419204
transform 1 0 7544 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1618419204
transform -1 0 7268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_58
timestamp 1618419204
transform 1 0 6440 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_67
timestamp 1618419204
transform 1 0 7268 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79
timestamp 1618419204
transform 1 0 8372 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _369_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 9108 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_87
timestamp 1618419204
transform 1 0 9108 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1618419204
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1618419204
transform -1 0 9844 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1618419204
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb1
timestamp 1619507013
transform 1 0 9476 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_1_98
timestamp 1618419204
transform 1 0 10120 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95
timestamp 1618419204
transform 1 0 9844 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1618419204
transform 1 0 10212 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_102
timestamp 1618419204
transform 1 0 10488 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1618419204
transform 1 0 10580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[11\].id.delayenb1
timestamp 1619507013
transform 1 0 10580 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[11\].id.delayen1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 10948 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_1_115
timestamp 1618419204
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1618419204
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117
timestamp 1618419204
transform 1 0 11868 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1618419204
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1618419204
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1618419204
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_122
timestamp 1618419204
transform 1 0 12328 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1619507013
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129
timestamp 1618419204
transform 1 0 12972 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125
timestamp 1618419204
transform 1 0 12604 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1618419204
transform -1 0 12972 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb1
timestamp 1619507013
transform 1 0 13340 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp 1618419204
transform -1 0 13892 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1618419204
transform 1 0 13892 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_140
timestamp 1618419204
transform 1 0 13984 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen1
timestamp 1618419204
transform 1 0 14260 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_1_148
timestamp 1618419204
transform 1 0 14720 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1618419204
transform 1 0 14536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144
timestamp 1618419204
transform 1 0 14352 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1618419204
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_156
timestamp 1618419204
transform 1 0 15456 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_157
timestamp 1618419204
transform 1 0 15548 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1618419204
transform 1 0 15180 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1618419204
transform 1 0 14904 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1618419204
transform 1 0 15548 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1618419204
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_170
timestamp 1618419204
transform 1 0 16744 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_166
timestamp 1618419204
transform 1 0 16376 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_170
timestamp 1618419204
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1618419204
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 15640 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrbp_2  idiv8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 17296 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1618419204
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1618419204
transform 1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1618419204
transform 1 0 17572 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1618419204
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_183
timestamp 1618419204
transform 1 0 17940 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_191 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_196
timestamp 1618419204
transform 1 0 19136 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_204
timestamp 1618419204
transform 1 0 19872 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_202
timestamp 1618419204
transform 1 0 19688 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1618419204
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_218
timestamp 1618419204
transform 1 0 21160 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_212
timestamp 1618419204
transform 1 0 20608 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_221
timestamp 1618419204
transform 1 0 21436 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_217
timestamp 1618419204
transform 1 0 21068 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_212
timestamp 1618419204
transform 1 0 20608 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output43
timestamp 1618419204
transform -1 0 21068 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1619507013
transform -1 0 21160 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1618419204
transform -1 0 21804 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1618419204
transform -1 0 21804 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_200
timestamp 1618419204
transform 1 0 19504 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1618419204
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1618419204
transform -1 0 1656 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_6
timestamp 1618419204
transform 1 0 1656 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1618419204
transform 1 0 2760 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1618419204
transform 1 0 4232 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1618419204
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_26
timestamp 1618419204
transform 1 0 3496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_30
timestamp 1618419204
transform 1 0 3864 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_38
timestamp 1618419204
transform 1 0 4600 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_4  irb
timestamp 1619507013
transform -1 0 7084 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_2_50
timestamp 1618419204
transform 1 0 5704 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_58
timestamp 1618419204
transform 1 0 6440 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1618419204
transform 1 0 7084 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1618419204
transform 1 0 9476 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen1
timestamp 1618419204
transform 1 0 8188 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1618419204
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_82
timestamp 1618419204
transform 1 0 8648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1618419204
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_94
timestamp 1618419204
transform 1 0 9752 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1618419204
transform 1 0 10856 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1618419204
transform 1 0 12052 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_115
timestamp 1618419204
transform 1 0 11684 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_122
timestamp 1618419204
transform 1 0 12328 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1618419204
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1618419204
transform 1 0 12696 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1618419204
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1618419204
transform 1 0 14076 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_144
timestamp 1618419204
transform 1 0 14352 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen0
timestamp 1618419204
transform -1 0 16376 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb0
timestamp 1619507013
transform -1 0 15548 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_157
timestamp 1618419204
transform 1 0 15548 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1618419204
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1618419204
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_190
timestamp 1618419204
transform 1 0 18584 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_198
timestamp 1618419204
transform 1 0 19320 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1618419204
transform -1 0 21804 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1618419204
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1618419204
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_201
timestamp 1618419204
transform 1 0 19596 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_213
timestamp 1618419204
transform 1 0 20700 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_218
timestamp 1618419204
transform 1 0 21160 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1618419204
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1618419204
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1618419204
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1618419204
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1618419204
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen0
timestamp 1618419204
transform 1 0 7912 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1618419204
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1618419204
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1618419204
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_70
timestamp 1618419204
transform 1 0 7544 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _356_
timestamp 1618419204
transform -1 0 10304 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 9016 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_79
timestamp 1618419204
transform 1 0 8372 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_86
timestamp 1618419204
transform 1 0 9016 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_90
timestamp 1618419204
transform 1 0 9384 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1618419204
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1618419204
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_100
timestamp 1618419204
transform 1 0 10304 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_112
timestamp 1618419204
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1618419204
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_122
timestamp 1618419204
transform 1 0 12328 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1618419204
transform 1 0 14720 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_134
timestamp 1618419204
transform 1 0 13432 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_146
timestamp 1618419204
transform 1 0 14536 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1618419204
transform -1 0 15732 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1618419204
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_151
timestamp 1618419204
transform 1 0 14996 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1618419204
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_172
timestamp 1618419204
transform 1 0 16928 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrbp_1  idiv16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 18124 0 1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_3_184
timestamp 1618419204
transform 1 0 18032 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1618419204
transform -1 0 21804 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1618419204
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_220
timestamp 1618419204
transform 1 0 21344 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1618419204
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1618419204
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1618419204
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrbp_2  idiv4
timestamp 1618419204
transform -1 0 7084 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1618419204
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1618419204
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_30
timestamp 1618419204
transform 1 0 3864 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_38
timestamp 1618419204
transform 1 0 4600 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _368_
timestamp 1618419204
transform 1 0 7820 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_65
timestamp 1618419204
transform 1 0 7084 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1618419204
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_82
timestamp 1618419204
transform 1 0 8648 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_87
timestamp 1618419204
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_99
timestamp 1618419204
transform 1 0 10212 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_4  ringosc.dstage\[11\].id.delayen0
timestamp 1619507013
transform 1 0 10488 0 -1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_12  FILLER_4_113
timestamp 1618419204
transform 1 0 11500 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1618419204
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_125
timestamp 1618419204
transform 1 0 12604 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_137
timestamp 1618419204
transform 1 0 13708 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144
timestamp 1618419204
transform 1 0 14352 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_156
timestamp 1618419204
transform 1 0 15456 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_168
timestamp 1618419204
transform 1 0 16560 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1618419204
transform 1 0 17940 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_180
timestamp 1618419204
transform 1 0 17664 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_192
timestamp 1618419204
transform 1 0 18768 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1618419204
transform -1 0 21804 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1618419204
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_201
timestamp 1618419204
transform 1 0 19596 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_213
timestamp 1618419204
transform 1 0 20700 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_221
timestamp 1618419204
transform 1 0 21436 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfrbp_2  idiv2
timestamp 1618419204
transform 1 0 2944 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1618419204
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1618419204
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1618419204
transform 1 0 2484 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_19
timestamp 1618419204
transform 1 0 2852 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1618419204
transform 1 0 5152 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb0
timestamp 1619507013
transform 1 0 7544 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1618419204
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_56
timestamp 1618419204
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1618419204
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb0
timestamp 1619507013
transform 1 0 10212 0 1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_12  FILLER_5_77
timestamp 1618419204
transform 1 0 8188 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_89
timestamp 1618419204
transform 1 0 9292 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_97
timestamp 1618419204
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb0
timestamp 1619507013
transform 1 0 12420 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1618419204
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_110
timestamp 1618419204
transform 1 0 11224 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_115
timestamp 1618419204
transform 1 0 11684 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen0
timestamp 1618419204
transform 1 0 13432 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1618419204
transform -1 0 14720 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_130
timestamp 1618419204
transform 1 0 13064 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_139
timestamp 1618419204
transform 1 0 13892 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_148
timestamp 1618419204
transform 1 0 14720 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1618419204
transform 1 0 15088 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1618419204
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_155
timestamp 1618419204
transform 1 0 15364 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_167
timestamp 1618419204
transform 1 0 16468 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_172
timestamp 1618419204
transform 1 0 16928 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1619507013
transform 1 0 18492 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1618419204
transform 1 0 17296 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_185
timestamp 1618419204
transform 1 0 18124 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_192
timestamp 1618419204
transform 1 0 18768 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1618419204
transform -1 0 21804 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_204
timestamp 1618419204
transform 1 0 19872 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_216
timestamp 1618419204
transform 1 0 20976 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_7
timestamp 1618419204
transform 1 0 1748 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output41
timestamp 1618419204
transform -1 0 1748 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1618419204
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1618419204
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_23
timestamp 1618419204
transform 1 0 3220 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_15
timestamp 1618419204
transform 1 0 2484 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_19
timestamp 1618419204
transform 1 0 2852 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_15
timestamp 1618419204
transform 1 0 2484 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  ringosc.ibufp11
timestamp 1619507013
transform -1 0 2852 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  ringosc.ibufp10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 3588 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1618419204
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[5\].id.delayen1
timestamp 1618419204
transform 1 0 5520 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1618419204
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1618419204
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1618419204
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1618419204
transform 1 0 4968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1618419204
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_39
timestamp 1618419204
transform 1 0 4692 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_47
timestamp 1618419204
transform 1 0 5428 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1618419204
transform -1 0 7176 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1618419204
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1618419204
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_54
timestamp 1618419204
transform 1 0 6072 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_66
timestamp 1618419204
transform 1 0 7176 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_53
timestamp 1618419204
transform 1 0 5980 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_58
timestamp 1618419204
transform 1 0 6440 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_65
timestamp 1618419204
transform 1 0 7084 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.delayen1
timestamp 1618419204
transform 1 0 9844 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1618419204
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_78
timestamp 1618419204
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_87
timestamp 1618419204
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_99
timestamp 1618419204
transform 1 0 10212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_77
timestamp 1618419204
transform 1 0 8188 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_89
timestamp 1618419204
transform 1 0 9292 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1618419204
transform -1 0 12880 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1618419204
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_111
timestamp 1618419204
transform 1 0 11316 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_123
timestamp 1618419204
transform 1 0 12420 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_100
timestamp 1618419204
transform 1 0 10304 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_112
timestamp 1618419204
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_115
timestamp 1618419204
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_136
timestamp 1618419204
transform 1 0 13616 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_128
timestamp 1618419204
transform 1 0 12880 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1618419204
transform -1 0 13616 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_139
timestamp 1618419204
transform 1 0 13892 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_144
timestamp 1618419204
transform 1 0 14352 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_142
timestamp 1618419204
transform 1 0 14168 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1618419204
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb1
timestamp 1619507013
transform 1 0 14720 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen1
timestamp 1618419204
transform 1 0 14628 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1618419204
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1618419204
transform 1 0 16100 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1618419204
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_155
timestamp 1618419204
transform 1 0 15364 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_172
timestamp 1618419204
transform 1 0 16928 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_152
timestamp 1618419204
transform 1 0 15088 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_164
timestamp 1618419204
transform 1 0 16192 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_170
timestamp 1618419204
transform 1 0 16744 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_172
timestamp 1618419204
transform 1 0 16928 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1619507013
transform -1 0 18768 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _322_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 18032 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _323_
timestamp 1618419204
transform -1 0 18124 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _325_
timestamp 1618419204
transform 1 0 18400 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_176
timestamp 1618419204
transform 1 0 17296 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_185
timestamp 1618419204
transform 1 0 18124 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_192
timestamp 1618419204
transform 1 0 18768 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_184
timestamp 1618419204
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1618419204
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1618419204
transform -1 0 21804 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1618419204
transform -1 0 21804 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1618419204
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1619507013
transform -1 0 21160 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_201
timestamp 1618419204
transform 1 0 19596 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_213
timestamp 1618419204
transform 1 0 20700 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_218
timestamp 1618419204
transform 1 0 21160 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1618419204
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_220
timestamp 1618419204
transform 1 0 21344 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1618419204
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1618419204
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1618419204
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb0
timestamp 1619507013
transform 1 0 4232 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[5\].id.delayenb1
timestamp 1619507013
transform -1 0 6256 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1618419204
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1618419204
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_30
timestamp 1618419204
transform 1 0 3864 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_45
timestamp 1618419204
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1618419204
transform 1 0 7820 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1618419204
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_68
timestamp 1618419204
transform 1 0 7360 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_72
timestamp 1618419204
transform 1 0 7728 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.iss.delayenb1
timestamp 1619507013
transform 1 0 9844 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1618419204
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_82
timestamp 1618419204
transform 1 0 8648 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_87
timestamp 1618419204
transform 1 0 9108 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1618419204
transform 1 0 10856 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_102
timestamp 1618419204
transform 1 0 10488 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1618419204
transform 1 0 11132 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1618419204
transform 1 0 12236 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1618419204
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_133
timestamp 1618419204
transform 1 0 13340 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1618419204
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1618419204
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1618419204
transform 1 0 15548 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_156
timestamp 1618419204
transform 1 0 15456 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_166
timestamp 1618419204
transform 1 0 16376 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _324_
timestamp 1618419204
transform -1 0 18124 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_174
timestamp 1618419204
transform 1 0 17112 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_185
timestamp 1618419204
transform 1 0 18124 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp 1618419204
transform 1 0 19228 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1618419204
transform -1 0 21804 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1618419204
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_201
timestamp 1618419204
transform 1 0 19596 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_213
timestamp 1618419204
transform 1 0 20700 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_221
timestamp 1618419204
transform 1 0 21436 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1618419204
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1618419204
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1618419204
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1619507013
transform 1 0 4692 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1618419204
transform -1 0 4048 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1618419204
transform 1 0 3588 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_32
timestamp 1618419204
transform 1 0 4048 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_38
timestamp 1618419204
transform 1 0 4600 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_46
timestamp 1618419204
transform 1 0 5336 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1618419204
transform -1 0 5980 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 7728 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1618419204
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_53
timestamp 1618419204
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1618419204
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_70
timestamp 1618419204
transform 1 0 7544 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.delayen0
timestamp 1619507013
transform 1 0 8556 0 1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb0
timestamp 1619507013
transform 1 0 9936 0 1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_9_77
timestamp 1618419204
transform 1 0 8188 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_92
timestamp 1618419204
transform 1 0 9568 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb0
timestamp 1619507013
transform 1 0 12236 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1618419204
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_107
timestamp 1618419204
transform 1 0 10948 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1618419204
transform 1 0 11500 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_115
timestamp 1618419204
transform 1 0 11684 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen0
timestamp 1618419204
transform 1 0 13248 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1618419204
transform -1 0 14352 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_128
timestamp 1618419204
transform 1 0 12880 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_137
timestamp 1618419204
transform 1 0 13708 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_144
timestamp 1618419204
transform 1 0 14352 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1618419204
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_156
timestamp 1618419204
transform 1 0 15456 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_168
timestamp 1618419204
transform 1 0 16560 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_172
timestamp 1618419204
transform 1 0 16928 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1618419204
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1618419204
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1618419204
transform -1 0 21804 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1618419204
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_220
timestamp 1618419204
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb0
timestamp 1619507013
transform 1 0 2116 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1618419204
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1618419204
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_18
timestamp 1618419204
transform 1 0 2760 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1618419204
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_26
timestamp 1618419204
transform 1 0 3496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1618419204
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1618419204
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 8096 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_10_54
timestamp 1618419204
transform 1 0 6072 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_62
timestamp 1618419204
transform 1 0 6808 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1618419204
transform -1 0 9936 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1618419204
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1618419204
transform 1 0 8096 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1618419204
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_87
timestamp 1618419204
transform 1 0 9108 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_96
timestamp 1618419204
transform 1 0 9936 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1618419204
transform -1 0 13248 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_108
timestamp 1618419204
transform 1 0 11040 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_120
timestamp 1618419204
transform 1 0 12144 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb1
timestamp 1619507013
transform 1 0 14720 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1618419204
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_132
timestamp 1618419204
transform 1 0 13248 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_140
timestamp 1618419204
transform 1 0 13984 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_144
timestamp 1618419204
transform 1 0 14352 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1618419204
transform -1 0 16560 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_155
timestamp 1618419204
transform 1 0 15364 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_163
timestamp 1618419204
transform 1 0 16100 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_168
timestamp 1618419204
transform 1 0 16560 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1618419204
transform -1 0 18492 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_180
timestamp 1618419204
transform 1 0 17664 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_189
timestamp 1618419204
transform 1 0 18492 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp 1618419204
transform 1 0 19228 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1618419204
transform -1 0 21804 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1618419204
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1618419204
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_213
timestamp 1618419204
transform 1 0 20700 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_221
timestamp 1618419204
transform 1 0 21436 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _360_
timestamp 1618419204
transform 1 0 2116 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1619507013
transform 1 0 3312 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1618419204
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1618419204
transform -1 0 1656 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_6
timestamp 1618419204
transform 1 0 1656 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_10
timestamp 1618419204
transform 1 0 2024 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_20
timestamp 1618419204
transform 1 0 2944 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_31
timestamp 1618419204
transform 1 0 3956 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_43
timestamp 1618419204
transform 1 0 5060 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1
timestamp 1619507013
transform -1 0 7176 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.reseten0
timestamp 1619507013
transform 1 0 7544 0 1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1618419204
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_55
timestamp 1618419204
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_58
timestamp 1618419204
transform 1 0 6440 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_62
timestamp 1618419204
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_66
timestamp 1618419204
transform 1 0 7176 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _306_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 9476 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_11_81
timestamp 1618419204
transform 1 0 8556 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_89
timestamp 1618419204
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_96
timestamp 1618419204
transform 1 0 9936 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 12052 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1618419204
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_108
timestamp 1618419204
transform 1 0 11040 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115
timestamp 1618419204
transform 1 0 11684 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_124
timestamp 1618419204
transform 1 0 12512 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen1
timestamp 1618419204
transform 1 0 14168 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_11_136
timestamp 1618419204
transform 1 0 13616 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_147
timestamp 1618419204
transform 1 0 14628 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1618419204
transform 1 0 14996 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1618419204
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_154
timestamp 1618419204
transform 1 0 15272 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_166
timestamp 1618419204
transform 1 0 16376 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_170
timestamp 1618419204
transform 1 0 16744 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_172
timestamp 1618419204
transform 1 0 16928 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1618419204
transform 1 0 19136 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen0
timestamp 1618419204
transform 1 0 17296 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb1
timestamp 1619507013
transform 1 0 18124 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_11_181
timestamp 1618419204
transform 1 0 17756 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_192
timestamp 1618419204
transform 1 0 18768 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1618419204
transform -1 0 21804 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1618419204
transform 1 0 20884 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_199
timestamp 1618419204
transform 1 0 19412 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_211
timestamp 1618419204
transform 1 0 20516 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_218
timestamp 1618419204
transform 1 0 21160 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1618419204
transform 1 0 2668 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1618419204
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1618419204
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_15
timestamp 1618419204
transform 1 0 2484 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1618419204
transform 1 0 2944 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 4508 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _372_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 6440 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1618419204
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_28
timestamp 1618419204
transform 1 0 3680 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_30
timestamp 1618419204
transform 1 0 3864 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_36
timestamp 1618419204
transform 1 0 4416 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_43
timestamp 1618419204
transform 1 0 5060 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 6808 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 8188 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_58
timestamp 1618419204
transform 1 0 6440 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_69
timestamp 1618419204
transform 1 0 7452 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _321_
timestamp 1619507013
transform -1 0 10028 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1618419204
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_77
timestamp 1618419204
transform 1 0 8188 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1618419204
transform 1 0 8924 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1618419204
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1618419204
transform 1 0 10028 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0
timestamp 1618419204
transform 1 0 11408 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1618419204
transform 1 0 12144 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_109
timestamp 1618419204
transform 1 0 11132 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_116
timestamp 1618419204
transform 1 0 11776 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_123
timestamp 1618419204
transform 1 0 12420 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1618419204
transform 1 0 14812 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1618419204
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_135
timestamp 1618419204
transform 1 0 13524 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_144
timestamp 1618419204
transform 1 0 14352 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_148
timestamp 1618419204
transform 1 0 14720 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb0
timestamp 1619507013
transform 1 0 16192 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_12_158
timestamp 1618419204
transform 1 0 15640 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_171
timestamp 1618419204
transform 1 0 16836 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1618419204
transform 1 0 17204 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen1
timestamp 1618419204
transform 1 0 18216 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_12_179
timestamp 1618419204
transform 1 0 17572 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_185
timestamp 1618419204
transform 1 0 18124 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_191
timestamp 1618419204
transform 1 0 18676 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1618419204
transform -1 0 21804 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1618419204
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_199
timestamp 1618419204
transform 1 0 19412 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1618419204
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_213
timestamp 1618419204
transform 1 0 20700 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_221
timestamp 1618419204
transform 1 0 21436 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1618419204
transform 1 0 1748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1618419204
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1618419204
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1618419204
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1618419204
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb1
timestamp 1619507013
transform 1 0 1748 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen1
timestamp 1618419204
transform 1 0 1840 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_13_14
timestamp 1618419204
transform 1 0 2392 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1618419204
transform 1 0 2760 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_13
timestamp 1618419204
transform 1 0 2300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_21
timestamp 1618419204
transform 1 0 3036 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _354_
timestamp 1618419204
transform -1 0 5888 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _377_
timestamp 1618419204
transform -1 0 5428 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1618419204
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_33
timestamp 1618419204
transform 1 0 4140 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_37
timestamp 1618419204
transform 1 0 4508 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1618419204
transform 1 0 5428 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_25
timestamp 1618419204
transform 1 0 3404 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1618419204
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_42
timestamp 1618419204
transform 1 0 4968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_52
timestamp 1618419204
transform 1 0 5888 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_58
timestamp 1618419204
transform 1 0 6440 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_55
timestamp 1618419204
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1618419204
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1618419204
transform 1 0 6256 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_72
timestamp 1618419204
transform 1 0 7728 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1618419204
transform 1 0 7084 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_66
timestamp 1618419204
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1619507013
transform -1 0 7728 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_8  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 8832 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__o21a_1  _312_
timestamp 1619507013
transform -1 0 10212 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _319_
timestamp 1619507013
transform 1 0 8096 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1618419204
transform -1 0 10212 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1618419204
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_84
timestamp 1618419204
transform 1 0 8832 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_99
timestamp 1618419204
transform 1 0 10212 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_82
timestamp 1618419204
transform 1 0 8648 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_87
timestamp 1618419204
transform 1 0 9108 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_99
timestamp 1618419204
transform 1 0 10212 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen1
timestamp 1618419204
transform 1 0 11500 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb1
timestamp 1619507013
transform 1 0 12052 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1618419204
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_111
timestamp 1618419204
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1618419204
transform 1 0 11684 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_111
timestamp 1618419204
transform 1 0 11316 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_118
timestamp 1618419204
transform 1 0 11960 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_135
timestamp 1618419204
transform 1 0 13524 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_126
timestamp 1618419204
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_133
timestamp 1618419204
transform 1 0 13340 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_126
timestamp 1618419204
transform 1 0 12696 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 1618419204
transform 1 0 13064 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb0
timestamp 1619507013
transform 1 0 12880 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_13_141
timestamp 1618419204
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1618419204
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _347_
timestamp 1618419204
transform -1 0 14536 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_144
timestamp 1618419204
transform 1 0 14352 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_146
timestamp 1618419204
transform 1 0 14536 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1618419204
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_158
timestamp 1618419204
transform 1 0 15640 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_170
timestamp 1618419204
transform 1 0 16744 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1618419204
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_156
timestamp 1618419204
transform 1 0 15456 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_168
timestamp 1618419204
transform 1 0 16560 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen1
timestamp 1618419204
transform -1 0 18676 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb1
timestamp 1619507013
transform -1 0 17848 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1618419204
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1618419204
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_174
timestamp 1618419204
transform 1 0 17112 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_182
timestamp 1618419204
transform 1 0 17848 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_191
timestamp 1618419204
transform 1 0 18676 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_199
timestamp 1618419204
transform 1 0 19412 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1618419204
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_218
timestamp 1618419204
transform 1 0 21160 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_213
timestamp 1618419204
transform 1 0 20700 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_220
timestamp 1618419204
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1618419204
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1618419204
transform -1 0 21804 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1618419204
transform -1 0 21804 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1618419204
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1618419204
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1618419204
transform 1 0 2576 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1618419204
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output39
timestamp 1618419204
transform -1 0 1748 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_7
timestamp 1618419204
transform 1 0 1748 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_15
timestamp 1618419204
transform 1 0 2484 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_20
timestamp 1618419204
transform 1 0 2944 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _314_
timestamp 1619507013
transform 1 0 4600 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_32
timestamp 1618419204
transform 1 0 4048 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1618419204
transform 1 0 5152 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _300_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 7728 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1618419204
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_56
timestamp 1618419204
transform 1 0 6256 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_58
timestamp 1618419204
transform 1 0 6440 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_66
timestamp 1618419204
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_72
timestamp 1618419204
transform 1 0 7728 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1619507013
transform 1 0 9568 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  repeater46
timestamp 1619507013
transform -1 0 9200 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_78
timestamp 1618419204
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_88
timestamp 1618419204
transform 1 0 9200 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_95
timestamp 1618419204
transform 1 0 9844 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1618419204
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_107
timestamp 1618419204
transform 1 0 10948 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1618419204
transform 1 0 11500 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_115
timestamp 1618419204
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen0
timestamp 1618419204
transform 1 0 13064 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb0
timestamp 1619507013
transform 1 0 14812 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_15_127
timestamp 1618419204
transform 1 0 12788 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1618419204
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_147
timestamp 1618419204
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen0
timestamp 1618419204
transform 1 0 15824 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1618419204
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_156
timestamp 1618419204
transform 1 0 15456 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_165
timestamp 1618419204
transform 1 0 16284 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_172
timestamp 1618419204
transform 1 0 16928 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp 1618419204
transform 1 0 17664 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _385_
timestamp 1619507013
transform 1 0 19136 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_15_189
timestamp 1618419204
transform 1 0 18492 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_195
timestamp 1618419204
transform 1 0 19044 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1618419204
transform -1 0 21804 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_217
timestamp 1618419204
transform 1 0 21068 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_221
timestamp 1618419204
transform 1 0 21436 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1618419204
transform 1 0 1564 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen1
timestamp 1618419204
transform -1 0 3404 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1618419204
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1618419204
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_14
timestamp 1618419204
transform 1 0 2392 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1618419204
transform 1 0 4232 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1618419204
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_25
timestamp 1618419204
transform 1 0 3404 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_30
timestamp 1618419204
transform 1 0 3864 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_37
timestamp 1618419204
transform 1 0 4508 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_49
timestamp 1618419204
transform 1 0 5612 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1619507013
transform 1 0 6900 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 7544 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 5888 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_16_59
timestamp 1618419204
transform 1 0 6532 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_66
timestamp 1618419204
transform 1 0 7176 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _315_
timestamp 1619507013
transform 1 0 10028 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1618419204
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_77
timestamp 1618419204
transform 1 0 8188 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1618419204
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_87
timestamp 1618419204
transform 1 0 9108 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_95
timestamp 1618419204
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_2  _365_
timestamp 1618419204
transform 1 0 11224 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_102
timestamp 1618419204
transform 1 0 10488 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_119
timestamp 1618419204
transform 1 0 12052 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1618419204
transform -1 0 13432 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1618419204
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_134
timestamp 1618419204
transform 1 0 13432 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_142
timestamp 1618419204
transform 1 0 14168 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_144
timestamp 1618419204
transform 1 0 14352 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1618419204
transform 1 0 14904 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1618419204
transform -1 0 17020 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1618419204
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1618419204
transform 1 0 16376 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_173
timestamp 1618419204
transform 1 0 17020 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _373_
timestamp 1618419204
transform 1 0 18032 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1618419204
transform -1 0 17664 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_180
timestamp 1618419204
transform 1 0 17664 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_193
timestamp 1618419204
transform 1 0 18860 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1618419204
transform -1 0 20332 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1618419204
transform -1 0 21804 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1618419204
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_199
timestamp 1618419204
transform 1 0 19412 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_201
timestamp 1618419204
transform 1 0 19596 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_205
timestamp 1618419204
transform 1 0 19964 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1618419204
transform 1 0 20332 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_221
timestamp 1618419204
transform 1 0 21436 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb1
timestamp 1619507013
transform -1 0 3588 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1618419204
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1618419204
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 1618419204
transform 1 0 2484 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_19
timestamp 1618419204
transform 1 0 2852 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _308_
timestamp 1618419204
transform 1 0 5336 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1618419204
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_39
timestamp 1618419204
transform 1 0 4692 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_45
timestamp 1618419204
transform 1 0 5244 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _296_
timestamp 1618419204
transform -1 0 7268 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _298_
timestamp 1618419204
transform -1 0 8464 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1618419204
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_53
timestamp 1618419204
transform 1 0 5980 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_58
timestamp 1618419204
transform 1 0 6440 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_67
timestamp 1618419204
transform 1 0 7268 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _311_
timestamp 1619507013
transform 1 0 9292 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_80
timestamp 1618419204
transform 1 0 8464 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_88
timestamp 1618419204
transform 1 0 9200 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_98
timestamp 1618419204
transform 1 0 10120 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _317_
timestamp 1619507013
transform -1 0 11040 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1618419204
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_108
timestamp 1618419204
transform 1 0 11040 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_115
timestamp 1618419204
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_127
timestamp 1618419204
transform 1 0 12788 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_139
timestamp 1618419204
transform 1 0 13892 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1618419204
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_151
timestamp 1618419204
transform 1 0 14996 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_163
timestamp 1618419204
transform 1 0 16100 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_172
timestamp 1618419204
transform 1 0 16928 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1618419204
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1618419204
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1618419204
transform -1 0 21804 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1618419204
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_220
timestamp 1618419204
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1618419204
transform 1 0 3128 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1618419204
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1618419204
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_15
timestamp 1618419204
transform 1 0 2484 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_21
timestamp 1618419204
transform 1 0 3036 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _366_
timestamp 1618419204
transform 1 0 4968 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1618419204
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_25
timestamp 1618419204
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1618419204
transform 1 0 3864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _302_
timestamp 1618419204
transform 1 0 7544 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _304_
timestamp 1618419204
transform 1 0 6164 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_18_51
timestamp 1618419204
transform 1 0 5796 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_62
timestamp 1618419204
transform 1 0 6808 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_74
timestamp 1618419204
transform 1 0 7912 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1618419204
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1618419204
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_99
timestamp 1618419204
transform 1 0 10212 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1618419204
transform -1 0 12328 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_111
timestamp 1618419204
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_122
timestamp 1618419204
transform 1 0 12328 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _292_
timestamp 1618419204
transform 1 0 12696 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1618419204
transform -1 0 14996 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1618419204
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_131
timestamp 1618419204
transform 1 0 13156 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_144
timestamp 1618419204
transform 1 0 14352 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_151
timestamp 1618419204
transform 1 0 14996 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_163
timestamp 1618419204
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_175
timestamp 1618419204
transform 1 0 17204 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_187
timestamp 1618419204
transform 1 0 18308 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1618419204
transform 1 0 20608 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1618419204
transform -1 0 21804 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1618419204
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_199
timestamp 1618419204
transform 1 0 19412 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_201
timestamp 1618419204
transform 1 0 19596 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_209
timestamp 1618419204
transform 1 0 20332 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_215
timestamp 1618419204
transform 1 0 20884 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_221
timestamp 1618419204
transform 1 0 21436 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1618419204
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_7
timestamp 1618419204
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output40
timestamp 1618419204
transform -1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1618419204
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1618419204
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb0
timestamp 1619507013
transform 1 0 2116 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _364_
timestamp 1618419204
transform -1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_18
timestamp 1618419204
transform 1 0 2760 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen0
timestamp 1618419204
transform 1 0 3128 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_20_14
timestamp 1618419204
transform 1 0 2392 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_1  _293_
timestamp 1618419204
transform -1 0 5336 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1618419204
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1618419204
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_39
timestamp 1618419204
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_46
timestamp 1618419204
transform 1 0 5336 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_26
timestamp 1618419204
transform 1 0 3496 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1618419204
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_42
timestamp 1618419204
transform 1 0 4968 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _248_
timestamp 1618419204
transform 1 0 6072 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1619507013
transform 1 0 7268 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _254_
timestamp 1618419204
transform 1 0 7544 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1618419204
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_54
timestamp 1618419204
transform 1 0 6072 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1618419204
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_59
timestamp 1618419204
transform 1 0 6532 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_70
timestamp 1618419204
transform 1 0 7544 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_80
timestamp 1618419204
transform 1 0 8464 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_76
timestamp 1618419204
transform 1 0 8096 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_86
timestamp 1618419204
transform 1 0 9016 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_77
timestamp 1618419204
transform 1 0 8188 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1618419204
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _310_
timestamp 1619507013
transform -1 0 9016 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1619507013
transform 1 0 8188 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_87
timestamp 1618419204
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_92
timestamp 1618419204
transform 1 0 9568 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o41a_1  _316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 10488 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _309_
timestamp 1618419204
transform 1 0 9476 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_20_96
timestamp 1618419204
transform 1 0 9936 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_109
timestamp 1618419204
transform 1 0 11132 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_102
timestamp 1618419204
transform 1 0 10488 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 11132 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _290_
timestamp 1618419204
transform 1 0 11040 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_20_117
timestamp 1618419204
transform 1 0 11868 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_113
timestamp 1618419204
transform 1 0 11500 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_115
timestamp 1618419204
transform 1 0 11684 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1618419204
transform 1 0 11500 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1618419204
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _371_
timestamp 1618419204
transform -1 0 12788 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1618419204
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1618419204
transform 1 0 12604 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _401_
timestamp 1619507013
transform 1 0 13800 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1618419204
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1618419204
transform 1 0 13432 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_127
timestamp 1618419204
transform 1 0 12788 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_139
timestamp 1618419204
transform 1 0 13892 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1618419204
transform 1 0 14352 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _341_
timestamp 1618419204
transform -1 0 16468 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _386_
timestamp 1619507013
transform -1 0 17756 0 -1 13600
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1618419204
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_158
timestamp 1618419204
transform 1 0 15640 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_167
timestamp 1618419204
transform 1 0 16468 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_172
timestamp 1618419204
transform 1 0 16928 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_156
timestamp 1618419204
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_181
timestamp 1618419204
transform 1 0 17756 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_180
timestamp 1618419204
transform 1 0 17664 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _285_
timestamp 1618419204
transform -1 0 17664 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _279_
timestamp 1618419204
transform -1 0 18584 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_20_198
timestamp 1618419204
transform 1 0 19320 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_190
timestamp 1618419204
transform 1 0 18584 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_194
timestamp 1618419204
transform 1 0 18952 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_188
timestamp 1618419204
transform 1 0 18400 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _288_
timestamp 1618419204
transform 1 0 18492 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _400_
timestamp 1619507013
transform 1 0 19320 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__a22o_1  _200_
timestamp 1619507013
transform -1 0 20608 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1618419204
transform -1 0 21804 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1618419204
transform -1 0 21804 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1618419204
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_218
timestamp 1618419204
transform 1 0 21160 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_201
timestamp 1618419204
transform 1 0 19596 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_212
timestamp 1618419204
transform 1 0 20608 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_220
timestamp 1618419204
transform 1 0 21344 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1618419204
transform -1 0 3496 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1618419204
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1618419204
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_15
timestamp 1618419204
transform 1 0 2484 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_21
timestamp 1618419204
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_26
timestamp 1618419204
transform 1 0 3496 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_38
timestamp 1618419204
transform 1 0 4600 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _294_
timestamp 1618419204
transform 1 0 7820 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _305_
timestamp 1618419204
transform 1 0 6808 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1618419204
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_50
timestamp 1618419204
transform 1 0 5704 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_56
timestamp 1618419204
transform 1 0 6256 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_58
timestamp 1618419204
transform 1 0 6440 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_69
timestamp 1618419204
transform 1 0 7452 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1619507013
transform 1 0 8648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _320_
timestamp 1618419204
transform -1 0 10304 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_78
timestamp 1618419204
transform 1 0 8280 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_85
timestamp 1618419204
transform 1 0 8924 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 12052 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1618419204
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_100
timestamp 1618419204
transform 1 0 10304 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_112
timestamp 1618419204
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_115
timestamp 1618419204
transform 1 0 11684 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_124
timestamp 1618419204
transform 1 0 12512 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _199_
timestamp 1619507013
transform -1 0 14720 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_21_136
timestamp 1618419204
transform 1 0 13616 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_140
timestamp 1618419204
transform 1 0 13984 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_148
timestamp 1618419204
transform 1 0 14720 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1618419204
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1618419204
transform 1 0 15824 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_168
timestamp 1618419204
transform 1 0 16560 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_172
timestamp 1618419204
transform 1 0 16928 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _286_
timestamp 1618419204
transform 1 0 17296 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 19320 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_21_183
timestamp 1618419204
transform 1 0 17940 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_198
timestamp 1618419204
transform 1 0 19320 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1618419204
transform -1 0 21804 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1619507013
transform -1 0 21160 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_210
timestamp 1618419204
transform 1 0 20424 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_214
timestamp 1618419204
transform 1 0 20792 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_218
timestamp 1618419204
transform 1 0 21160 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1618419204
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1618419204
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1618419204
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  _392_
timestamp 1619507013
transform -1 0 6164 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1618419204
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1618419204
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_30
timestamp 1618419204
transform 1 0 3864 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1619507013
transform 1 0 7360 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1619507013
transform 1 0 6532 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_55
timestamp 1618419204
transform 1 0 6164 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_62
timestamp 1618419204
transform 1 0 6808 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_71
timestamp 1618419204
transform 1 0 7636 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1618419204
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_83
timestamp 1618419204
transform 1 0 8740 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_87
timestamp 1618419204
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1618419204
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_4  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 12328 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_22_111
timestamp 1618419204
transform 1 0 11316 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_119
timestamp 1618419204
transform 1 0 12052 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 14720 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1618419204
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1618419204
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1618419204
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_144
timestamp 1618419204
transform 1 0 14352 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1619507013
transform -1 0 16100 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_156
timestamp 1618419204
transform 1 0 15456 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_163
timestamp 1618419204
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1619507013
transform 1 0 17296 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1619507013
transform -1 0 19044 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1619507013
transform -1 0 18216 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_175
timestamp 1618419204
transform 1 0 17204 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_179
timestamp 1618419204
transform 1 0 17572 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_186
timestamp 1618419204
transform 1 0 18216 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_195
timestamp 1618419204
transform 1 0 19044 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _209_
timestamp 1618419204
transform 1 0 20148 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1618419204
transform -1 0 21804 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1618419204
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_199
timestamp 1618419204
transform 1 0 19412 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_201
timestamp 1618419204
transform 1 0 19596 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_215
timestamp 1618419204
transform 1 0 20884 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_221
timestamp 1618419204
transform 1 0 21436 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1618419204
transform 1 0 1564 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb1
timestamp 1619507013
transform -1 0 3496 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1618419204
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1618419204
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_14
timestamp 1618419204
transform 1 0 2392 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_18
timestamp 1618419204
transform 1 0 2760 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1618419204
transform 1 0 4876 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen1
timestamp 1618419204
transform 1 0 3864 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_23_26
timestamp 1618419204
transform 1 0 3496 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_35
timestamp 1618419204
transform 1 0 4324 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_44
timestamp 1618419204
transform 1 0 5152 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _246_
timestamp 1619507013
transform 1 0 6808 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1618419204
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_56
timestamp 1618419204
transform 1 0 6256 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_58
timestamp 1618419204
transform 1 0 6440 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1618419204
transform 1 0 7452 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _363_
timestamp 1618419204
transform 1 0 9384 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1618419204
transform 1 0 8556 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_89
timestamp 1618419204
transform 1 0 9292 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_99
timestamp 1618419204
transform 1 0 10212 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1619507013
transform 1 0 10580 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1618419204
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_106
timestamp 1618419204
transform 1 0 10856 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_115
timestamp 1618419204
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _223_
timestamp 1619507013
transform 1 0 14260 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 13064 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_127
timestamp 1618419204
transform 1 0 12788 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1618419204
transform 1 0 13800 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_142
timestamp 1618419204
transform 1 0 14168 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_147
timestamp 1618419204
transform 1 0 14628 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _207_
timestamp 1619507013
transform -1 0 15272 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1618419204
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_154
timestamp 1618419204
transform 1 0 15272 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_166
timestamp 1618419204
transform 1 0 16376 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_170
timestamp 1618419204
transform 1 0 16744 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_172
timestamp 1618419204
transform 1 0 16928 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1619507013
transform 1 0 18860 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_184
timestamp 1618419204
transform 1 0 18032 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_192
timestamp 1618419204
transform 1 0 18768 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_196
timestamp 1618419204
transform 1 0 19136 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _210_
timestamp 1619507013
transform -1 0 20240 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1618419204
transform -1 0 21804 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1619507013
transform -1 0 21160 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_200
timestamp 1618419204
transform 1 0 19504 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_208
timestamp 1618419204
transform 1 0 20240 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_214
timestamp 1618419204
transform 1 0 20792 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_218
timestamp 1618419204
transform 1 0 21160 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1619507013
transform 1 0 2024 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1618419204
transform -1 0 3312 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1618419204
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1618419204
transform -1 0 1656 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_6
timestamp 1618419204
transform 1 0 1656 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_17
timestamp 1618419204
transform 1 0 2668 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1618419204
transform 1 0 3312 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1618419204
transform 1 0 4232 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1618419204
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_28
timestamp 1618419204
transform 1 0 3680 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_30
timestamp 1618419204
transform 1 0 3864 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_37
timestamp 1618419204
transform 1 0 4508 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_49
timestamp 1618419204
transform 1 0 5612 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1619507013
transform 1 0 6992 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _273_
timestamp 1618419204
transform -1 0 6624 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_55
timestamp 1618419204
transform 1 0 6164 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_60
timestamp 1618419204
transform 1 0 6624 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_67
timestamp 1618419204
transform 1 0 7268 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _258_
timestamp 1619507013
transform -1 0 8648 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_2  _395_
timestamp 1619507013
transform 1 0 9936 0 -1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1618419204
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_82
timestamp 1618419204
transform 1 0 8648 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_87
timestamp 1618419204
transform 1 0 9108 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_95
timestamp 1618419204
transform 1 0 9844 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _221_
timestamp 1618419204
transform 1 0 12328 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_24_117
timestamp 1618419204
transform 1 0 11868 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_121
timestamp 1618419204
transform 1 0 12236 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _220_
timestamp 1618419204
transform 1 0 13156 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1618419204
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_127
timestamp 1618419204
transform 1 0 12788 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_139
timestamp 1618419204
transform 1 0 13892 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_144
timestamp 1618419204
transform 1 0 14352 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 16928 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_24_156
timestamp 1618419204
transform 1 0 15456 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_168
timestamp 1618419204
transform 1 0 16560 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_179
timestamp 1618419204
transform 1 0 17572 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_191
timestamp 1618419204
transform 1 0 18676 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2ai_1  _228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 20608 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1618419204
transform -1 0 21804 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1618419204
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_199
timestamp 1618419204
transform 1 0 19412 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_201
timestamp 1618419204
transform 1 0 19596 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_212
timestamp 1618419204
transform 1 0 20608 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_220
timestamp 1618419204
transform 1 0 21344 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb0
timestamp 1619507013
transform 1 0 1564 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1618419204
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1618419204
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_12
timestamp 1618419204
transform 1 0 2208 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_24
timestamp 1618419204
transform 1 0 3312 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_36
timestamp 1618419204
transform 1 0 4416 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_48
timestamp 1618419204
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1619507013
transform -1 0 5980 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 7544 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1618419204
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_53
timestamp 1618419204
transform 1 0 5980 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_58
timestamp 1618419204
transform 1 0 6440 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_70
timestamp 1618419204
transform 1 0 7544 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _260_
timestamp 1618419204
transform 1 0 8464 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _261_
timestamp 1618419204
transform -1 0 9936 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_78
timestamp 1618419204
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_88
timestamp 1618419204
transform 1 0 9200 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_96
timestamp 1618419204
transform 1 0 9936 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 12880 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1618419204
transform -1 0 11224 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1618419204
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_104
timestamp 1618419204
transform 1 0 10672 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_110
timestamp 1618419204
transform 1 0 11224 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_115
timestamp 1618419204
transform 1 0 11684 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1618419204
transform 1 0 12052 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _213_
timestamp 1618419204
transform -1 0 15180 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_128
timestamp 1618419204
transform 1 0 12880 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 1618419204
transform 1 0 13984 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_144
timestamp 1618419204
transform 1 0 14352 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _206_
timestamp 1619507013
transform 1 0 15548 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1618419204
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1618419204
transform 1 0 15180 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 1618419204
transform 1 0 15824 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_168
timestamp 1618419204
transform 1 0 16560 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_172
timestamp 1618419204
transform 1 0 16928 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _384_
timestamp 1619507013
transform 1 0 17296 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_25_196
timestamp 1618419204
transform 1 0 19136 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _208_
timestamp 1619507013
transform 1 0 20424 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _227_
timestamp 1618419204
transform -1 0 20056 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1618419204
transform -1 0 21804 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1618419204
transform 1 0 20056 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_215
timestamp 1618419204
transform 1 0 20884 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_221
timestamp 1618419204
transform 1 0 21436 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1618419204
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1618419204
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1618419204
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1618419204
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1618419204
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1618419204
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _244_
timestamp 1619507013
transform 1 0 5336 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1618419204
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1618419204
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1618419204
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_42
timestamp 1618419204
transform 1 0 4968 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1618419204
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_39
timestamp 1618419204
transform 1 0 4692 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_45
timestamp 1618419204
transform 1 0 5244 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_58
timestamp 1618419204
transform 1 0 6440 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_53
timestamp 1618419204
transform 1 0 5980 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_55
timestamp 1618419204
transform 1 0 6164 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_50
timestamp 1618419204
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1618419204
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _270_
timestamp 1618419204
transform 1 0 5796 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _250_
timestamp 1619507013
transform -1 0 7544 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1619507013
transform 1 0 6532 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_70
timestamp 1618419204
transform 1 0 7544 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_74
timestamp 1618419204
transform 1 0 7912 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_62
timestamp 1618419204
transform 1 0 6808 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1618419204
transform 1 0 8924 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_79
timestamp 1618419204
transform 1 0 8372 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1618419204
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1619507013
transform -1 0 8372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1619507013
transform 1 0 8096 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_97
timestamp 1618419204
transform 1 0 10028 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_91
timestamp 1618419204
transform 1 0 9476 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1619507013
transform 1 0 10120 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_79
timestamp 1618419204
transform 1 0 8372 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_99
timestamp 1618419204
transform 1 0 10212 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1618419204
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1619507013
transform 1 0 12144 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_2  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 12052 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1618419204
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_111
timestamp 1618419204
transform 1 0 11316 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_119
timestamp 1618419204
transform 1 0 12052 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_123
timestamp 1618419204
transform 1 0 12420 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_101
timestamp 1618419204
transform 1 0 10396 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1618419204
transform 1 0 11500 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_115
timestamp 1618419204
transform 1 0 11684 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _219_
timestamp 1618419204
transform 1 0 14720 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _402_
timestamp 1619507013
transform -1 0 16284 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1618419204
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_135
timestamp 1618419204
transform 1 0 13524 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_144
timestamp 1618419204
transform 1 0 14352 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_131
timestamp 1618419204
transform 1 0 13156 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_143
timestamp 1618419204
transform 1 0 14260 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__a311o_1  _289_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 17572 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1618419204
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1618419204
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_166
timestamp 1618419204
transform 1 0 16376 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_170
timestamp 1618419204
transform 1 0 16744 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_165
timestamp 1618419204
transform 1 0 16284 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1618419204
transform 1 0 16928 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1619507013
transform -1 0 19136 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _343_
timestamp 1618419204
transform -1 0 18216 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _399_
timestamp 1619507013
transform 1 0 19320 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_26_179
timestamp 1618419204
transform 1 0 17572 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_186
timestamp 1618419204
transform 1 0 18216 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_192
timestamp 1618419204
transform 1 0 18768 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_196
timestamp 1618419204
transform 1 0 19136 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1618419204
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_196
timestamp 1618419204
transform 1 0 19136 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _201_
timestamp 1619507013
transform 1 0 19964 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1618419204
transform -1 0 21804 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1618419204
transform -1 0 21804 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1618419204
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_201
timestamp 1618419204
transform 1 0 19596 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_212
timestamp 1618419204
transform 1 0 20608 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_220
timestamp 1618419204
transform 1 0 21344 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_218
timestamp 1618419204
transform 1 0 21160 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1618419204
transform -1 0 3404 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1618419204
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1618419204
transform -1 0 1656 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_6
timestamp 1618419204
transform 1 0 1656 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_18
timestamp 1618419204
transform 1 0 2760 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 4600 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1618419204
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_25
timestamp 1618419204
transform 1 0 3404 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_30
timestamp 1618419204
transform 1 0 3864 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_46
timestamp 1618419204
transform 1 0 5336 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1619507013
transform 1 0 6808 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _256_
timestamp 1619507013
transform 1 0 7820 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _269_
timestamp 1618419204
transform -1 0 6440 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_28_52
timestamp 1618419204
transform 1 0 5888 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_58
timestamp 1618419204
transform 1 0 6440 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_65
timestamp 1618419204
transform 1 0 7084 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _394_
timestamp 1619507013
transform 1 0 9476 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1618419204
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_81
timestamp 1618419204
transform 1 0 8556 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 1618419204
transform 1 0 8924 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_87
timestamp 1618419204
transform 1 0 9108 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _237_
timestamp 1618419204
transform 1 0 12236 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_28_112
timestamp 1618419204
transform 1 0 11408 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_120
timestamp 1618419204
transform 1 0 12144 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _198_
timestamp 1619507013
transform 1 0 14720 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1619507013
transform 1 0 13064 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1618419204
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_126
timestamp 1618419204
transform 1 0 12696 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_133
timestamp 1618419204
transform 1 0 13340 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1618419204
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_144
timestamp 1618419204
transform 1 0 14352 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_155
timestamp 1618419204
transform 1 0 15364 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_167
timestamp 1618419204
transform 1 0 16468 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_179
timestamp 1618419204
transform 1 0 17572 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_191
timestamp 1618419204
transform 1 0 18676 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp 1618419204
transform 1 0 20700 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1618419204
transform -1 0 21804 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1618419204
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_199
timestamp 1618419204
transform 1 0 19412 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_201
timestamp 1618419204
transform 1 0 19596 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_216
timestamp 1618419204
transform 1 0 20976 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_2  _391_
timestamp 1619507013
transform -1 0 4600 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1618419204
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1618419204
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_15
timestamp 1618419204
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  _274_
timestamp 1618419204
transform -1 0 5704 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_29_38
timestamp 1618419204
transform 1 0 4600 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_44
timestamp 1618419204
transform 1 0 5152 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1618419204
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1618419204
transform 1 0 5704 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_56
timestamp 1618419204
transform 1 0 6256 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_58
timestamp 1618419204
transform 1 0 6440 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_70
timestamp 1618419204
transform 1 0 7544 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _252_
timestamp 1619507013
transform 1 0 8464 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _266_
timestamp 1618419204
transform -1 0 9844 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 1618419204
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_87
timestamp 1618419204
transform 1 0 9108 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_95
timestamp 1618419204
transform 1 0 9844 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_99
timestamp 1618419204
transform 1 0 10212 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _238_
timestamp 1619507013
transform 1 0 12144 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp 1618419204
transform -1 0 10580 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1618419204
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_103
timestamp 1618419204
transform 1 0 10580 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_111
timestamp 1618419204
transform 1 0 11316 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_115
timestamp 1618419204
transform 1 0 11684 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_119
timestamp 1618419204
transform 1 0 12052 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1618419204
transform 1 0 13708 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1618419204
transform 1 0 14812 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1618419204
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_161
timestamp 1618419204
transform 1 0 15916 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1618419204
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_172
timestamp 1618419204
transform 1 0 16928 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1619507013
transform -1 0 18676 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _231_
timestamp 1618419204
transform -1 0 19872 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1618419204
transform -1 0 17572 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_179
timestamp 1618419204
transform 1 0 17572 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_187
timestamp 1618419204
transform 1 0 18308 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_191
timestamp 1618419204
transform 1 0 18676 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1618419204
transform -1 0 21804 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1618419204
transform 1 0 20884 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_204
timestamp 1618419204
transform 1 0 19872 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_212
timestamp 1618419204
transform 1 0 20608 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_218
timestamp 1618419204
transform 1 0 21160 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1618419204
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1618419204
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1618419204
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _242_
timestamp 1618419204
transform -1 0 5704 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1618419204
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1618419204
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_30
timestamp 1618419204
transform 1 0 3864 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_42
timestamp 1618419204
transform 1 0 4968 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1619507013
transform 1 0 6532 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _263_
timestamp 1618419204
transform 1 0 7820 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_50
timestamp 1618419204
transform 1 0 5704 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_58
timestamp 1618419204
transform 1 0 6440 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_62
timestamp 1618419204
transform 1 0 6808 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_70
timestamp 1618419204
transform 1 0 7544 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1619507013
transform 1 0 9476 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1618419204
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_77
timestamp 1618419204
transform 1 0 8188 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1618419204
transform 1 0 8924 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_87
timestamp 1618419204
transform 1 0 9108 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_94
timestamp 1618419204
transform 1 0 9752 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__a41o_2  _234_
timestamp 1619507013
transform 1 0 12236 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_30_106
timestamp 1618419204
transform 1 0 10856 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_118
timestamp 1618419204
transform 1 0 11960 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _236_
timestamp 1618419204
transform -1 0 13800 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1618419204
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_130
timestamp 1618419204
transform 1 0 13064 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_138
timestamp 1618419204
transform 1 0 13800 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_142
timestamp 1618419204
transform 1 0 14168 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_144
timestamp 1618419204
transform 1 0 14352 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _283_
timestamp 1618419204
transform 1 0 15456 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_2  _387_
timestamp 1619507013
transform 1 0 16652 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_30_165
timestamp 1618419204
transform 1 0 16284 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_190
timestamp 1618419204
transform 1 0 18584 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_198
timestamp 1618419204
transform 1 0 19320 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _229_
timestamp 1618419204
transform -1 0 21160 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 19964 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1618419204
transform -1 0 21804 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1618419204
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_201
timestamp 1618419204
transform 1 0 19596 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_211
timestamp 1618419204
transform 1 0 20516 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_218
timestamp 1618419204
transform 1 0 21160 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1618419204
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1618419204
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1618419204
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1619507013
transform 1 0 4508 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _240_
timestamp 1619507013
transform 1 0 5152 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_31_27
timestamp 1618419204
transform 1 0 3588 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_35
timestamp 1618419204
transform 1 0 4324 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_40
timestamp 1618419204
transform 1 0 4784 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _251_
timestamp 1619507013
transform 1 0 7360 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1618419204
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_51
timestamp 1618419204
transform 1 0 5796 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_58
timestamp 1618419204
transform 1 0 6440 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_66
timestamp 1618419204
transform 1 0 7176 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1619507013
transform 1 0 9568 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _265_
timestamp 1618419204
transform 1 0 8464 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_75
timestamp 1618419204
transform 1 0 8004 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_79
timestamp 1618419204
transform 1 0 8372 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_88
timestamp 1618419204
transform 1 0 9200 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_95
timestamp 1618419204
transform 1 0 9844 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1619507013
transform -1 0 12788 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1618419204
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_107
timestamp 1618419204
transform 1 0 10948 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 1618419204
transform 1 0 11500 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_115
timestamp 1618419204
transform 1 0 11684 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_123
timestamp 1618419204
transform 1 0 12420 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _216_
timestamp 1618419204
transform -1 0 14996 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _218_
timestamp 1618419204
transform -1 0 13800 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_127
timestamp 1618419204
transform 1 0 12788 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_138
timestamp 1618419204
transform 1 0 13800 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _214_
timestamp 1618419204
transform 1 0 15364 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1618419204
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_151
timestamp 1618419204
transform 1 0 14996 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_160
timestamp 1618419204
transform 1 0 15824 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_168
timestamp 1618419204
transform 1 0 16560 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_172
timestamp 1618419204
transform 1 0 16928 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp 1618419204
transform -1 0 17848 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _383_
timestamp 1619507013
transform 1 0 19320 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_31_178
timestamp 1618419204
transform 1 0 17480 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_182
timestamp 1618419204
transform 1 0 17848 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_194
timestamp 1618419204
transform 1 0 18952 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1618419204
transform -1 0 21804 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_218
timestamp 1618419204
transform 1 0 21160 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1618419204
transform -1 0 3404 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1618419204
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1618419204
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_15
timestamp 1618419204
transform 1 0 2484 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_21
timestamp 1618419204
transform 1 0 3036 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_1  _277_
timestamp 1618419204
transform 1 0 4692 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1618419204
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_25
timestamp 1618419204
transform 1 0 3404 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_30
timestamp 1618419204
transform 1 0 3864 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_38
timestamp 1618419204
transform 1 0 4600 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_47
timestamp 1618419204
transform 1 0 5428 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _262_
timestamp 1618419204
transform 1 0 7728 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _276_
timestamp 1618419204
transform 1 0 5796 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1618419204
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_68
timestamp 1618419204
transform 1 0 7360 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1618419204
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_77
timestamp 1618419204
transform 1 0 8188 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_85
timestamp 1618419204
transform 1 0 8924 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_87
timestamp 1618419204
transform 1 0 9108 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_99
timestamp 1618419204
transform 1 0 10212 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1618419204
transform -1 0 10580 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_103
timestamp 1618419204
transform 1 0 10580 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_115
timestamp 1618419204
transform 1 0 11684 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_1  _215_
timestamp 1618419204
transform -1 0 15456 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1618419204
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_127
timestamp 1618419204
transform 1 0 12788 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_139
timestamp 1618419204
transform 1 0 13892 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_144
timestamp 1618419204
transform 1 0 14352 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _282_
timestamp 1619507013
transform -1 0 16468 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_156
timestamp 1618419204
transform 1 0 15456 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_162
timestamp 1618419204
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_167
timestamp 1618419204
transform 1 0 16468 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_179
timestamp 1618419204
transform 1 0 17572 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_191
timestamp 1618419204
transform 1 0 18676 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp 1618419204
transform 1 0 20424 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1618419204
transform -1 0 21804 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1618419204
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_199
timestamp 1618419204
transform 1 0 19412 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_201
timestamp 1618419204
transform 1 0 19596 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_209
timestamp 1618419204
transform 1 0 20332 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_213
timestamp 1618419204
transform 1 0 20700 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_221
timestamp 1618419204
transform 1 0 21436 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _390_
timestamp 1619507013
transform 1 0 2484 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1618419204
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1618419204
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1619507013
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_6
timestamp 1618419204
transform 1 0 1656 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_14
timestamp 1618419204
transform 1 0 2392 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1618419204
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1618419204
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1618419204
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_35
timestamp 1618419204
transform 1 0 4324 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1618419204
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_42
timestamp 1618419204
transform 1 0 4968 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_48
timestamp 1618419204
transform 1 0 5520 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_43
timestamp 1618419204
transform 1 0 5060 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _241_
timestamp 1618419204
transform 1 0 5244 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1619507013
transform -1 0 5428 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_47
timestamp 1618419204
transform 1 0 5428 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_30
timestamp 1618419204
transform 1 0 3864 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_59
timestamp 1618419204
transform 1 0 6532 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_56
timestamp 1618419204
transform 1 0 6256 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1618419204
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_74
timestamp 1618419204
transform 1 0 7912 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_65
timestamp 1618419204
transform 1 0 7084 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_70
timestamp 1618419204
transform 1 0 7544 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_1  _268_
timestamp 1618419204
transform 1 0 7176 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _267_
timestamp 1618419204
transform -1 0 7912 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1618419204
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_58
timestamp 1618419204
transform 1 0 6440 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1619507013
transform 1 0 8280 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _398_
timestamp 1619507013
transform 1 0 9384 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1618419204
transform 1 0 9016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_86
timestamp 1618419204
transform 1 0 9016 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_81
timestamp 1618419204
transform 1 0 8556 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_85
timestamp 1618419204
transform 1 0 8924 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_87
timestamp 1618419204
transform 1 0 9108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_99
timestamp 1618419204
transform 1 0 10212 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _202_
timestamp 1619507013
transform -1 0 12420 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform 1 0 12052 0 1 20128
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1618419204
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_110
timestamp 1618419204
transform 1 0 11224 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_115
timestamp 1618419204
transform 1 0 11684 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_111
timestamp 1618419204
transform 1 0 11316 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_115
timestamp 1618419204
transform 1 0 11684 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_123
timestamp 1618419204
transform 1 0 12420 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1619507013
transform -1 0 14352 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _195_
timestamp 1619507013
transform 1 0 14720 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _205_
timestamp 1619507013
transform 1 0 14720 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1618419204
transform 1 0 14260 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_129
timestamp 1618419204
transform 1 0 12972 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_144
timestamp 1618419204
transform 1 0 14352 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_135
timestamp 1618419204
transform 1 0 13524 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_144
timestamp 1618419204
transform 1 0 14352 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1619507013
transform -1 0 16008 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _388_
timestamp 1619507013
transform 1 0 16192 0 -1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1618419204
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_155
timestamp 1618419204
transform 1 0 15364 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_162
timestamp 1618419204
transform 1 0 16008 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_170
timestamp 1618419204
transform 1 0 16744 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_172
timestamp 1618419204
transform 1 0 16928 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_155
timestamp 1618419204
transform 1 0 15364 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_163
timestamp 1618419204
transform 1 0 16100 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _339_
timestamp 1618419204
transform 1 0 17296 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _382_
timestamp 1619507013
transform 1 0 19044 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_33_179
timestamp 1618419204
transform 1 0 17572 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1618419204
transform 1 0 18676 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_185
timestamp 1618419204
transform 1 0 18124 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_197
timestamp 1618419204
transform 1 0 19228 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1618419204
transform -1 0 21804 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1618419204
transform -1 0 21804 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1618419204
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output42
timestamp 1618419204
transform 1 0 20792 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_215
timestamp 1618419204
transform 1 0 20884 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_221
timestamp 1618419204
transform 1 0 21436 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_201
timestamp 1618419204
transform 1 0 19596 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1618419204
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_218
timestamp 1618419204
transform 1 0 21160 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _349_
timestamp 1618419204
transform 1 0 1748 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1618419204
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1618419204
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_10
timestamp 1618419204
transform 1 0 2024 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_22
timestamp 1618419204
transform 1 0 3128 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _389_
timestamp 1619507013
transform 1 0 3864 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _393_
timestamp 1619507013
transform 1 0 6808 0 1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1618419204
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_50
timestamp 1618419204
transform 1 0 5704 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_56
timestamp 1618419204
transform 1 0 6256 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_58
timestamp 1618419204
transform 1 0 6440 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _396_
timestamp 1619507013
transform 1 0 9108 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_35_83
timestamp 1618419204
transform 1 0 8740 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _397_
timestamp 1619507013
transform -1 0 13892 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1618419204
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_107
timestamp 1618419204
transform 1 0 10948 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 1618419204
transform 1 0 11500 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_115
timestamp 1618419204
transform 1 0 11684 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _403_
timestamp 1619507013
transform -1 0 16100 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_35_139
timestamp 1618419204
transform 1 0 13892 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1618419204
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_163
timestamp 1618419204
transform 1 0 16100 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_172
timestamp 1618419204
transform 1 0 16928 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _381_
timestamp 1619507013
transform 1 0 17388 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_35_176
timestamp 1618419204
transform 1 0 17296 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_197
timestamp 1618419204
transform 1 0 19228 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 21160 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1618419204
transform -1 0 21804 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_201
timestamp 1618419204
transform 1 0 19596 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_218
timestamp 1618419204
transform 1 0 21160 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1618419204
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1618419204
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1618419204
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _278_
timestamp 1619507013
transform 1 0 4784 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1618419204
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1618419204
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_30
timestamp 1618419204
transform 1 0 3864 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_38
timestamp 1618419204
transform 1 0 4600 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_47
timestamp 1618419204
transform 1 0 5428 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1618419204
transform -1 0 7820 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_59
timestamp 1618419204
transform 1 0 6532 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_67
timestamp 1618419204
transform 1 0 7268 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_73
timestamp 1618419204
transform 1 0 7820 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 1618419204
transform -1 0 10120 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1618419204
transform 1 0 9016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_85
timestamp 1618419204
transform 1 0 8924 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_87
timestamp 1618419204
transform 1 0 9108 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_98
timestamp 1618419204
transform 1 0 10120 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _203_
timestamp 1619507013
transform 1 0 11684 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _204_
timestamp 1618419204
transform -1 0 11132 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_36_109
timestamp 1618419204
transform 1 0 11132 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_122
timestamp 1618419204
transform 1 0 12328 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1618419204
transform 1 0 12696 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1618419204
transform 1 0 14260 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1618419204
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1618419204
transform 1 0 14076 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_144
timestamp 1618419204
transform 1 0 14352 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp 1618419204
transform 1 0 15180 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_152
timestamp 1618419204
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_156
timestamp 1618419204
transform 1 0 15456 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1618419204
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp 1618419204
transform -1 0 18584 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_180
timestamp 1618419204
transform 1 0 17664 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_186
timestamp 1618419204
transform 1 0 18216 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_190
timestamp 1618419204
transform 1 0 18584 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_198
timestamp 1618419204
transform 1 0 19320 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _345_
timestamp 1618419204
transform -1 0 20240 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1618419204
transform -1 0 21804 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1618419204
transform 1 0 19504 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1619507013
transform -1 0 21160 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_201
timestamp 1618419204
transform 1 0 19596 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_208
timestamp 1618419204
transform 1 0 20240 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_214
timestamp 1618419204
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_218
timestamp 1618419204
transform 1 0 21160 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1618419204
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1619507013
transform 1 0 2760 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1618419204
transform 1 0 2116 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output44
timestamp 1618419204
transform -1 0 1748 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_7
timestamp 1618419204
transform 1 0 1748 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_14
timestamp 1618419204
transform 1 0 2392 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_21
timestamp 1618419204
transform 1 0 3036 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _338_
timestamp 1618419204
transform -1 0 4968 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1618419204
transform 1 0 3772 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1619507013
transform 1 0 5336 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_30
timestamp 1618419204
transform 1 0 3864 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_38
timestamp 1618419204
transform 1 0 4600 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_42
timestamp 1618419204
transform 1 0 4968 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_49
timestamp 1618419204
transform 1 0 5612 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1618419204
transform 1 0 6440 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1619507013
transform 1 0 7820 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1619507013
transform -1 0 7176 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_57
timestamp 1618419204
transform 1 0 6348 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_59
timestamp 1618419204
transform 1 0 6532 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_66
timestamp 1618419204
transform 1 0 7176 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_72
timestamp 1618419204
transform 1 0 7728 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1618419204
transform 1 0 9108 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1619507013
transform 1 0 9660 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_76
timestamp 1618419204
transform 1 0 8096 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_84
timestamp 1618419204
transform 1 0 8832 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_88
timestamp 1618419204
transform 1 0 9200 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_92
timestamp 1618419204
transform 1 0 9568 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_96
timestamp 1618419204
transform 1 0 9936 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1618419204
transform 1 0 11776 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1618419204
transform 1 0 12236 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_108
timestamp 1618419204
transform 1 0 11040 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_117
timestamp 1618419204
transform 1 0 11868 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_124
timestamp 1618419204
transform 1 0 12512 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1618419204
transform 1 0 14444 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1619507013
transform 1 0 12880 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_131
timestamp 1618419204
transform 1 0 13156 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_143
timestamp 1618419204
transform 1 0 14260 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_146
timestamp 1618419204
transform 1 0 14536 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1619507013
transform -1 0 15180 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1619507013
transform -1 0 16744 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_153
timestamp 1618419204
transform 1 0 15180 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_165
timestamp 1618419204
transform 1 0 16284 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_170
timestamp 1618419204
transform 1 0 16744 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1618419204
transform 1 0 17112 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1619507013
transform -1 0 19412 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1618419204
transform 1 0 17940 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_175
timestamp 1618419204
transform 1 0 17204 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_186
timestamp 1618419204
transform 1 0 18216 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_194
timestamp 1618419204
transform 1 0 18952 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1618419204
transform -1 0 21804 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1618419204
transform 1 0 19780 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1618419204
transform -1 0 21160 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_199
timestamp 1618419204
transform 1 0 19412 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_204
timestamp 1618419204
transform 1 0 19872 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_212
timestamp 1618419204
transform 1 0 20608 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_218
timestamp 1618419204
transform 1 0 21160 0 1 22304
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 10208 800 10328 6 clockc
port 0 nsew signal tristate
rlabel metal3 s 0 12928 800 13048 6 clockd[0]
port 1 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 clockd[1]
port 2 nsew signal tristate
rlabel metal3 s 22179 20408 22979 20528 6 clockd[2]
port 3 nsew signal tristate
rlabel metal2 s 20718 0 20774 800 6 clockd[3]
port 4 nsew signal tristate
rlabel metal3 s 0 23128 800 23248 6 clockp[0]
port 5 nsew signal tristate
rlabel metal2 s 1858 0 1914 800 6 clockp[1]
port 6 nsew signal tristate
rlabel metal2 s 15658 0 15714 800 6 dco
port 7 nsew signal input
rlabel metal3 s 22179 15648 22979 15768 6 div[0]
port 8 nsew signal input
rlabel metal2 s 19798 24323 19854 25123 6 div[1]
port 9 nsew signal input
rlabel metal2 s 7838 24323 7894 25123 6 div[2]
port 10 nsew signal input
rlabel metal2 s 478 0 534 800 6 div[3]
port 11 nsew signal input
rlabel metal2 s 14738 24323 14794 25123 6 div[4]
port 12 nsew signal input
rlabel metal2 s 16578 24323 16634 25123 6 ext_trim[0]
port 13 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 ext_trim[10]
port 14 nsew signal input
rlabel metal2 s 2778 24323 2834 25123 6 ext_trim[11]
port 15 nsew signal input
rlabel metal3 s 22179 5448 22979 5568 6 ext_trim[12]
port 16 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 ext_trim[13]
port 17 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 ext_trim[14]
port 18 nsew signal input
rlabel metal3 s 22179 17688 22979 17808 6 ext_trim[15]
port 19 nsew signal input
rlabel metal2 s 4618 24323 4674 25123 6 ext_trim[16]
port 20 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 ext_trim[17]
port 21 nsew signal input
rlabel metal2 s 5998 24323 6054 25123 6 ext_trim[18]
port 22 nsew signal input
rlabel metal3 s 22179 10208 22979 10328 6 ext_trim[19]
port 23 nsew signal input
rlabel metal2 s 12898 24323 12954 25123 6 ext_trim[1]
port 24 nsew signal input
rlabel metal2 s 11518 24323 11574 25123 6 ext_trim[20]
port 25 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 ext_trim[21]
port 26 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 ext_trim[22]
port 27 nsew signal input
rlabel metal3 s 22179 23128 22979 23248 6 ext_trim[23]
port 28 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 ext_trim[24]
port 29 nsew signal input
rlabel metal2 s 9678 24323 9734 25123 6 ext_trim[25]
port 30 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 ext_trim[2]
port 31 nsew signal input
rlabel metal3 s 22179 8168 22979 8288 6 ext_trim[3]
port 32 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 ext_trim[4]
port 33 nsew signal input
rlabel metal3 s 22179 12928 22979 13048 6 ext_trim[5]
port 34 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 ext_trim[6]
port 35 nsew signal input
rlabel metal2 s 938 24323 994 25123 6 ext_trim[7]
port 36 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 ext_trim[8]
port 37 nsew signal input
rlabel metal3 s 22179 2728 22979 2848 6 ext_trim[9]
port 38 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 extclk_sel
port 39 nsew signal input
rlabel metal2 s 17958 24323 18014 25123 6 osc
port 40 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 reset
port 41 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 sel[0]
port 42 nsew signal input
rlabel metal2 s 21638 24323 21694 25123 6 sel[1]
port 43 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 sel[2]
port 44 nsew signal input
rlabel metal4 s 18194 2128 18514 22896 6 VPWR
port 45 nsew power bidirectional
rlabel metal4 s 11294 2128 11614 22896 6 VPWR
port 46 nsew power bidirectional
rlabel metal4 s 4394 2128 4714 22896 6 VPWR
port 47 nsew power bidirectional
rlabel metal5 s 1104 19195 21804 19515 6 VPWR
port 48 nsew power bidirectional
rlabel metal5 s 1104 12304 21804 12624 6 VPWR
port 49 nsew power bidirectional
rlabel metal5 s 1104 5413 21804 5733 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 14744 2128 15064 22896 6 VGND
port 51 nsew ground bidirectional
rlabel metal4 s 7844 2128 8164 22896 6 VGND
port 52 nsew ground bidirectional
rlabel metal5 s 1104 15749 21804 16069 6 VGND
port 53 nsew ground bidirectional
rlabel metal5 s 1104 8859 21804 9179 6 VGND
port 54 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 22979 25123
<< end >>
