magic
tech sky130A
magscale 1 2
timestamp 1623853968
<< obsli1 >>
rect 1104 2159 16836 17969
<< obsm1 >>
rect 474 2048 17098 18000
<< metal2 >>
rect 478 19371 534 20171
rect 2318 19371 2374 20171
rect 3698 19371 3754 20171
rect 5538 19371 5594 20171
rect 6918 19371 6974 20171
rect 8758 19371 8814 20171
rect 10138 19371 10194 20171
rect 11978 19371 12034 20171
rect 13818 19371 13874 20171
rect 15198 19371 15254 20171
rect 17038 19371 17094 20171
rect 478 0 534 800
rect 1858 0 1914 800
rect 3698 0 3754 800
rect 5078 0 5134 800
rect 6918 0 6974 800
rect 8298 0 8354 800
rect 10138 0 10194 800
rect 11518 0 11574 800
rect 13358 0 13414 800
rect 15198 0 15254 800
rect 16578 0 16634 800
<< obsm2 >>
rect 590 19315 2262 19371
rect 2430 19315 3642 19371
rect 3810 19315 5482 19371
rect 5650 19315 6862 19371
rect 7030 19315 8702 19371
rect 8870 19315 10082 19371
rect 10250 19315 11922 19371
rect 12090 19315 13762 19371
rect 13930 19315 15142 19371
rect 15310 19315 16982 19371
rect 480 856 17092 19315
rect 590 800 1802 856
rect 1970 800 3642 856
rect 3810 800 5022 856
rect 5190 800 6862 856
rect 7030 800 8242 856
rect 8410 800 10082 856
rect 10250 800 11462 856
rect 11630 800 13302 856
rect 13470 800 15142 856
rect 15310 800 16522 856
rect 16690 800 17092 856
<< metal3 >>
rect 17227 18368 18027 18488
rect 0 17008 800 17128
rect 17227 15648 18027 15768
rect 0 14968 800 15088
rect 17227 13608 18027 13728
rect 0 12248 800 12368
rect 17227 10888 18027 11008
rect 0 10208 800 10328
rect 17227 8168 18027 8288
rect 0 7488 800 7608
rect 17227 6128 18027 6248
rect 0 5448 800 5568
rect 17227 3408 18027 3528
rect 0 2728 800 2848
rect 17227 1368 18027 1488
<< obsm3 >>
rect 800 18288 17147 18461
rect 800 17208 17227 18288
rect 880 16928 17227 17208
rect 800 15848 17227 16928
rect 800 15568 17147 15848
rect 800 15168 17227 15568
rect 880 14888 17227 15168
rect 800 13808 17227 14888
rect 800 13528 17147 13808
rect 800 12448 17227 13528
rect 880 12168 17227 12448
rect 800 11088 17227 12168
rect 800 10808 17147 11088
rect 800 10408 17227 10808
rect 880 10128 17227 10408
rect 800 8368 17227 10128
rect 800 8088 17147 8368
rect 800 7688 17227 8088
rect 880 7408 17227 7688
rect 800 6328 17227 7408
rect 800 6048 17147 6328
rect 800 5648 17227 6048
rect 880 5368 17227 5648
rect 800 3608 17227 5368
rect 800 3328 17147 3608
rect 800 2928 17227 3328
rect 880 2648 17227 2928
rect 800 1568 17227 2648
rect 800 1395 17147 1568
<< metal4 >>
rect 3566 2128 3886 18000
rect 6188 2128 6508 18000
rect 8810 2128 9130 18000
rect 11432 2128 11752 18000
rect 14054 2128 14374 18000
<< metal5 >>
rect 1104 15115 16836 15435
rect 1104 12485 16836 12805
rect 1104 9856 16836 10176
rect 1104 7227 16836 7547
rect 1104 4597 16836 4917
<< obsm5 >>
rect 1104 13125 16836 14795
rect 1104 10496 16836 12165
rect 1104 7867 16836 9536
<< labels >>
rlabel metal2 s 6918 0 6974 800 6 clockp[0]
port 1 nsew signal output
rlabel metal2 s 6918 19371 6974 20171 6 clockp[1]
port 2 nsew signal output
rlabel metal2 s 10138 19371 10194 20171 6 dco
port 3 nsew signal input
rlabel metal2 s 13818 19371 13874 20171 6 div[0]
port 4 nsew signal input
rlabel metal3 s 17227 3408 18027 3528 6 div[1]
port 5 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 div[2]
port 6 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 div[3]
port 7 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 div[4]
port 8 nsew signal input
rlabel metal2 s 17038 19371 17094 20171 6 enable
port 9 nsew signal input
rlabel metal2 s 8758 19371 8814 20171 6 ext_trim[0]
port 10 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 ext_trim[10]
port 11 nsew signal input
rlabel metal2 s 478 0 534 800 6 ext_trim[11]
port 12 nsew signal input
rlabel metal2 s 3698 19371 3754 20171 6 ext_trim[12]
port 13 nsew signal input
rlabel metal2 s 5538 19371 5594 20171 6 ext_trim[13]
port 14 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 ext_trim[14]
port 15 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 ext_trim[15]
port 16 nsew signal input
rlabel metal3 s 17227 10888 18027 11008 6 ext_trim[16]
port 17 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 ext_trim[17]
port 18 nsew signal input
rlabel metal3 s 17227 1368 18027 1488 6 ext_trim[18]
port 19 nsew signal input
rlabel metal2 s 15198 19371 15254 20171 6 ext_trim[19]
port 20 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 ext_trim[1]
port 21 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 ext_trim[20]
port 22 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 ext_trim[21]
port 23 nsew signal input
rlabel metal3 s 17227 15648 18027 15768 6 ext_trim[22]
port 24 nsew signal input
rlabel metal2 s 2318 19371 2374 20171 6 ext_trim[23]
port 25 nsew signal input
rlabel metal2 s 478 19371 534 20171 6 ext_trim[24]
port 26 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 ext_trim[25]
port 27 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 ext_trim[2]
port 28 nsew signal input
rlabel metal2 s 11978 19371 12034 20171 6 ext_trim[3]
port 29 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 ext_trim[4]
port 30 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 ext_trim[5]
port 31 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 ext_trim[6]
port 32 nsew signal input
rlabel metal3 s 17227 13608 18027 13728 6 ext_trim[7]
port 33 nsew signal input
rlabel metal3 s 17227 6128 18027 6248 6 ext_trim[8]
port 34 nsew signal input
rlabel metal3 s 17227 18368 18027 18488 6 ext_trim[9]
port 35 nsew signal input
rlabel metal3 s 17227 8168 18027 8288 6 osc
port 36 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 resetb
port 37 nsew signal input
rlabel metal4 s 14054 2128 14374 18000 6 VPWR
port 38 nsew power bidirectional
rlabel metal4 s 8810 2128 9130 18000 6 VPWR
port 39 nsew power bidirectional
rlabel metal4 s 3566 2128 3886 18000 6 VPWR
port 40 nsew power bidirectional
rlabel metal5 s 1104 15115 16836 15435 6 VPWR
port 41 nsew power bidirectional
rlabel metal5 s 1104 9856 16836 10176 6 VPWR
port 42 nsew power bidirectional
rlabel metal5 s 1104 4597 16836 4917 6 VPWR
port 43 nsew power bidirectional
rlabel metal4 s 11432 2128 11752 18000 6 VGND
port 44 nsew ground bidirectional
rlabel metal4 s 6188 2128 6508 18000 6 VGND
port 45 nsew ground bidirectional
rlabel metal5 s 1104 12485 16836 12805 6 VGND
port 46 nsew ground bidirectional
rlabel metal5 s 1104 7227 16836 7547 6 VGND
port 47 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 18027 20171
string LEFview TRUE
string GDS_FILE /openLANE_flow/designs/digital_pll/runs/check_run/results/magic/digital_pll.gds
string GDS_END 1267362
string GDS_START 478372
<< end >>

