magic
tech sky130A
magscale 1 2
timestamp 1623890261
<< checkpaint >>
rect -3932 -3932 21178 23322
<< locali >>
rect 5641 16031 5675 16201
rect 4905 12223 4939 12393
rect 3801 8415 3835 8585
rect 7941 5151 7975 5253
<< viali >>
rect 1593 16745 1627 16779
rect 5089 16745 5123 16779
rect 11161 16745 11195 16779
rect 15485 16677 15519 16711
rect 15669 16677 15703 16711
rect 1409 16609 1443 16643
rect 5273 16609 5307 16643
rect 11253 16609 11287 16643
rect 5641 16201 5675 16235
rect 10977 16201 11011 16235
rect 4905 16133 4939 16167
rect 2145 16065 2179 16099
rect 4721 16065 4755 16099
rect 8309 16133 8343 16167
rect 8401 16133 8435 16167
rect 7941 16065 7975 16099
rect 8769 16065 8803 16099
rect 10793 16065 10827 16099
rect 4997 15997 5031 16031
rect 5273 15997 5307 16031
rect 5365 15997 5399 16031
rect 5641 15997 5675 16031
rect 5733 15997 5767 16031
rect 6653 15997 6687 16031
rect 7297 15997 7331 16031
rect 7849 15997 7883 16031
rect 8585 15997 8619 16031
rect 10149 15997 10183 16031
rect 10241 15997 10275 16031
rect 11069 15997 11103 16031
rect 11391 15997 11425 16031
rect 11494 15997 11528 16031
rect 12909 15997 12943 16031
rect 13277 15997 13311 16031
rect 2421 15929 2455 15963
rect 5457 15929 5491 15963
rect 7757 15929 7791 15963
rect 9229 15929 9263 15963
rect 9505 15929 9539 15963
rect 10701 15929 10735 15963
rect 12725 15929 12759 15963
rect 3893 15861 3927 15895
rect 4721 15861 4755 15895
rect 5181 15861 5215 15895
rect 5917 15861 5951 15895
rect 6561 15861 6595 15895
rect 8309 15861 8343 15895
rect 8677 15861 8711 15895
rect 13461 15861 13495 15895
rect 13737 15861 13771 15895
rect 13829 15861 13863 15895
rect 2881 15657 2915 15691
rect 3525 15657 3559 15691
rect 4721 15657 4755 15691
rect 7021 15657 7055 15691
rect 9505 15657 9539 15691
rect 13553 15657 13587 15691
rect 4445 15589 4479 15623
rect 5089 15589 5123 15623
rect 13001 15589 13035 15623
rect 3157 15521 3191 15555
rect 3249 15521 3283 15555
rect 3709 15521 3743 15555
rect 4077 15521 4111 15555
rect 4225 15521 4259 15555
rect 4353 15521 4387 15555
rect 4583 15521 4617 15555
rect 6745 15521 6779 15555
rect 7021 15521 7055 15555
rect 9597 15521 9631 15555
rect 12541 15521 12575 15555
rect 13093 15521 13127 15555
rect 13553 15521 13587 15555
rect 13829 15521 13863 15555
rect 14381 15521 14415 15555
rect 14933 15521 14967 15555
rect 15209 15521 15243 15555
rect 2881 15453 2915 15487
rect 3065 15453 3099 15487
rect 4813 15453 4847 15487
rect 13185 15453 13219 15487
rect 14197 15453 14231 15487
rect 3341 15385 3375 15419
rect 15025 15385 15059 15419
rect 6561 15317 6595 15351
rect 13829 15317 13863 15351
rect 14933 15317 14967 15351
rect 8493 15113 8527 15147
rect 9137 15113 9171 15147
rect 11713 15045 11747 15079
rect 9505 14977 9539 15011
rect 6561 14909 6595 14943
rect 8493 14909 8527 14943
rect 9045 14909 9079 14943
rect 9137 14909 9171 14943
rect 6469 14841 6503 14875
rect 11897 14841 11931 14875
rect 4813 14569 4847 14603
rect 5273 14569 5307 14603
rect 7941 14569 7975 14603
rect 8309 14569 8343 14603
rect 8401 14569 8435 14603
rect 11621 14569 11655 14603
rect 13645 14569 13679 14603
rect 14381 14569 14415 14603
rect 4169 14501 4203 14535
rect 4399 14501 4433 14535
rect 7389 14501 7423 14535
rect 10977 14501 11011 14535
rect 13185 14501 13219 14535
rect 1961 14433 1995 14467
rect 3433 14433 3467 14467
rect 3525 14433 3559 14467
rect 4077 14433 4111 14467
rect 4261 14433 4295 14467
rect 4997 14433 5031 14467
rect 5181 14433 5215 14467
rect 5549 14433 5583 14467
rect 6929 14433 6963 14467
rect 7481 14433 7515 14467
rect 8217 14433 8251 14467
rect 10517 14433 10551 14467
rect 11069 14433 11103 14467
rect 12817 14433 12851 14467
rect 13001 14433 13035 14467
rect 4537 14365 4571 14399
rect 5273 14365 5307 14399
rect 5457 14365 5491 14399
rect 7573 14365 7607 14399
rect 11253 14365 11287 14399
rect 13277 14365 13311 14399
rect 7941 14297 7975 14331
rect 8033 14297 8067 14331
rect 11621 14297 11655 14331
rect 13645 14297 13679 14331
rect 2145 14229 2179 14263
rect 3341 14229 3375 14263
rect 3617 14229 3651 14263
rect 3893 14229 3927 14263
rect 14473 14229 14507 14263
rect 5917 14025 5951 14059
rect 7113 14025 7147 14059
rect 9229 14025 9263 14059
rect 9597 14025 9631 14059
rect 11805 14025 11839 14059
rect 13921 14025 13955 14059
rect 4721 13957 4755 13991
rect 4997 13957 5031 13991
rect 9781 13957 9815 13991
rect 13737 13957 13771 13991
rect 14841 13957 14875 13991
rect 2973 13889 3007 13923
rect 4537 13889 4571 13923
rect 5181 13889 5215 13923
rect 9689 13889 9723 13923
rect 3249 13821 3283 13855
rect 3520 13821 3554 13855
rect 3617 13821 3651 13855
rect 3709 13821 3743 13855
rect 3837 13821 3871 13855
rect 3985 13821 4019 13855
rect 4261 13821 4295 13855
rect 4353 13821 4387 13855
rect 4629 13821 4663 13855
rect 4905 13821 4939 13855
rect 5089 13821 5123 13855
rect 5365 13821 5399 13855
rect 5641 13821 5675 13855
rect 5733 13821 5767 13855
rect 6009 13821 6043 13855
rect 7205 13821 7239 13855
rect 9505 13821 9539 13855
rect 9965 13821 9999 13855
rect 13185 13821 13219 13855
rect 13737 13821 13771 13855
rect 14105 13821 14139 13855
rect 14197 13821 14231 13855
rect 14657 13821 14691 13855
rect 14749 13821 14783 13855
rect 15209 13821 15243 13855
rect 1501 13685 1535 13719
rect 3341 13685 3375 13719
rect 4077 13685 4111 13719
rect 5457 13685 5491 13719
rect 11713 13685 11747 13719
rect 14841 13685 14875 13719
rect 4813 13481 4847 13515
rect 5641 13481 5675 13515
rect 11621 13481 11655 13515
rect 13369 13481 13403 13515
rect 9505 13413 9539 13447
rect 11069 13413 11103 13447
rect 12173 13413 12207 13447
rect 15301 13413 15335 13447
rect 4997 13345 5031 13379
rect 5089 13345 5123 13379
rect 5181 13345 5215 13379
rect 5365 13345 5399 13379
rect 5457 13345 5491 13379
rect 5641 13345 5675 13379
rect 6285 13345 6319 13379
rect 6929 13345 6963 13379
rect 7113 13345 7147 13379
rect 7849 13345 7883 13379
rect 8585 13345 8619 13379
rect 8861 13345 8895 13379
rect 9413 13345 9447 13379
rect 10149 13345 10183 13379
rect 10609 13345 10643 13379
rect 11161 13345 11195 13379
rect 11897 13345 11931 13379
rect 12357 13345 12391 13379
rect 12873 13345 12907 13379
rect 13001 13345 13035 13379
rect 13185 13345 13219 13379
rect 6377 13277 6411 13311
rect 7665 13277 7699 13311
rect 7765 13277 7799 13311
rect 7941 13277 7975 13311
rect 9321 13277 9355 13311
rect 9965 13277 9999 13311
rect 10333 13277 10367 13311
rect 11253 13277 11287 13311
rect 8125 13209 8159 13243
rect 9873 13209 9907 13243
rect 11621 13209 11655 13243
rect 11713 13209 11747 13243
rect 13093 13209 13127 13243
rect 15117 13209 15151 13243
rect 7205 13141 7239 13175
rect 8677 13141 8711 13175
rect 12449 13141 12483 13175
rect 13737 12869 13771 12903
rect 14105 12869 14139 12903
rect 7757 12801 7791 12835
rect 2329 12733 2363 12767
rect 3709 12733 3743 12767
rect 5641 12733 5675 12767
rect 5825 12733 5859 12767
rect 6561 12733 6595 12767
rect 6745 12733 6779 12767
rect 7113 12733 7147 12767
rect 7389 12733 7423 12767
rect 8125 12733 8159 12767
rect 13369 12733 13403 12767
rect 14289 12733 14323 12767
rect 3893 12665 3927 12699
rect 7205 12665 7239 12699
rect 7941 12665 7975 12699
rect 8309 12665 8343 12699
rect 14565 12665 14599 12699
rect 2145 12597 2179 12631
rect 4077 12597 4111 12631
rect 5733 12597 5767 12631
rect 13737 12597 13771 12631
rect 14381 12597 14415 12631
rect 4905 12393 4939 12427
rect 9781 12393 9815 12427
rect 11529 12393 11563 12427
rect 12725 12393 12759 12427
rect 4169 12325 4203 12359
rect 4261 12325 4295 12359
rect 3249 12257 3283 12291
rect 3525 12257 3559 12291
rect 3709 12257 3743 12291
rect 4077 12257 4111 12291
rect 4379 12257 4413 12291
rect 4629 12257 4663 12291
rect 6101 12325 6135 12359
rect 7389 12325 7423 12359
rect 9873 12325 9907 12359
rect 12969 12325 13003 12359
rect 13185 12325 13219 12359
rect 13737 12325 13771 12359
rect 4997 12257 5031 12291
rect 5181 12257 5215 12291
rect 5457 12257 5491 12291
rect 5917 12257 5951 12291
rect 6009 12257 6043 12291
rect 6285 12257 6319 12291
rect 6469 12257 6503 12291
rect 6561 12257 6595 12291
rect 6745 12257 6779 12291
rect 7297 12257 7331 12291
rect 7757 12257 7791 12291
rect 8033 12257 8067 12291
rect 8217 12257 8251 12291
rect 8493 12257 8527 12291
rect 9137 12257 9171 12291
rect 9322 12257 9356 12291
rect 9597 12257 9631 12291
rect 10057 12257 10091 12291
rect 10333 12257 10367 12291
rect 11437 12257 11471 12291
rect 12265 12257 12299 12291
rect 12541 12257 12575 12291
rect 13277 12257 13311 12291
rect 13829 12257 13863 12291
rect 14381 12257 14415 12291
rect 14909 12257 14943 12291
rect 15025 12257 15059 12291
rect 2973 12189 3007 12223
rect 3617 12189 3651 12223
rect 4537 12189 4571 12223
rect 4905 12189 4939 12223
rect 5263 12189 5297 12223
rect 5641 12189 5675 12223
rect 6929 12189 6963 12223
rect 7849 12189 7883 12223
rect 8401 12189 8435 12223
rect 15393 12189 15427 12223
rect 3893 12121 3927 12155
rect 5365 12121 5399 12155
rect 5733 12121 5767 12155
rect 7941 12121 7975 12155
rect 9413 12121 9447 12155
rect 9505 12121 9539 12155
rect 10149 12121 10183 12155
rect 10241 12121 10275 12155
rect 12357 12121 12391 12155
rect 12449 12121 12483 12155
rect 1501 12053 1535 12087
rect 4721 12053 4755 12087
rect 7573 12053 7607 12087
rect 12817 12053 12851 12087
rect 13001 12053 13035 12087
rect 14933 12053 14967 12087
rect 15025 12053 15059 12087
rect 6561 11849 6595 11883
rect 9505 11849 9539 11883
rect 10517 11849 10551 11883
rect 11069 11849 11103 11883
rect 8861 11781 8895 11815
rect 10701 11713 10735 11747
rect 12173 11713 12207 11747
rect 12357 11713 12391 11747
rect 6101 11645 6135 11679
rect 8769 11645 8803 11679
rect 8953 11645 8987 11679
rect 9045 11645 9079 11679
rect 9226 11645 9260 11679
rect 9321 11645 9355 11679
rect 9505 11645 9539 11679
rect 9965 11645 9999 11679
rect 10517 11645 10551 11679
rect 11069 11645 11103 11679
rect 12541 11645 12575 11679
rect 12633 11645 12667 11679
rect 6745 11577 6779 11611
rect 6929 11577 6963 11611
rect 6193 11509 6227 11543
rect 8585 11509 8619 11543
rect 9689 11509 9723 11543
rect 5365 11305 5399 11339
rect 7573 11305 7607 11339
rect 10977 11305 11011 11339
rect 15301 11237 15335 11271
rect 4261 11169 4295 11203
rect 4445 11169 4479 11203
rect 6837 11169 6871 11203
rect 7021 11169 7055 11203
rect 7205 11169 7239 11203
rect 7297 11169 7331 11203
rect 7665 11169 7699 11203
rect 9321 11169 9355 11203
rect 9597 11169 9631 11203
rect 9781 11169 9815 11203
rect 10885 11169 10919 11203
rect 1409 11101 1443 11135
rect 5457 11101 5491 11135
rect 5549 11101 5583 11135
rect 7757 11101 7791 11135
rect 9505 11101 9539 11135
rect 7113 11033 7147 11067
rect 9137 11033 9171 11067
rect 9413 11033 9447 11067
rect 15117 11033 15151 11067
rect 1672 10965 1706 10999
rect 3157 10965 3191 10999
rect 4261 10965 4295 10999
rect 4629 10965 4663 10999
rect 4997 10965 5031 10999
rect 2145 10761 2179 10795
rect 2789 10761 2823 10795
rect 2881 10761 2915 10795
rect 4997 10761 5031 10795
rect 8125 10761 8159 10795
rect 8677 10761 8711 10795
rect 9505 10761 9539 10795
rect 3065 10693 3099 10727
rect 8217 10693 8251 10727
rect 9137 10693 9171 10727
rect 10977 10693 11011 10727
rect 11069 10693 11103 10727
rect 12081 10693 12115 10727
rect 14289 10693 14323 10727
rect 14381 10693 14415 10727
rect 2743 10625 2777 10659
rect 4537 10625 4571 10659
rect 9008 10625 9042 10659
rect 9229 10625 9263 10659
rect 10609 10625 10643 10659
rect 11989 10625 12023 10659
rect 13921 10625 13955 10659
rect 1961 10557 1995 10591
rect 2973 10557 3007 10591
rect 3249 10557 3283 10591
rect 3341 10557 3375 10591
rect 3709 10557 3743 10591
rect 3939 10557 3973 10591
rect 4077 10557 4111 10591
rect 4353 10557 4387 10591
rect 4445 10557 4479 10591
rect 4721 10557 4755 10591
rect 4813 10557 4847 10591
rect 5089 10557 5123 10591
rect 5273 10557 5307 10591
rect 5365 10557 5399 10591
rect 5457 10557 5491 10591
rect 7941 10557 7975 10591
rect 8309 10557 8343 10591
rect 8401 10557 8435 10591
rect 9965 10557 9999 10591
rect 10517 10557 10551 10591
rect 11253 10557 11287 10591
rect 11897 10557 11931 10591
rect 12173 10557 12207 10591
rect 13277 10557 13311 10591
rect 13829 10557 13863 10591
rect 14565 10557 14599 10591
rect 2605 10489 2639 10523
rect 3617 10489 3651 10523
rect 4169 10489 4203 10523
rect 8861 10489 8895 10523
rect 10425 10489 10459 10523
rect 13737 10489 13771 10523
rect 3801 10421 3835 10455
rect 5733 10421 5767 10455
rect 10977 10421 11011 10455
rect 11713 10421 11747 10455
rect 14289 10421 14323 10455
rect 14657 10421 14691 10455
rect 14749 10421 14783 10455
rect 3617 10217 3651 10251
rect 6193 10217 6227 10251
rect 5365 10149 5399 10183
rect 13461 10149 13495 10183
rect 13645 10149 13679 10183
rect 3709 10081 3743 10115
rect 4445 10081 4479 10115
rect 4721 10081 4755 10115
rect 4813 10081 4847 10115
rect 5825 10081 5859 10115
rect 6252 10081 6286 10115
rect 6561 10081 6595 10115
rect 7573 10081 7607 10115
rect 7665 10081 7699 10115
rect 10241 10081 10275 10115
rect 10517 10081 10551 10115
rect 12081 10081 12115 10115
rect 12541 10081 12575 10115
rect 12633 10081 12667 10115
rect 12817 10081 12851 10115
rect 13001 10081 13035 10115
rect 13093 10081 13127 10115
rect 13369 10081 13403 10115
rect 14381 10081 14415 10115
rect 14933 10081 14967 10115
rect 15025 10081 15059 10115
rect 15761 10081 15795 10115
rect 4261 10013 4295 10047
rect 5733 10013 5767 10047
rect 7481 10013 7515 10047
rect 7757 10013 7791 10047
rect 10333 10013 10367 10047
rect 12173 10013 12207 10047
rect 15393 10013 15427 10047
rect 10425 9945 10459 9979
rect 12265 9945 12299 9979
rect 6377 9877 6411 9911
rect 6745 9877 6779 9911
rect 7297 9877 7331 9911
rect 10057 9877 10091 9911
rect 11805 9877 11839 9911
rect 12357 9877 12391 9911
rect 12909 9877 12943 9911
rect 13829 9877 13863 9911
rect 14933 9877 14967 9911
rect 15025 9877 15059 9911
rect 15577 9877 15611 9911
rect 2973 9673 3007 9707
rect 8217 9673 8251 9707
rect 11069 9673 11103 9707
rect 3249 9605 3283 9639
rect 6745 9537 6779 9571
rect 1409 9469 1443 9503
rect 2053 9469 2087 9503
rect 2697 9469 2731 9503
rect 2789 9469 2823 9503
rect 3065 9469 3099 9503
rect 3341 9469 3375 9503
rect 6469 9469 6503 9503
rect 8769 9469 8803 9503
rect 9597 9469 9631 9503
rect 15301 9469 15335 9503
rect 8401 9401 8435 9435
rect 8585 9401 8619 9435
rect 10977 9401 11011 9435
rect 15117 9401 15151 9435
rect 1593 9333 1627 9367
rect 2237 9333 2271 9367
rect 2513 9333 2547 9367
rect 9781 9333 9815 9367
rect 9781 9129 9815 9163
rect 10609 9129 10643 9163
rect 1685 9061 1719 9095
rect 6193 9061 6227 9095
rect 9597 9061 9631 9095
rect 10701 9061 10735 9095
rect 3893 8993 3927 9027
rect 4077 8993 4111 9027
rect 4537 8993 4571 9027
rect 4721 8993 4755 9027
rect 5181 8993 5215 9027
rect 5917 8993 5951 9027
rect 6377 8993 6411 9027
rect 9137 8993 9171 9027
rect 9689 8993 9723 9027
rect 10241 8993 10275 9027
rect 12541 8993 12575 9027
rect 13093 8993 13127 9027
rect 13277 8993 13311 9027
rect 13553 8993 13587 9027
rect 1409 8925 1443 8959
rect 10149 8925 10183 8959
rect 13001 8925 13035 8959
rect 9781 8857 9815 8891
rect 10609 8857 10643 8891
rect 10793 8857 10827 8891
rect 3157 8789 3191 8823
rect 3893 8789 3927 8823
rect 4261 8789 4295 8823
rect 4813 8789 4847 8823
rect 5273 8789 5307 8823
rect 5825 8789 5859 8823
rect 6009 8789 6043 8823
rect 13277 8789 13311 8823
rect 13737 8789 13771 8823
rect 3801 8585 3835 8619
rect 4721 8585 4755 8619
rect 10517 8585 10551 8619
rect 2421 8517 2455 8551
rect 4629 8517 4663 8551
rect 5641 8517 5675 8551
rect 13093 8517 13127 8551
rect 13553 8517 13587 8551
rect 15209 8517 15243 8551
rect 15301 8517 15335 8551
rect 4169 8449 4203 8483
rect 5089 8449 5123 8483
rect 7389 8449 7423 8483
rect 14013 8449 14047 8483
rect 14841 8449 14875 8483
rect 2237 8381 2271 8415
rect 2421 8381 2455 8415
rect 3801 8381 3835 8415
rect 3893 8381 3927 8415
rect 4077 8381 4111 8415
rect 4261 8381 4295 8415
rect 4445 8381 4479 8415
rect 4905 8381 4939 8415
rect 5181 8381 5215 8415
rect 5273 8381 5307 8415
rect 5457 8381 5491 8415
rect 5917 8381 5951 8415
rect 6009 8381 6043 8415
rect 6101 8381 6135 8415
rect 6285 8381 6319 8415
rect 6561 8381 6595 8415
rect 6653 8381 6687 8415
rect 6929 8381 6963 8415
rect 7113 8381 7147 8415
rect 7757 8381 7791 8415
rect 9965 8381 9999 8415
rect 10517 8381 10551 8415
rect 11805 8381 11839 8415
rect 13277 8381 13311 8415
rect 14197 8381 14231 8415
rect 14749 8381 14783 8415
rect 15485 8381 15519 8415
rect 6837 8313 6871 8347
rect 8401 8313 8435 8347
rect 13461 8313 13495 8347
rect 14657 8313 14691 8347
rect 7757 8245 7791 8279
rect 8217 8245 8251 8279
rect 15209 8245 15243 8279
rect 8585 8041 8619 8075
rect 8677 8041 8711 8075
rect 9689 8041 9723 8075
rect 13461 8041 13495 8075
rect 14749 8041 14783 8075
rect 2973 7973 3007 8007
rect 4261 7973 4295 8007
rect 7757 7973 7791 8007
rect 9597 7973 9631 8007
rect 1869 7905 1903 7939
rect 2329 7905 2363 7939
rect 2697 7905 2731 7939
rect 3157 7905 3191 7939
rect 3341 7905 3375 7939
rect 4353 7905 4387 7939
rect 4905 7905 4939 7939
rect 5089 7905 5123 7939
rect 5641 7905 5675 7939
rect 5825 7905 5859 7939
rect 7297 7905 7331 7939
rect 7849 7905 7883 7939
rect 8585 7905 8619 7939
rect 8861 7905 8895 7939
rect 11805 7905 11839 7939
rect 13277 7905 13311 7939
rect 13645 7905 13679 7939
rect 14657 7905 14691 7939
rect 2237 7837 2271 7871
rect 2605 7837 2639 7871
rect 8217 7837 8251 7871
rect 13093 7837 13127 7871
rect 2513 7769 2547 7803
rect 14473 7769 14507 7803
rect 14841 7701 14875 7735
rect 2697 7497 2731 7531
rect 5181 7497 5215 7531
rect 8769 7497 8803 7531
rect 3341 7429 3375 7463
rect 10793 7429 10827 7463
rect 11069 7429 11103 7463
rect 15025 7429 15059 7463
rect 2053 7361 2087 7395
rect 2421 7361 2455 7395
rect 3525 7361 3559 7395
rect 10425 7361 10459 7395
rect 14657 7361 14691 7395
rect 2513 7293 2547 7327
rect 2789 7293 2823 7327
rect 3157 7293 3191 7327
rect 3433 7293 3467 7327
rect 5089 7293 5123 7327
rect 8217 7293 8251 7327
rect 8769 7293 8803 7327
rect 11253 7293 11287 7327
rect 14013 7293 14047 7327
rect 14565 7293 14599 7327
rect 2973 7225 3007 7259
rect 3065 7225 3099 7259
rect 14473 7225 14507 7259
rect 10793 7157 10827 7191
rect 11345 7157 11379 7191
rect 11437 7157 11471 7191
rect 15025 7157 15059 7191
rect 3893 6953 3927 6987
rect 4077 6953 4111 6987
rect 6561 6953 6595 6987
rect 5181 6885 5215 6919
rect 5825 6885 5859 6919
rect 9597 6885 9631 6919
rect 10701 6885 10735 6919
rect 4074 6817 4108 6851
rect 4629 6817 4663 6851
rect 4721 6817 4755 6851
rect 4905 6817 4939 6851
rect 5365 6817 5399 6851
rect 5457 6817 5491 6851
rect 5917 6817 5951 6851
rect 6193 6817 6227 6851
rect 6285 6817 6319 6851
rect 6837 6817 6871 6851
rect 7205 6817 7239 6851
rect 7297 6817 7331 6851
rect 9781 6817 9815 6851
rect 10241 6817 10275 6851
rect 10793 6817 10827 6851
rect 11253 6817 11287 6851
rect 11989 6817 12023 6851
rect 13185 6817 13219 6851
rect 4537 6749 4571 6783
rect 5089 6749 5123 6783
rect 6745 6749 6779 6783
rect 7113 6749 7147 6783
rect 11345 6749 11379 6783
rect 12265 6749 12299 6783
rect 12909 6749 12943 6783
rect 5181 6681 5215 6715
rect 6469 6681 6503 6715
rect 4445 6613 4479 6647
rect 7389 6613 7423 6647
rect 4077 6409 4111 6443
rect 4905 6409 4939 6443
rect 7021 6409 7055 6443
rect 7573 6409 7607 6443
rect 7757 6409 7791 6443
rect 5365 6273 5399 6307
rect 6101 6273 6135 6307
rect 13185 6273 13219 6307
rect 2145 6205 2179 6239
rect 2513 6205 2547 6239
rect 2697 6205 2731 6239
rect 2881 6205 2915 6239
rect 3893 6205 3927 6239
rect 4077 6205 4111 6239
rect 5089 6205 5123 6239
rect 5273 6205 5307 6239
rect 5457 6205 5491 6239
rect 5641 6205 5675 6239
rect 5733 6205 5767 6239
rect 5917 6205 5951 6239
rect 6009 6205 6043 6239
rect 7202 6205 7236 6239
rect 7665 6205 7699 6239
rect 8033 6205 8067 6239
rect 8125 6205 8159 6239
rect 8309 6205 8343 6239
rect 9597 6205 9631 6239
rect 11713 6205 11747 6239
rect 12081 6205 12115 6239
rect 12173 6205 12207 6239
rect 12909 6205 12943 6239
rect 13645 6205 13679 6239
rect 2789 6137 2823 6171
rect 5825 6137 5859 6171
rect 7757 6137 7791 6171
rect 8217 6137 8251 6171
rect 11897 6137 11931 6171
rect 13093 6137 13127 6171
rect 1961 6069 1995 6103
rect 3065 6069 3099 6103
rect 7205 6069 7239 6103
rect 7941 6069 7975 6103
rect 9781 6069 9815 6103
rect 13829 6069 13863 6103
rect 1409 5865 1443 5899
rect 6837 5865 6871 5899
rect 9137 5865 9171 5899
rect 2881 5797 2915 5831
rect 4169 5797 4203 5831
rect 6469 5797 6503 5831
rect 8585 5797 8619 5831
rect 3893 5729 3927 5763
rect 4077 5729 4111 5763
rect 4261 5729 4295 5763
rect 6285 5729 6319 5763
rect 6561 5729 6595 5763
rect 6653 5729 6687 5763
rect 8309 5729 8343 5763
rect 8493 5729 8527 5763
rect 8677 5729 8711 5763
rect 11253 5729 11287 5763
rect 12357 5729 12391 5763
rect 14473 5729 14507 5763
rect 3157 5661 3191 5695
rect 10609 5661 10643 5695
rect 10885 5661 10919 5695
rect 8861 5593 8895 5627
rect 12173 5593 12207 5627
rect 4445 5525 4479 5559
rect 11253 5525 11287 5559
rect 14473 5525 14507 5559
rect 3249 5321 3283 5355
rect 5365 5321 5399 5355
rect 6469 5321 6503 5355
rect 7941 5253 7975 5287
rect 10977 5253 11011 5287
rect 4721 5185 4755 5219
rect 4997 5185 5031 5219
rect 7021 5185 7055 5219
rect 12357 5185 12391 5219
rect 13829 5185 13863 5219
rect 5273 5117 5307 5151
rect 5825 5117 5859 5151
rect 6650 5117 6684 5151
rect 7113 5117 7147 5151
rect 7941 5117 7975 5151
rect 8217 5117 8251 5151
rect 9045 5117 9079 5151
rect 9413 5117 9447 5151
rect 10517 5117 10551 5151
rect 11161 5117 11195 5151
rect 12173 5117 12207 5151
rect 12449 5117 12483 5151
rect 13185 5117 13219 5151
rect 9229 5049 9263 5083
rect 9321 5049 9355 5083
rect 11253 5049 11287 5083
rect 11529 5049 11563 5083
rect 14105 5049 14139 5083
rect 5549 4981 5583 5015
rect 5733 4981 5767 5015
rect 6653 4981 6687 5015
rect 8033 4981 8067 5015
rect 9597 4981 9631 5015
rect 10333 4981 10367 5015
rect 11345 4981 11379 5015
rect 13001 4981 13035 5015
rect 15577 4981 15611 5015
rect 2605 4777 2639 4811
rect 2881 4777 2915 4811
rect 4169 4777 4203 4811
rect 6101 4777 6135 4811
rect 9413 4777 9447 4811
rect 11989 4777 12023 4811
rect 14197 4777 14231 4811
rect 2421 4709 2455 4743
rect 10885 4709 10919 4743
rect 11529 4709 11563 4743
rect 2053 4641 2087 4675
rect 2697 4641 2731 4675
rect 2973 4641 3007 4675
rect 4353 4641 4387 4675
rect 5457 4641 5491 4675
rect 6009 4641 6043 4675
rect 6929 4641 6963 4675
rect 11345 4641 11379 4675
rect 11621 4641 11655 4675
rect 11713 4641 11747 4675
rect 13737 4641 13771 4675
rect 14013 4641 14047 4675
rect 14841 4641 14875 4675
rect 15025 4641 15059 4675
rect 15577 4641 15611 4675
rect 5365 4573 5399 4607
rect 7205 4573 7239 4607
rect 8953 4573 8987 4607
rect 11161 4573 11195 4607
rect 13461 4573 13495 4607
rect 15669 4573 15703 4607
rect 11897 4505 11931 4539
rect 2237 4437 2271 4471
rect 2421 4437 2455 4471
rect 14565 4437 14599 4471
rect 1672 4233 1706 4267
rect 3157 4233 3191 4267
rect 15761 4233 15795 4267
rect 1409 4097 1443 4131
rect 5641 4097 5675 4131
rect 14013 4097 14047 4131
rect 5549 4029 5583 4063
rect 6101 4029 6135 4063
rect 7297 4029 7331 4063
rect 11713 4029 11747 4063
rect 11989 4029 12023 4063
rect 12081 4029 12115 4063
rect 11897 3961 11931 3995
rect 14289 3961 14323 3995
rect 7205 3893 7239 3927
rect 12265 3893 12299 3927
rect 4261 3689 4295 3723
rect 8585 3689 8619 3723
rect 12081 3689 12115 3723
rect 3985 3621 4019 3655
rect 9413 3621 9447 3655
rect 13553 3621 13587 3655
rect 4169 3553 4203 3587
rect 4353 3553 4387 3587
rect 6285 3553 6319 3587
rect 6469 3553 6503 3587
rect 6837 3553 6871 3587
rect 7481 3553 7515 3587
rect 8677 3553 8711 3587
rect 9137 3553 9171 3587
rect 9321 3553 9355 3587
rect 9505 3553 9539 3587
rect 10057 3553 10091 3587
rect 13829 3553 13863 3587
rect 6561 3485 6595 3519
rect 6653 3485 6687 3519
rect 7293 3485 7327 3519
rect 7389 3485 7423 3519
rect 7573 3485 7607 3519
rect 10241 3485 10275 3519
rect 10517 3485 10551 3519
rect 11989 3485 12023 3519
rect 4537 3349 4571 3383
rect 7021 3349 7055 3383
rect 7113 3349 7147 3383
rect 9689 3349 9723 3383
rect 9873 3349 9907 3383
rect 1593 3145 1627 3179
rect 6193 3145 6227 3179
rect 9137 3145 9171 3179
rect 9321 3145 9355 3179
rect 11161 3145 11195 3179
rect 14565 3145 14599 3179
rect 14933 3145 14967 3179
rect 3893 3077 3927 3111
rect 5825 3077 5859 3111
rect 6101 3077 6135 3111
rect 6653 3077 6687 3111
rect 3157 3009 3191 3043
rect 3617 3009 3651 3043
rect 4813 3009 4847 3043
rect 6285 3009 6319 3043
rect 7389 3009 7423 3043
rect 10793 3009 10827 3043
rect 11069 3009 11103 3043
rect 12817 3009 12851 3043
rect 13093 3009 13127 3043
rect 1409 2941 1443 2975
rect 2237 2941 2271 2975
rect 2881 2941 2915 2975
rect 3065 2941 3099 2975
rect 3249 2941 3283 2975
rect 3433 2941 3467 2975
rect 3525 2941 3559 2975
rect 3709 2941 3743 2975
rect 4077 2941 4111 2975
rect 4445 2941 4479 2975
rect 4537 2941 4571 2975
rect 4905 2941 4939 2975
rect 5181 2941 5215 2975
rect 5733 2941 5767 2975
rect 6009 2941 6043 2975
rect 6561 2941 6595 2975
rect 6837 2941 6871 2975
rect 11345 2941 11379 2975
rect 14749 2941 14783 2975
rect 2697 2873 2731 2907
rect 4169 2873 4203 2907
rect 4261 2873 4295 2907
rect 7665 2873 7699 2907
rect 11529 2873 11563 2907
rect 2421 2805 2455 2839
rect 4997 2805 5031 2839
rect 7021 2805 7055 2839
rect 3157 2601 3191 2635
rect 5641 2601 5675 2635
rect 5917 2601 5951 2635
rect 6745 2601 6779 2635
rect 7481 2601 7515 2635
rect 8585 2601 8619 2635
rect 11253 2601 11287 2635
rect 12173 2601 12207 2635
rect 13921 2601 13955 2635
rect 15577 2601 15611 2635
rect 1685 2533 1719 2567
rect 4169 2533 4203 2567
rect 6193 2533 6227 2567
rect 7113 2533 7147 2567
rect 7297 2533 7331 2567
rect 1409 2465 1443 2499
rect 5733 2465 5767 2499
rect 6837 2465 6871 2499
rect 8401 2465 8435 2499
rect 11069 2465 11103 2499
rect 11989 2465 12023 2499
rect 13737 2465 13771 2499
rect 15761 2465 15795 2499
rect 3893 2397 3927 2431
rect 6009 2329 6043 2363
<< metal1 >>
rect 1104 16890 16100 16912
rect 1104 16838 5980 16890
rect 6032 16838 6044 16890
rect 6096 16838 6108 16890
rect 6160 16838 6172 16890
rect 6224 16838 10979 16890
rect 11031 16838 11043 16890
rect 11095 16838 11107 16890
rect 11159 16838 11171 16890
rect 11223 16838 16100 16890
rect 1104 16816 16100 16838
rect 1581 16779 1639 16785
rect 1581 16745 1593 16779
rect 1627 16776 1639 16779
rect 2314 16776 2320 16788
rect 1627 16748 2320 16776
rect 1627 16745 1639 16748
rect 1581 16739 1639 16745
rect 2314 16736 2320 16748
rect 2372 16736 2378 16788
rect 4522 16736 4528 16788
rect 4580 16776 4586 16788
rect 5077 16779 5135 16785
rect 5077 16776 5089 16779
rect 4580 16748 5089 16776
rect 4580 16736 4586 16748
rect 5077 16745 5089 16748
rect 5123 16745 5135 16779
rect 5077 16739 5135 16745
rect 11149 16779 11207 16785
rect 11149 16745 11161 16779
rect 11195 16776 11207 16779
rect 11330 16776 11336 16788
rect 11195 16748 11336 16776
rect 11195 16745 11207 16748
rect 11149 16739 11207 16745
rect 11330 16736 11336 16748
rect 11388 16736 11394 16788
rect 6730 16668 6736 16720
rect 6788 16708 6794 16720
rect 15473 16711 15531 16717
rect 15473 16708 15485 16711
rect 6788 16680 15485 16708
rect 6788 16668 6794 16680
rect 15473 16677 15485 16680
rect 15519 16677 15531 16711
rect 15473 16671 15531 16677
rect 15657 16711 15715 16717
rect 15657 16677 15669 16711
rect 15703 16708 15715 16711
rect 16574 16708 16580 16720
rect 15703 16680 16580 16708
rect 15703 16677 15715 16680
rect 15657 16671 15715 16677
rect 16574 16668 16580 16680
rect 16632 16668 16638 16720
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 5074 16600 5080 16652
rect 5132 16640 5138 16652
rect 5261 16643 5319 16649
rect 5261 16640 5273 16643
rect 5132 16612 5273 16640
rect 5132 16600 5138 16612
rect 5261 16609 5273 16612
rect 5307 16609 5319 16643
rect 11238 16640 11244 16652
rect 11199 16612 11244 16640
rect 5261 16603 5319 16609
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 1104 16346 16100 16368
rect 1104 16294 3481 16346
rect 3533 16294 3545 16346
rect 3597 16294 3609 16346
rect 3661 16294 3673 16346
rect 3725 16294 8480 16346
rect 8532 16294 8544 16346
rect 8596 16294 8608 16346
rect 8660 16294 8672 16346
rect 8724 16294 13478 16346
rect 13530 16294 13542 16346
rect 13594 16294 13606 16346
rect 13658 16294 13670 16346
rect 13722 16294 16100 16346
rect 1104 16272 16100 16294
rect 3786 16192 3792 16244
rect 3844 16232 3850 16244
rect 5629 16235 5687 16241
rect 5629 16232 5641 16235
rect 3844 16204 5641 16232
rect 3844 16192 3850 16204
rect 5629 16201 5641 16204
rect 5675 16201 5687 16235
rect 5629 16195 5687 16201
rect 10965 16235 11023 16241
rect 10965 16201 10977 16235
rect 11011 16232 11023 16235
rect 11238 16232 11244 16244
rect 11011 16204 11244 16232
rect 11011 16201 11023 16204
rect 10965 16195 11023 16201
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 3418 16124 3424 16176
rect 3476 16164 3482 16176
rect 4430 16164 4436 16176
rect 3476 16136 4436 16164
rect 3476 16124 3482 16136
rect 4430 16124 4436 16136
rect 4488 16164 4494 16176
rect 4893 16167 4951 16173
rect 4893 16164 4905 16167
rect 4488 16136 4905 16164
rect 4488 16124 4494 16136
rect 4893 16133 4905 16136
rect 4939 16133 4951 16167
rect 4893 16127 4951 16133
rect 8297 16167 8355 16173
rect 8297 16133 8309 16167
rect 8343 16164 8355 16167
rect 8389 16167 8447 16173
rect 8389 16164 8401 16167
rect 8343 16136 8401 16164
rect 8343 16133 8355 16136
rect 8297 16127 8355 16133
rect 8389 16133 8401 16136
rect 8435 16133 8447 16167
rect 8389 16127 8447 16133
rect 2133 16099 2191 16105
rect 2133 16065 2145 16099
rect 2179 16096 2191 16099
rect 3142 16096 3148 16108
rect 2179 16068 3148 16096
rect 2179 16065 2191 16068
rect 2133 16059 2191 16065
rect 3142 16056 3148 16068
rect 3200 16056 3206 16108
rect 4706 16096 4712 16108
rect 4667 16068 4712 16096
rect 4706 16056 4712 16068
rect 4764 16056 4770 16108
rect 6546 16096 6552 16108
rect 5000 16068 6552 16096
rect 3510 15988 3516 16040
rect 3568 15988 3574 16040
rect 5000 16037 5028 16068
rect 6546 16056 6552 16068
rect 6604 16056 6610 16108
rect 7929 16099 7987 16105
rect 7929 16096 7941 16099
rect 7300 16068 7941 16096
rect 4985 16031 5043 16037
rect 4985 15997 4997 16031
rect 5031 15997 5043 16031
rect 4985 15991 5043 15997
rect 5074 15988 5080 16040
rect 5132 16028 5138 16040
rect 5261 16031 5319 16037
rect 5261 16028 5273 16031
rect 5132 16000 5273 16028
rect 5132 15988 5138 16000
rect 5261 15997 5273 16000
rect 5307 15997 5319 16031
rect 5261 15991 5319 15997
rect 5350 15988 5356 16040
rect 5408 16028 5414 16040
rect 5629 16031 5687 16037
rect 5408 16000 5453 16028
rect 5408 15988 5414 16000
rect 5629 15997 5641 16031
rect 5675 16028 5687 16031
rect 5721 16031 5779 16037
rect 5721 16028 5733 16031
rect 5675 16000 5733 16028
rect 5675 15997 5687 16000
rect 5629 15991 5687 15997
rect 5721 15997 5733 16000
rect 5767 15997 5779 16031
rect 6638 16028 6644 16040
rect 6599 16000 6644 16028
rect 5721 15991 5779 15997
rect 6638 15988 6644 16000
rect 6696 15988 6702 16040
rect 7006 15988 7012 16040
rect 7064 16028 7070 16040
rect 7300 16037 7328 16068
rect 7929 16065 7941 16068
rect 7975 16065 7987 16099
rect 7929 16059 7987 16065
rect 8757 16099 8815 16105
rect 8757 16065 8769 16099
rect 8803 16096 8815 16099
rect 10781 16099 10839 16105
rect 10781 16096 10793 16099
rect 8803 16068 10793 16096
rect 8803 16065 8815 16068
rect 8757 16059 8815 16065
rect 10781 16065 10793 16068
rect 10827 16065 10839 16099
rect 10781 16059 10839 16065
rect 7285 16031 7343 16037
rect 7285 16028 7297 16031
rect 7064 16000 7297 16028
rect 7064 15988 7070 16000
rect 7285 15997 7297 16000
rect 7331 15997 7343 16031
rect 7285 15991 7343 15997
rect 7837 16031 7895 16037
rect 7837 15997 7849 16031
rect 7883 16028 7895 16031
rect 8573 16031 8631 16037
rect 8573 16028 8585 16031
rect 7883 16000 8585 16028
rect 7883 15997 7895 16000
rect 7837 15991 7895 15997
rect 8573 15997 8585 16000
rect 8619 15997 8631 16031
rect 8573 15991 8631 15997
rect 2406 15960 2412 15972
rect 2367 15932 2412 15960
rect 2406 15920 2412 15932
rect 2464 15920 2470 15972
rect 4246 15920 4252 15972
rect 4304 15960 4310 15972
rect 5445 15963 5503 15969
rect 5445 15960 5457 15963
rect 4304 15932 5457 15960
rect 4304 15920 4310 15932
rect 5445 15929 5457 15932
rect 5491 15929 5503 15963
rect 5445 15923 5503 15929
rect 7745 15963 7803 15969
rect 7745 15929 7757 15963
rect 7791 15929 7803 15963
rect 8588 15960 8616 15991
rect 9858 15988 9864 16040
rect 9916 16028 9922 16040
rect 10137 16031 10195 16037
rect 10137 16028 10149 16031
rect 9916 16000 10149 16028
rect 9916 15988 9922 16000
rect 10137 15997 10149 16000
rect 10183 16028 10195 16031
rect 10229 16031 10287 16037
rect 10229 16028 10241 16031
rect 10183 16000 10241 16028
rect 10183 15997 10195 16000
rect 10137 15991 10195 15997
rect 10229 15997 10241 16000
rect 10275 15997 10287 16031
rect 10229 15991 10287 15997
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 16028 11115 16031
rect 11379 16031 11437 16037
rect 11379 16028 11391 16031
rect 11103 16000 11391 16028
rect 11103 15997 11115 16000
rect 11057 15991 11115 15997
rect 11379 15997 11391 16000
rect 11425 15997 11437 16031
rect 11379 15991 11437 15997
rect 11482 16031 11540 16037
rect 11482 15997 11494 16031
rect 11528 16028 11540 16031
rect 12897 16031 12955 16037
rect 11528 15997 11560 16028
rect 11482 15991 11560 15997
rect 12897 15997 12909 16031
rect 12943 16028 12955 16031
rect 13262 16028 13268 16040
rect 12943 16000 13268 16028
rect 12943 15997 12955 16000
rect 12897 15991 12955 15997
rect 9214 15960 9220 15972
rect 8588 15932 9220 15960
rect 7745 15923 7803 15929
rect 3881 15895 3939 15901
rect 3881 15861 3893 15895
rect 3927 15892 3939 15895
rect 4614 15892 4620 15904
rect 3927 15864 4620 15892
rect 3927 15861 3939 15864
rect 3881 15855 3939 15861
rect 4614 15852 4620 15864
rect 4672 15852 4678 15904
rect 4709 15895 4767 15901
rect 4709 15861 4721 15895
rect 4755 15892 4767 15895
rect 5074 15892 5080 15904
rect 4755 15864 5080 15892
rect 4755 15861 4767 15864
rect 4709 15855 4767 15861
rect 5074 15852 5080 15864
rect 5132 15852 5138 15904
rect 5166 15852 5172 15904
rect 5224 15892 5230 15904
rect 5224 15864 5269 15892
rect 5224 15852 5230 15864
rect 5810 15852 5816 15904
rect 5868 15892 5874 15904
rect 5905 15895 5963 15901
rect 5905 15892 5917 15895
rect 5868 15864 5917 15892
rect 5868 15852 5874 15864
rect 5905 15861 5917 15864
rect 5951 15861 5963 15895
rect 6546 15892 6552 15904
rect 6507 15864 6552 15892
rect 5905 15855 5963 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 7760 15892 7788 15923
rect 9214 15920 9220 15932
rect 9272 15920 9278 15972
rect 9493 15963 9551 15969
rect 9493 15929 9505 15963
rect 9539 15960 9551 15963
rect 10689 15963 10747 15969
rect 10689 15960 10701 15963
rect 9539 15932 10701 15960
rect 9539 15929 9551 15932
rect 9493 15923 9551 15929
rect 10689 15929 10701 15932
rect 10735 15960 10747 15963
rect 11532 15960 11560 15991
rect 13262 15988 13268 16000
rect 13320 15988 13326 16040
rect 12713 15963 12771 15969
rect 12713 15960 12725 15963
rect 10735 15932 12725 15960
rect 10735 15929 10747 15932
rect 10689 15923 10747 15929
rect 12713 15929 12725 15932
rect 12759 15929 12771 15963
rect 12713 15923 12771 15929
rect 8297 15895 8355 15901
rect 8297 15892 8309 15895
rect 7760 15864 8309 15892
rect 8297 15861 8309 15864
rect 8343 15892 8355 15895
rect 8665 15895 8723 15901
rect 8665 15892 8677 15895
rect 8343 15864 8677 15892
rect 8343 15861 8355 15864
rect 8297 15855 8355 15861
rect 8665 15861 8677 15864
rect 8711 15861 8723 15895
rect 8665 15855 8723 15861
rect 13449 15895 13507 15901
rect 13449 15861 13461 15895
rect 13495 15892 13507 15895
rect 13538 15892 13544 15904
rect 13495 15864 13544 15892
rect 13495 15861 13507 15864
rect 13449 15855 13507 15861
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 13722 15892 13728 15904
rect 13683 15864 13728 15892
rect 13722 15852 13728 15864
rect 13780 15852 13786 15904
rect 13814 15852 13820 15904
rect 13872 15892 13878 15904
rect 13872 15864 13917 15892
rect 13872 15852 13878 15864
rect 1104 15802 16100 15824
rect 1104 15750 5980 15802
rect 6032 15750 6044 15802
rect 6096 15750 6108 15802
rect 6160 15750 6172 15802
rect 6224 15750 10979 15802
rect 11031 15750 11043 15802
rect 11095 15750 11107 15802
rect 11159 15750 11171 15802
rect 11223 15750 16100 15802
rect 1104 15728 16100 15750
rect 2406 15648 2412 15700
rect 2464 15688 2470 15700
rect 2869 15691 2927 15697
rect 2869 15688 2881 15691
rect 2464 15660 2881 15688
rect 2464 15648 2470 15660
rect 2869 15657 2881 15660
rect 2915 15657 2927 15691
rect 3510 15688 3516 15700
rect 3471 15660 3516 15688
rect 2869 15651 2927 15657
rect 3510 15648 3516 15660
rect 3568 15648 3574 15700
rect 4154 15648 4160 15700
rect 4212 15648 4218 15700
rect 4706 15688 4712 15700
rect 4667 15660 4712 15688
rect 4706 15648 4712 15660
rect 4764 15648 4770 15700
rect 5166 15688 5172 15700
rect 4816 15660 5172 15688
rect 4172 15620 4200 15648
rect 3160 15592 4200 15620
rect 4433 15623 4491 15629
rect 3160 15561 3188 15592
rect 4433 15589 4445 15623
rect 4479 15620 4491 15623
rect 4816 15620 4844 15660
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 7006 15688 7012 15700
rect 6967 15660 7012 15688
rect 7006 15648 7012 15660
rect 7064 15648 7070 15700
rect 9214 15648 9220 15700
rect 9272 15688 9278 15700
rect 9493 15691 9551 15697
rect 9493 15688 9505 15691
rect 9272 15660 9505 15688
rect 9272 15648 9278 15660
rect 9493 15657 9505 15660
rect 9539 15657 9551 15691
rect 13541 15691 13599 15697
rect 13541 15688 13553 15691
rect 9493 15651 9551 15657
rect 13004 15660 13553 15688
rect 5074 15620 5080 15632
rect 4479 15592 4844 15620
rect 5035 15592 5080 15620
rect 4479 15589 4491 15592
rect 4433 15583 4491 15589
rect 5074 15580 5080 15592
rect 5132 15580 5138 15632
rect 5810 15580 5816 15632
rect 5868 15580 5874 15632
rect 13004 15629 13032 15660
rect 13541 15657 13553 15660
rect 13587 15688 13599 15691
rect 13722 15688 13728 15700
rect 13587 15660 13728 15688
rect 13587 15657 13599 15660
rect 13541 15651 13599 15657
rect 13722 15648 13728 15660
rect 13780 15648 13786 15700
rect 12989 15623 13047 15629
rect 12989 15589 13001 15623
rect 13035 15589 13047 15623
rect 13262 15620 13268 15632
rect 12989 15583 13047 15589
rect 13096 15592 13268 15620
rect 3145 15555 3203 15561
rect 3145 15521 3157 15555
rect 3191 15521 3203 15555
rect 3145 15515 3203 15521
rect 3237 15555 3295 15561
rect 3237 15521 3249 15555
rect 3283 15552 3295 15555
rect 3418 15552 3424 15564
rect 3283 15524 3424 15552
rect 3283 15521 3295 15524
rect 3237 15515 3295 15521
rect 2866 15484 2872 15496
rect 2827 15456 2872 15484
rect 2866 15444 2872 15456
rect 2924 15444 2930 15496
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 3252 15484 3280 15515
rect 3418 15512 3424 15524
rect 3476 15512 3482 15564
rect 3697 15555 3755 15561
rect 3697 15521 3709 15555
rect 3743 15552 3755 15555
rect 3786 15552 3792 15564
rect 3743 15524 3792 15552
rect 3743 15521 3755 15524
rect 3697 15515 3755 15521
rect 3786 15512 3792 15524
rect 3844 15512 3850 15564
rect 4246 15561 4252 15564
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15521 4123 15555
rect 4065 15515 4123 15521
rect 4213 15555 4252 15561
rect 4213 15521 4225 15555
rect 4213 15515 4252 15521
rect 3099 15456 3280 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 3329 15419 3387 15425
rect 3329 15385 3341 15419
rect 3375 15416 3387 15419
rect 4080 15416 4108 15515
rect 4246 15512 4252 15515
rect 4304 15512 4310 15564
rect 4338 15512 4344 15564
rect 4396 15552 4402 15564
rect 4571 15555 4629 15561
rect 4396 15524 4441 15552
rect 4396 15512 4402 15524
rect 4571 15521 4583 15555
rect 4617 15552 4629 15555
rect 4706 15552 4712 15564
rect 4617 15524 4712 15552
rect 4617 15521 4629 15524
rect 4571 15515 4629 15521
rect 4706 15512 4712 15524
rect 4764 15512 4770 15564
rect 6454 15512 6460 15564
rect 6512 15552 6518 15564
rect 6733 15555 6791 15561
rect 6733 15552 6745 15555
rect 6512 15524 6745 15552
rect 6512 15512 6518 15524
rect 6733 15521 6745 15524
rect 6779 15521 6791 15555
rect 7006 15552 7012 15564
rect 6967 15524 7012 15552
rect 6733 15515 6791 15521
rect 7006 15512 7012 15524
rect 7064 15512 7070 15564
rect 9582 15552 9588 15564
rect 9543 15524 9588 15552
rect 9582 15512 9588 15524
rect 9640 15512 9646 15564
rect 12434 15512 12440 15564
rect 12492 15552 12498 15564
rect 13096 15561 13124 15592
rect 13262 15580 13268 15592
rect 13320 15620 13326 15632
rect 13320 15592 14964 15620
rect 13320 15580 13326 15592
rect 12529 15555 12587 15561
rect 12529 15552 12541 15555
rect 12492 15524 12541 15552
rect 12492 15512 12498 15524
rect 12529 15521 12541 15524
rect 12575 15521 12587 15555
rect 12529 15515 12587 15521
rect 13081 15555 13139 15561
rect 13081 15521 13093 15555
rect 13127 15521 13139 15555
rect 13538 15552 13544 15564
rect 13499 15524 13544 15552
rect 13081 15515 13139 15521
rect 4801 15487 4859 15493
rect 4801 15484 4813 15487
rect 4356 15456 4813 15484
rect 4246 15416 4252 15428
rect 3375 15388 4252 15416
rect 3375 15385 3387 15388
rect 3329 15379 3387 15385
rect 4246 15376 4252 15388
rect 4304 15376 4310 15428
rect 3234 15308 3240 15360
rect 3292 15348 3298 15360
rect 4356 15348 4384 15456
rect 4801 15453 4813 15456
rect 4847 15453 4859 15487
rect 12544 15484 12572 15515
rect 13538 15512 13544 15524
rect 13596 15512 13602 15564
rect 13814 15552 13820 15564
rect 13775 15524 13820 15552
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 14936 15561 14964 15592
rect 14369 15555 14427 15561
rect 14369 15552 14381 15555
rect 14200 15524 14381 15552
rect 14200 15496 14228 15524
rect 14369 15521 14381 15524
rect 14415 15521 14427 15555
rect 14369 15515 14427 15521
rect 14921 15555 14979 15561
rect 14921 15521 14933 15555
rect 14967 15521 14979 15555
rect 14921 15515 14979 15521
rect 15197 15555 15255 15561
rect 15197 15521 15209 15555
rect 15243 15521 15255 15555
rect 15197 15515 15255 15521
rect 13173 15487 13231 15493
rect 13173 15484 13185 15487
rect 12544 15456 13185 15484
rect 4801 15447 4859 15453
rect 13173 15453 13185 15456
rect 13219 15453 13231 15487
rect 14182 15484 14188 15496
rect 14143 15456 14188 15484
rect 13173 15447 13231 15453
rect 14182 15444 14188 15456
rect 14240 15444 14246 15496
rect 15212 15484 15240 15515
rect 14936 15456 15240 15484
rect 3292 15320 4384 15348
rect 3292 15308 3298 15320
rect 4706 15308 4712 15360
rect 4764 15348 4770 15360
rect 5258 15348 5264 15360
rect 4764 15320 5264 15348
rect 4764 15308 4770 15320
rect 5258 15308 5264 15320
rect 5316 15308 5322 15360
rect 5810 15308 5816 15360
rect 5868 15348 5874 15360
rect 6549 15351 6607 15357
rect 6549 15348 6561 15351
rect 5868 15320 6561 15348
rect 5868 15308 5874 15320
rect 6549 15317 6561 15320
rect 6595 15348 6607 15351
rect 6638 15348 6644 15360
rect 6595 15320 6644 15348
rect 6595 15317 6607 15320
rect 6549 15311 6607 15317
rect 6638 15308 6644 15320
rect 6696 15308 6702 15360
rect 14936 15357 14964 15456
rect 15010 15376 15016 15428
rect 15068 15416 15074 15428
rect 15068 15388 15113 15416
rect 15068 15376 15074 15388
rect 13817 15351 13875 15357
rect 13817 15317 13829 15351
rect 13863 15348 13875 15351
rect 14921 15351 14979 15357
rect 14921 15348 14933 15351
rect 13863 15320 14933 15348
rect 13863 15317 13875 15320
rect 13817 15311 13875 15317
rect 14921 15317 14933 15320
rect 14967 15317 14979 15351
rect 14921 15311 14979 15317
rect 1104 15258 16100 15280
rect 1104 15206 3481 15258
rect 3533 15206 3545 15258
rect 3597 15206 3609 15258
rect 3661 15206 3673 15258
rect 3725 15206 8480 15258
rect 8532 15206 8544 15258
rect 8596 15206 8608 15258
rect 8660 15206 8672 15258
rect 8724 15206 13478 15258
rect 13530 15206 13542 15258
rect 13594 15206 13606 15258
rect 13658 15206 13670 15258
rect 13722 15206 16100 15258
rect 1104 15184 16100 15206
rect 4338 15104 4344 15156
rect 4396 15144 4402 15156
rect 4982 15144 4988 15156
rect 4396 15116 4988 15144
rect 4396 15104 4402 15116
rect 4982 15104 4988 15116
rect 5040 15104 5046 15156
rect 8481 15147 8539 15153
rect 8481 15113 8493 15147
rect 8527 15144 8539 15147
rect 9125 15147 9183 15153
rect 9125 15144 9137 15147
rect 8527 15116 9137 15144
rect 8527 15113 8539 15116
rect 8481 15107 8539 15113
rect 9125 15113 9137 15116
rect 9171 15144 9183 15147
rect 9582 15144 9588 15156
rect 9171 15116 9588 15144
rect 9171 15113 9183 15116
rect 9125 15107 9183 15113
rect 9582 15104 9588 15116
rect 9640 15104 9646 15156
rect 11701 15079 11759 15085
rect 11701 15076 11713 15079
rect 8588 15048 11713 15076
rect 4614 14900 4620 14952
rect 4672 14940 4678 14952
rect 6549 14943 6607 14949
rect 6549 14940 6561 14943
rect 4672 14912 6561 14940
rect 4672 14900 4678 14912
rect 6549 14909 6561 14912
rect 6595 14940 6607 14943
rect 7650 14940 7656 14952
rect 6595 14912 7656 14940
rect 6595 14909 6607 14912
rect 6549 14903 6607 14909
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 8202 14900 8208 14952
rect 8260 14940 8266 14952
rect 8481 14943 8539 14949
rect 8481 14940 8493 14943
rect 8260 14912 8493 14940
rect 8260 14900 8266 14912
rect 8481 14909 8493 14912
rect 8527 14940 8539 14943
rect 8588 14940 8616 15048
rect 11701 15045 11713 15048
rect 11747 15045 11759 15079
rect 11701 15039 11759 15045
rect 9493 15011 9551 15017
rect 9493 15008 9505 15011
rect 9048 14980 9505 15008
rect 9048 14952 9076 14980
rect 9493 14977 9505 14980
rect 9539 14977 9551 15011
rect 9493 14971 9551 14977
rect 9030 14940 9036 14952
rect 8527 14912 8616 14940
rect 8991 14912 9036 14940
rect 8527 14909 8539 14912
rect 8481 14903 8539 14909
rect 9030 14900 9036 14912
rect 9088 14900 9094 14952
rect 9122 14900 9128 14952
rect 9180 14940 9186 14952
rect 9180 14912 9225 14940
rect 9180 14900 9186 14912
rect 4154 14832 4160 14884
rect 4212 14872 4218 14884
rect 6454 14872 6460 14884
rect 4212 14844 6460 14872
rect 4212 14832 4218 14844
rect 6454 14832 6460 14844
rect 6512 14872 6518 14884
rect 8846 14872 8852 14884
rect 6512 14844 8852 14872
rect 6512 14832 6518 14844
rect 8846 14832 8852 14844
rect 8904 14832 8910 14884
rect 11606 14832 11612 14884
rect 11664 14872 11670 14884
rect 11885 14875 11943 14881
rect 11885 14872 11897 14875
rect 11664 14844 11897 14872
rect 11664 14832 11670 14844
rect 11885 14841 11897 14844
rect 11931 14841 11943 14875
rect 11885 14835 11943 14841
rect 1104 14714 16100 14736
rect 1104 14662 5980 14714
rect 6032 14662 6044 14714
rect 6096 14662 6108 14714
rect 6160 14662 6172 14714
rect 6224 14662 10979 14714
rect 11031 14662 11043 14714
rect 11095 14662 11107 14714
rect 11159 14662 11171 14714
rect 11223 14662 16100 14714
rect 1104 14640 16100 14662
rect 4801 14603 4859 14609
rect 4801 14600 4813 14603
rect 4264 14572 4813 14600
rect 3786 14532 3792 14544
rect 2746 14504 3792 14532
rect 1946 14464 1952 14476
rect 1907 14436 1952 14464
rect 1946 14424 1952 14436
rect 2004 14464 2010 14476
rect 2746 14464 2774 14504
rect 3786 14492 3792 14504
rect 3844 14492 3850 14544
rect 4157 14535 4215 14541
rect 4157 14501 4169 14535
rect 4203 14532 4215 14535
rect 4264 14532 4292 14572
rect 4801 14569 4813 14572
rect 4847 14569 4859 14603
rect 4801 14563 4859 14569
rect 5261 14603 5319 14609
rect 5261 14569 5273 14603
rect 5307 14600 5319 14603
rect 5350 14600 5356 14612
rect 5307 14572 5356 14600
rect 5307 14569 5319 14572
rect 5261 14563 5319 14569
rect 4430 14541 4436 14544
rect 4203 14504 4292 14532
rect 4387 14535 4436 14541
rect 4203 14501 4215 14504
rect 4157 14495 4215 14501
rect 4387 14501 4399 14535
rect 4433 14501 4436 14535
rect 4387 14495 4436 14501
rect 4430 14492 4436 14495
rect 4488 14492 4494 14544
rect 4816 14532 4844 14563
rect 5350 14560 5356 14572
rect 5408 14560 5414 14612
rect 7929 14603 7987 14609
rect 7929 14600 7941 14603
rect 7392 14572 7941 14600
rect 7392 14541 7420 14572
rect 7929 14569 7941 14572
rect 7975 14600 7987 14603
rect 8297 14603 8355 14609
rect 8297 14600 8309 14603
rect 7975 14572 8309 14600
rect 7975 14569 7987 14572
rect 7929 14563 7987 14569
rect 8297 14569 8309 14572
rect 8343 14569 8355 14603
rect 8297 14563 8355 14569
rect 8389 14603 8447 14609
rect 8389 14569 8401 14603
rect 8435 14600 8447 14603
rect 9122 14600 9128 14612
rect 8435 14572 9128 14600
rect 8435 14569 8447 14572
rect 8389 14563 8447 14569
rect 9122 14560 9128 14572
rect 9180 14560 9186 14612
rect 11606 14600 11612 14612
rect 10980 14572 11612 14600
rect 10980 14541 11008 14572
rect 11606 14560 11612 14572
rect 11664 14560 11670 14612
rect 13633 14603 13691 14609
rect 13633 14569 13645 14603
rect 13679 14600 13691 14603
rect 13814 14600 13820 14612
rect 13679 14572 13820 14600
rect 13679 14569 13691 14572
rect 13633 14563 13691 14569
rect 13814 14560 13820 14572
rect 13872 14600 13878 14612
rect 14369 14603 14427 14609
rect 14369 14600 14381 14603
rect 13872 14572 14381 14600
rect 13872 14560 13878 14572
rect 14369 14569 14381 14572
rect 14415 14569 14427 14603
rect 14369 14563 14427 14569
rect 7377 14535 7435 14541
rect 4816 14504 5304 14532
rect 2004 14436 2774 14464
rect 3421 14467 3479 14473
rect 2004 14424 2010 14436
rect 3421 14433 3433 14467
rect 3467 14433 3479 14467
rect 3421 14427 3479 14433
rect 3513 14467 3571 14473
rect 3513 14433 3525 14467
rect 3559 14464 3571 14467
rect 3970 14464 3976 14476
rect 3559 14436 3976 14464
rect 3559 14433 3571 14436
rect 3513 14427 3571 14433
rect 3436 14396 3464 14427
rect 3970 14424 3976 14436
rect 4028 14424 4034 14476
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 4249 14467 4307 14473
rect 4111 14436 4200 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 3436 14368 4108 14396
rect 4080 14340 4108 14368
rect 4062 14288 4068 14340
rect 4120 14288 4126 14340
rect 2133 14263 2191 14269
rect 2133 14229 2145 14263
rect 2179 14260 2191 14263
rect 2222 14260 2228 14272
rect 2179 14232 2228 14260
rect 2179 14229 2191 14232
rect 2133 14223 2191 14229
rect 2222 14220 2228 14232
rect 2280 14220 2286 14272
rect 3326 14260 3332 14272
rect 3287 14232 3332 14260
rect 3326 14220 3332 14232
rect 3384 14220 3390 14272
rect 3605 14263 3663 14269
rect 3605 14229 3617 14263
rect 3651 14260 3663 14263
rect 3786 14260 3792 14272
rect 3651 14232 3792 14260
rect 3651 14229 3663 14232
rect 3605 14223 3663 14229
rect 3786 14220 3792 14232
rect 3844 14220 3850 14272
rect 3878 14220 3884 14272
rect 3936 14260 3942 14272
rect 4172 14260 4200 14436
rect 4249 14433 4261 14467
rect 4295 14433 4307 14467
rect 4985 14467 5043 14473
rect 4985 14464 4997 14467
rect 4249 14427 4307 14433
rect 4816 14436 4997 14464
rect 4264 14396 4292 14427
rect 4338 14396 4344 14408
rect 4264 14368 4344 14396
rect 4338 14356 4344 14368
rect 4396 14356 4402 14408
rect 4525 14399 4583 14405
rect 4525 14365 4537 14399
rect 4571 14365 4583 14399
rect 4525 14359 4583 14365
rect 4246 14288 4252 14340
rect 4304 14328 4310 14340
rect 4540 14328 4568 14359
rect 4304 14300 4568 14328
rect 4816 14328 4844 14436
rect 4985 14433 4997 14436
rect 5031 14433 5043 14467
rect 4985 14427 5043 14433
rect 5169 14467 5227 14473
rect 5169 14433 5181 14467
rect 5215 14433 5227 14467
rect 5169 14427 5227 14433
rect 4890 14356 4896 14408
rect 4948 14396 4954 14408
rect 5184 14396 5212 14427
rect 5276 14405 5304 14504
rect 7377 14501 7389 14535
rect 7423 14501 7435 14535
rect 7377 14495 7435 14501
rect 10965 14535 11023 14541
rect 10965 14501 10977 14535
rect 11011 14501 11023 14535
rect 10965 14495 11023 14501
rect 13173 14535 13231 14541
rect 13173 14501 13185 14535
rect 13219 14532 13231 14535
rect 14182 14532 14188 14544
rect 13219 14504 14188 14532
rect 13219 14501 13231 14504
rect 13173 14495 13231 14501
rect 14182 14492 14188 14504
rect 14240 14492 14246 14544
rect 5537 14467 5595 14473
rect 5537 14433 5549 14467
rect 5583 14464 5595 14467
rect 5718 14464 5724 14476
rect 5583 14436 5724 14464
rect 5583 14433 5595 14436
rect 5537 14427 5595 14433
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 6917 14467 6975 14473
rect 6917 14433 6929 14467
rect 6963 14433 6975 14467
rect 6917 14427 6975 14433
rect 7469 14467 7527 14473
rect 7469 14433 7481 14467
rect 7515 14464 7527 14467
rect 8202 14464 8208 14476
rect 7515 14436 8208 14464
rect 7515 14433 7527 14436
rect 7469 14427 7527 14433
rect 4948 14368 5212 14396
rect 5261 14399 5319 14405
rect 4948 14356 4954 14368
rect 5261 14365 5273 14399
rect 5307 14365 5319 14399
rect 5261 14359 5319 14365
rect 5350 14356 5356 14408
rect 5408 14396 5414 14408
rect 5445 14399 5503 14405
rect 5445 14396 5457 14399
rect 5408 14368 5457 14396
rect 5408 14356 5414 14368
rect 5445 14365 5457 14368
rect 5491 14365 5503 14399
rect 6932 14396 6960 14427
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 10505 14467 10563 14473
rect 10505 14433 10517 14467
rect 10551 14433 10563 14467
rect 10505 14427 10563 14433
rect 11057 14467 11115 14473
rect 11057 14433 11069 14467
rect 11103 14464 11115 14467
rect 11330 14464 11336 14476
rect 11103 14436 11336 14464
rect 11103 14433 11115 14436
rect 11057 14427 11115 14433
rect 7558 14396 7564 14408
rect 6932 14368 7564 14396
rect 5445 14359 5503 14365
rect 7558 14356 7564 14368
rect 7616 14356 7622 14408
rect 10520 14396 10548 14427
rect 11330 14424 11336 14436
rect 11388 14424 11394 14476
rect 12158 14424 12164 14476
rect 12216 14464 12222 14476
rect 12805 14467 12863 14473
rect 12805 14464 12817 14467
rect 12216 14436 12817 14464
rect 12216 14424 12222 14436
rect 12805 14433 12817 14436
rect 12851 14433 12863 14467
rect 12986 14464 12992 14476
rect 12947 14436 12992 14464
rect 12805 14427 12863 14433
rect 12986 14424 12992 14436
rect 13044 14424 13050 14476
rect 11241 14399 11299 14405
rect 11241 14396 11253 14399
rect 10520 14368 11253 14396
rect 11241 14365 11253 14368
rect 11287 14396 11299 14399
rect 12176 14396 12204 14424
rect 11287 14368 12204 14396
rect 13265 14399 13323 14405
rect 11287 14365 11299 14368
rect 11241 14359 11299 14365
rect 13265 14365 13277 14399
rect 13311 14396 13323 14399
rect 13354 14396 13360 14408
rect 13311 14368 13360 14396
rect 13311 14365 13323 14368
rect 13265 14359 13323 14365
rect 13354 14356 13360 14368
rect 13412 14356 13418 14408
rect 5534 14328 5540 14340
rect 4816 14300 5540 14328
rect 4304 14288 4310 14300
rect 5534 14288 5540 14300
rect 5592 14288 5598 14340
rect 7929 14331 7987 14337
rect 7929 14297 7941 14331
rect 7975 14328 7987 14331
rect 8021 14331 8079 14337
rect 8021 14328 8033 14331
rect 7975 14300 8033 14328
rect 7975 14297 7987 14300
rect 7929 14291 7987 14297
rect 8021 14297 8033 14300
rect 8067 14297 8079 14331
rect 8021 14291 8079 14297
rect 11609 14331 11667 14337
rect 11609 14297 11621 14331
rect 11655 14328 11667 14331
rect 11790 14328 11796 14340
rect 11655 14300 11796 14328
rect 11655 14297 11667 14300
rect 11609 14291 11667 14297
rect 11790 14288 11796 14300
rect 11848 14288 11854 14340
rect 13633 14331 13691 14337
rect 13633 14297 13645 14331
rect 13679 14328 13691 14331
rect 13906 14328 13912 14340
rect 13679 14300 13912 14328
rect 13679 14297 13691 14300
rect 13633 14291 13691 14297
rect 13906 14288 13912 14300
rect 13964 14288 13970 14340
rect 5626 14260 5632 14272
rect 3936 14232 3981 14260
rect 4172 14232 5632 14260
rect 3936 14220 3942 14232
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 14461 14263 14519 14269
rect 14461 14229 14473 14263
rect 14507 14260 14519 14263
rect 14826 14260 14832 14272
rect 14507 14232 14832 14260
rect 14507 14229 14519 14232
rect 14461 14223 14519 14229
rect 14826 14220 14832 14232
rect 14884 14220 14890 14272
rect 1104 14170 16100 14192
rect 1104 14118 3481 14170
rect 3533 14118 3545 14170
rect 3597 14118 3609 14170
rect 3661 14118 3673 14170
rect 3725 14118 8480 14170
rect 8532 14118 8544 14170
rect 8596 14118 8608 14170
rect 8660 14118 8672 14170
rect 8724 14118 13478 14170
rect 13530 14118 13542 14170
rect 13594 14118 13606 14170
rect 13658 14118 13670 14170
rect 13722 14118 16100 14170
rect 1104 14096 16100 14118
rect 5905 14059 5963 14065
rect 5905 14056 5917 14059
rect 5092 14028 5917 14056
rect 3878 13988 3884 14000
rect 3252 13960 3884 13988
rect 2961 13923 3019 13929
rect 2961 13889 2973 13923
rect 3007 13920 3019 13923
rect 3252 13920 3280 13960
rect 3878 13948 3884 13960
rect 3936 13948 3942 14000
rect 4062 13988 4068 14000
rect 3988 13960 4068 13988
rect 3007 13892 3280 13920
rect 3007 13889 3019 13892
rect 2961 13883 3019 13889
rect 3326 13880 3332 13932
rect 3384 13920 3390 13932
rect 3988 13920 4016 13960
rect 4062 13948 4068 13960
rect 4120 13988 4126 14000
rect 4709 13991 4767 13997
rect 4709 13988 4721 13991
rect 4120 13960 4721 13988
rect 4120 13948 4126 13960
rect 4709 13957 4721 13960
rect 4755 13957 4767 13991
rect 4982 13988 4988 14000
rect 4943 13960 4988 13988
rect 4709 13951 4767 13957
rect 4982 13948 4988 13960
rect 5040 13948 5046 14000
rect 3384 13892 3648 13920
rect 3384 13880 3390 13892
rect 3234 13812 3240 13864
rect 3292 13852 3298 13864
rect 3620 13861 3648 13892
rect 3712 13892 4016 13920
rect 3712 13861 3740 13892
rect 4154 13880 4160 13932
rect 4212 13880 4218 13932
rect 4525 13923 4583 13929
rect 4525 13889 4537 13923
rect 4571 13920 4583 13923
rect 5092 13920 5120 14028
rect 5905 14025 5917 14028
rect 5951 14025 5963 14059
rect 5905 14019 5963 14025
rect 7006 14016 7012 14068
rect 7064 14056 7070 14068
rect 7101 14059 7159 14065
rect 7101 14056 7113 14059
rect 7064 14028 7113 14056
rect 7064 14016 7070 14028
rect 7101 14025 7113 14028
rect 7147 14025 7159 14059
rect 7101 14019 7159 14025
rect 9030 14016 9036 14068
rect 9088 14056 9094 14068
rect 9217 14059 9275 14065
rect 9217 14056 9229 14059
rect 9088 14028 9229 14056
rect 9088 14016 9094 14028
rect 9217 14025 9229 14028
rect 9263 14025 9275 14059
rect 9217 14019 9275 14025
rect 9398 14016 9404 14068
rect 9456 14056 9462 14068
rect 9585 14059 9643 14065
rect 9585 14056 9597 14059
rect 9456 14028 9597 14056
rect 9456 14016 9462 14028
rect 9585 14025 9597 14028
rect 9631 14056 9643 14059
rect 11790 14056 11796 14068
rect 9631 14028 10916 14056
rect 11751 14028 11796 14056
rect 9631 14025 9643 14028
rect 9585 14019 9643 14025
rect 7024 13988 7052 14016
rect 9766 13988 9772 14000
rect 5184 13960 7052 13988
rect 9727 13960 9772 13988
rect 5184 13929 5212 13960
rect 9766 13948 9772 13960
rect 9824 13948 9830 14000
rect 10888 13988 10916 14028
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 13906 14056 13912 14068
rect 13867 14028 13912 14056
rect 13906 14016 13912 14028
rect 13964 14016 13970 14068
rect 12066 13988 12072 14000
rect 10888 13960 12072 13988
rect 12066 13948 12072 13960
rect 12124 13988 12130 14000
rect 12986 13988 12992 14000
rect 12124 13960 12992 13988
rect 12124 13948 12130 13960
rect 12986 13948 12992 13960
rect 13044 13948 13050 14000
rect 13725 13991 13783 13997
rect 13725 13957 13737 13991
rect 13771 13988 13783 13991
rect 13814 13988 13820 14000
rect 13771 13960 13820 13988
rect 13771 13957 13783 13960
rect 13725 13951 13783 13957
rect 13814 13948 13820 13960
rect 13872 13948 13878 14000
rect 14826 13988 14832 14000
rect 14787 13960 14832 13988
rect 14826 13948 14832 13960
rect 14884 13948 14890 14000
rect 4571 13892 5120 13920
rect 5169 13923 5227 13929
rect 4571 13889 4583 13892
rect 4525 13883 4583 13889
rect 3508 13855 3566 13861
rect 3292 13824 3337 13852
rect 3292 13812 3298 13824
rect 3508 13821 3520 13855
rect 3554 13821 3566 13855
rect 3508 13815 3566 13821
rect 3605 13855 3663 13861
rect 3605 13821 3617 13855
rect 3651 13821 3663 13855
rect 3605 13815 3663 13821
rect 3697 13855 3755 13861
rect 3697 13821 3709 13855
rect 3743 13821 3755 13855
rect 3697 13815 3755 13821
rect 2222 13744 2228 13796
rect 2280 13744 2286 13796
rect 1486 13716 1492 13728
rect 1447 13688 1492 13716
rect 1486 13676 1492 13688
rect 1544 13676 1550 13728
rect 2866 13676 2872 13728
rect 2924 13716 2930 13728
rect 3329 13719 3387 13725
rect 3329 13716 3341 13719
rect 2924 13688 3341 13716
rect 2924 13676 2930 13688
rect 3329 13685 3341 13688
rect 3375 13685 3387 13719
rect 3528 13716 3556 13815
rect 3786 13812 3792 13864
rect 3844 13861 3850 13864
rect 3844 13855 3883 13861
rect 3871 13821 3883 13855
rect 3844 13815 3883 13821
rect 3973 13855 4031 13861
rect 3973 13821 3985 13855
rect 4019 13852 4031 13855
rect 4062 13852 4068 13864
rect 4019 13824 4068 13852
rect 4019 13821 4031 13824
rect 3973 13815 4031 13821
rect 3844 13812 3850 13815
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 4172 13852 4200 13880
rect 4724 13864 4752 13892
rect 5169 13889 5181 13923
rect 5215 13889 5227 13923
rect 5534 13920 5540 13932
rect 5169 13883 5227 13889
rect 5276 13892 5540 13920
rect 4249 13855 4307 13861
rect 4249 13852 4261 13855
rect 4172 13824 4261 13852
rect 4249 13821 4261 13824
rect 4295 13821 4307 13855
rect 4249 13815 4307 13821
rect 4341 13855 4399 13861
rect 4341 13821 4353 13855
rect 4387 13821 4399 13855
rect 4614 13852 4620 13864
rect 4575 13824 4620 13852
rect 4341 13815 4399 13821
rect 4356 13784 4384 13815
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 4706 13812 4712 13864
rect 4764 13812 4770 13864
rect 4890 13852 4896 13864
rect 4851 13824 4896 13852
rect 4890 13812 4896 13824
rect 4948 13812 4954 13864
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13852 5135 13855
rect 5276 13852 5304 13892
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 5810 13920 5816 13932
rect 5644 13892 5816 13920
rect 5123 13824 5304 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 5350 13812 5356 13864
rect 5408 13852 5414 13864
rect 5644 13861 5672 13892
rect 5810 13880 5816 13892
rect 5868 13880 5874 13932
rect 9214 13920 9220 13932
rect 7024 13892 9220 13920
rect 7024 13864 7052 13892
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 9306 13880 9312 13932
rect 9364 13920 9370 13932
rect 9677 13923 9735 13929
rect 9677 13920 9689 13923
rect 9364 13892 9689 13920
rect 9364 13880 9370 13892
rect 9677 13889 9689 13892
rect 9723 13889 9735 13923
rect 9677 13883 9735 13889
rect 14108 13892 14780 13920
rect 5629 13855 5687 13861
rect 5408 13824 5453 13852
rect 5408 13812 5414 13824
rect 5629 13821 5641 13855
rect 5675 13821 5687 13855
rect 5629 13815 5687 13821
rect 5721 13855 5779 13861
rect 5721 13821 5733 13855
rect 5767 13821 5779 13855
rect 5721 13815 5779 13821
rect 5997 13855 6055 13861
rect 5997 13821 6009 13855
rect 6043 13852 6055 13855
rect 6546 13852 6552 13864
rect 6043 13824 6552 13852
rect 6043 13821 6055 13824
rect 5997 13815 6055 13821
rect 5368 13784 5396 13812
rect 5736 13784 5764 13815
rect 6546 13812 6552 13824
rect 6604 13852 6610 13864
rect 7006 13852 7012 13864
rect 6604 13824 7012 13852
rect 6604 13812 6610 13824
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 7190 13852 7196 13864
rect 7151 13824 7196 13852
rect 7190 13812 7196 13824
rect 7248 13812 7254 13864
rect 9490 13852 9496 13864
rect 9451 13824 9496 13852
rect 9490 13812 9496 13824
rect 9548 13812 9554 13864
rect 9950 13852 9956 13864
rect 9911 13824 9956 13852
rect 9950 13812 9956 13824
rect 10008 13852 10014 13864
rect 13078 13852 13084 13864
rect 10008 13824 13084 13852
rect 10008 13812 10014 13824
rect 13078 13812 13084 13824
rect 13136 13812 13142 13864
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13852 13231 13855
rect 13354 13852 13360 13864
rect 13219 13824 13360 13852
rect 13219 13821 13231 13824
rect 13173 13815 13231 13821
rect 13354 13812 13360 13824
rect 13412 13812 13418 13864
rect 14108 13861 14136 13892
rect 13725 13855 13783 13861
rect 13725 13821 13737 13855
rect 13771 13852 13783 13855
rect 14093 13855 14151 13861
rect 14093 13852 14105 13855
rect 13771 13824 14105 13852
rect 13771 13821 13783 13824
rect 13725 13815 13783 13821
rect 14093 13821 14105 13824
rect 14139 13821 14151 13855
rect 14093 13815 14151 13821
rect 14185 13855 14243 13861
rect 14185 13821 14197 13855
rect 14231 13821 14243 13855
rect 14642 13852 14648 13864
rect 14603 13824 14648 13852
rect 14185 13815 14243 13821
rect 4356 13756 5764 13784
rect 10134 13744 10140 13796
rect 10192 13784 10198 13796
rect 14200 13784 14228 13815
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 14752 13861 14780 13892
rect 14737 13855 14795 13861
rect 14737 13821 14749 13855
rect 14783 13852 14795 13855
rect 15010 13852 15016 13864
rect 14783 13824 15016 13852
rect 14783 13821 14795 13824
rect 14737 13815 14795 13821
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 15197 13855 15255 13861
rect 15197 13821 15209 13855
rect 15243 13821 15255 13855
rect 15197 13815 15255 13821
rect 15212 13784 15240 13815
rect 10192 13756 15240 13784
rect 10192 13744 10198 13756
rect 3970 13716 3976 13728
rect 3528 13688 3976 13716
rect 3329 13679 3387 13685
rect 3970 13676 3976 13688
rect 4028 13716 4034 13728
rect 4065 13719 4123 13725
rect 4065 13716 4077 13719
rect 4028 13688 4077 13716
rect 4028 13676 4034 13688
rect 4065 13685 4077 13688
rect 4111 13685 4123 13719
rect 4065 13679 4123 13685
rect 4982 13676 4988 13728
rect 5040 13716 5046 13728
rect 5445 13719 5503 13725
rect 5445 13716 5457 13719
rect 5040 13688 5457 13716
rect 5040 13676 5046 13688
rect 5445 13685 5457 13688
rect 5491 13685 5503 13719
rect 11698 13716 11704 13728
rect 11659 13688 11704 13716
rect 5445 13679 5503 13685
rect 11698 13676 11704 13688
rect 11756 13676 11762 13728
rect 14642 13676 14648 13728
rect 14700 13716 14706 13728
rect 14829 13719 14887 13725
rect 14829 13716 14841 13719
rect 14700 13688 14841 13716
rect 14700 13676 14706 13688
rect 14829 13685 14841 13688
rect 14875 13685 14887 13719
rect 14829 13679 14887 13685
rect 1104 13626 16100 13648
rect 1104 13574 5980 13626
rect 6032 13574 6044 13626
rect 6096 13574 6108 13626
rect 6160 13574 6172 13626
rect 6224 13574 10979 13626
rect 11031 13574 11043 13626
rect 11095 13574 11107 13626
rect 11159 13574 11171 13626
rect 11223 13574 16100 13626
rect 1104 13552 16100 13574
rect 4801 13515 4859 13521
rect 4801 13481 4813 13515
rect 4847 13512 4859 13515
rect 4890 13512 4896 13524
rect 4847 13484 4896 13512
rect 4847 13481 4859 13484
rect 4801 13475 4859 13481
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 5626 13512 5632 13524
rect 5587 13484 5632 13512
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 5810 13472 5816 13524
rect 5868 13512 5874 13524
rect 7742 13512 7748 13524
rect 5868 13484 7748 13512
rect 5868 13472 5874 13484
rect 4908 13444 4936 13472
rect 4908 13416 5488 13444
rect 4706 13336 4712 13388
rect 4764 13376 4770 13388
rect 4985 13379 5043 13385
rect 4985 13376 4997 13379
rect 4764 13348 4997 13376
rect 4764 13336 4770 13348
rect 4985 13345 4997 13348
rect 5031 13345 5043 13379
rect 4985 13339 5043 13345
rect 5077 13379 5135 13385
rect 5077 13345 5089 13379
rect 5123 13345 5135 13379
rect 5077 13339 5135 13345
rect 5169 13379 5227 13385
rect 5169 13345 5181 13379
rect 5215 13345 5227 13379
rect 5350 13376 5356 13388
rect 5311 13348 5356 13376
rect 5169 13339 5227 13345
rect 1486 13268 1492 13320
rect 1544 13308 1550 13320
rect 4430 13308 4436 13320
rect 1544 13280 4436 13308
rect 1544 13268 1550 13280
rect 4430 13268 4436 13280
rect 4488 13308 4494 13320
rect 5092 13308 5120 13339
rect 4488 13280 5120 13308
rect 5184 13308 5212 13339
rect 5350 13336 5356 13348
rect 5408 13336 5414 13388
rect 5460 13385 5488 13416
rect 5445 13379 5503 13385
rect 5445 13345 5457 13379
rect 5491 13345 5503 13379
rect 5445 13339 5503 13345
rect 5534 13336 5540 13388
rect 5592 13376 5598 13388
rect 5629 13379 5687 13385
rect 5629 13376 5641 13379
rect 5592 13348 5641 13376
rect 5592 13336 5598 13348
rect 5629 13345 5641 13348
rect 5675 13345 5687 13379
rect 6270 13376 6276 13388
rect 6231 13348 6276 13376
rect 5629 13339 5687 13345
rect 6270 13336 6276 13348
rect 6328 13376 6334 13388
rect 7116 13385 7144 13484
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 9766 13512 9772 13524
rect 8036 13484 9772 13512
rect 6917 13379 6975 13385
rect 6917 13376 6929 13379
rect 6328 13348 6929 13376
rect 6328 13336 6334 13348
rect 6917 13345 6929 13348
rect 6963 13345 6975 13379
rect 6917 13339 6975 13345
rect 7101 13379 7159 13385
rect 7101 13345 7113 13379
rect 7147 13376 7159 13379
rect 7837 13379 7895 13385
rect 7147 13348 7788 13376
rect 7147 13345 7159 13348
rect 7101 13339 7159 13345
rect 5718 13308 5724 13320
rect 5184 13280 5724 13308
rect 4488 13268 4494 13280
rect 5092 13240 5120 13280
rect 5718 13268 5724 13280
rect 5776 13308 5782 13320
rect 6365 13311 6423 13317
rect 6365 13308 6377 13311
rect 5776 13280 6377 13308
rect 5776 13268 5782 13280
rect 6365 13277 6377 13280
rect 6411 13308 6423 13311
rect 6546 13308 6552 13320
rect 6411 13280 6552 13308
rect 6411 13277 6423 13280
rect 6365 13271 6423 13277
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 6270 13240 6276 13252
rect 5092 13212 6276 13240
rect 6270 13200 6276 13212
rect 6328 13200 6334 13252
rect 6932 13240 6960 13339
rect 7650 13308 7656 13320
rect 7611 13280 7656 13308
rect 7650 13268 7656 13280
rect 7708 13268 7714 13320
rect 7760 13317 7788 13348
rect 7837 13345 7849 13379
rect 7883 13376 7895 13379
rect 8036 13376 8064 13484
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 11609 13515 11667 13521
rect 11609 13481 11621 13515
rect 11655 13512 11667 13515
rect 11698 13512 11704 13524
rect 11655 13484 11704 13512
rect 11655 13481 11667 13484
rect 11609 13475 11667 13481
rect 9493 13447 9551 13453
rect 9493 13444 9505 13447
rect 8588 13416 9505 13444
rect 7883 13348 8064 13376
rect 7883 13345 7895 13348
rect 7837 13339 7895 13345
rect 7753 13311 7811 13317
rect 7753 13277 7765 13311
rect 7799 13277 7811 13311
rect 7753 13271 7811 13277
rect 7852 13240 7880 13339
rect 8294 13336 8300 13388
rect 8352 13376 8358 13388
rect 8588 13385 8616 13416
rect 9493 13413 9505 13416
rect 9539 13413 9551 13447
rect 9493 13407 9551 13413
rect 11057 13447 11115 13453
rect 11057 13413 11069 13447
rect 11103 13444 11115 13447
rect 11624 13444 11652 13475
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 13354 13512 13360 13524
rect 13315 13484 13360 13512
rect 13354 13472 13360 13484
rect 13412 13472 13418 13524
rect 11103 13416 11652 13444
rect 12161 13447 12219 13453
rect 11103 13413 11115 13416
rect 11057 13407 11115 13413
rect 12161 13413 12173 13447
rect 12207 13444 12219 13447
rect 12250 13444 12256 13456
rect 12207 13416 12256 13444
rect 12207 13413 12219 13416
rect 12161 13407 12219 13413
rect 12250 13404 12256 13416
rect 12308 13404 12314 13456
rect 14642 13404 14648 13456
rect 14700 13444 14706 13456
rect 15289 13447 15347 13453
rect 15289 13444 15301 13447
rect 14700 13416 15301 13444
rect 14700 13404 14706 13416
rect 15289 13413 15301 13416
rect 15335 13413 15347 13447
rect 15289 13407 15347 13413
rect 8573 13379 8631 13385
rect 8573 13376 8585 13379
rect 8352 13348 8585 13376
rect 8352 13336 8358 13348
rect 8573 13345 8585 13348
rect 8619 13345 8631 13379
rect 8846 13376 8852 13388
rect 8807 13348 8852 13376
rect 8573 13339 8631 13345
rect 8846 13336 8852 13348
rect 8904 13336 8910 13388
rect 9030 13336 9036 13388
rect 9088 13376 9094 13388
rect 9401 13379 9459 13385
rect 9401 13376 9413 13379
rect 9088 13348 9413 13376
rect 9088 13336 9094 13348
rect 9401 13345 9413 13348
rect 9447 13345 9459 13379
rect 10042 13376 10048 13388
rect 9401 13339 9459 13345
rect 9646 13348 10048 13376
rect 7926 13268 7932 13320
rect 7984 13308 7990 13320
rect 9306 13308 9312 13320
rect 7984 13280 8029 13308
rect 9267 13280 9312 13308
rect 7984 13268 7990 13280
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 6932 13212 7880 13240
rect 8113 13243 8171 13249
rect 8113 13209 8125 13243
rect 8159 13240 8171 13243
rect 9646 13240 9674 13348
rect 10042 13336 10048 13348
rect 10100 13336 10106 13388
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13345 10195 13379
rect 10137 13339 10195 13345
rect 10597 13379 10655 13385
rect 10597 13345 10609 13379
rect 10643 13345 10655 13379
rect 10597 13339 10655 13345
rect 11149 13379 11207 13385
rect 11149 13345 11161 13379
rect 11195 13376 11207 13379
rect 11330 13376 11336 13388
rect 11195 13348 11336 13376
rect 11195 13345 11207 13348
rect 11149 13339 11207 13345
rect 9953 13311 10011 13317
rect 9953 13277 9965 13311
rect 9999 13277 10011 13311
rect 9953 13271 10011 13277
rect 8159 13212 9674 13240
rect 9861 13243 9919 13249
rect 8159 13209 8171 13212
rect 8113 13203 8171 13209
rect 9861 13209 9873 13243
rect 9907 13240 9919 13243
rect 9968 13240 9996 13271
rect 9907 13212 9996 13240
rect 10152 13240 10180 13339
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 10612 13308 10640 13339
rect 11330 13336 11336 13348
rect 11388 13376 11394 13388
rect 11885 13379 11943 13385
rect 11885 13376 11897 13379
rect 11388 13348 11897 13376
rect 11388 13336 11394 13348
rect 11885 13345 11897 13348
rect 11931 13345 11943 13379
rect 12342 13376 12348 13388
rect 12303 13348 12348 13376
rect 11885 13339 11943 13345
rect 12342 13336 12348 13348
rect 12400 13336 12406 13388
rect 12710 13336 12716 13388
rect 12768 13376 12774 13388
rect 12861 13379 12919 13385
rect 12861 13376 12873 13379
rect 12768 13348 12873 13376
rect 12768 13336 12774 13348
rect 12861 13345 12873 13348
rect 12907 13345 12919 13379
rect 12986 13376 12992 13388
rect 12947 13348 12992 13376
rect 12861 13339 12919 13345
rect 12986 13336 12992 13348
rect 13044 13336 13050 13388
rect 13078 13336 13084 13388
rect 13136 13376 13142 13388
rect 13173 13379 13231 13385
rect 13173 13376 13185 13379
rect 13136 13348 13185 13376
rect 13136 13336 13142 13348
rect 13173 13345 13185 13348
rect 13219 13345 13231 13379
rect 13173 13339 13231 13345
rect 11241 13311 11299 13317
rect 11241 13308 11253 13311
rect 10367 13280 11253 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 11241 13277 11253 13280
rect 11287 13277 11299 13311
rect 12434 13308 12440 13320
rect 11241 13271 11299 13277
rect 11348 13280 12440 13308
rect 11348 13240 11376 13280
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 10152 13212 11376 13240
rect 11609 13243 11667 13249
rect 9907 13209 9919 13212
rect 9861 13203 9919 13209
rect 7190 13172 7196 13184
rect 7151 13144 7196 13172
rect 7190 13132 7196 13144
rect 7248 13132 7254 13184
rect 8665 13175 8723 13181
rect 8665 13141 8677 13175
rect 8711 13172 8723 13175
rect 10152 13172 10180 13212
rect 11609 13209 11621 13243
rect 11655 13240 11667 13243
rect 11701 13243 11759 13249
rect 11701 13240 11713 13243
rect 11655 13212 11713 13240
rect 11655 13209 11667 13212
rect 11609 13203 11667 13209
rect 11701 13209 11713 13212
rect 11747 13209 11759 13243
rect 11701 13203 11759 13209
rect 12802 13200 12808 13252
rect 12860 13240 12866 13252
rect 13081 13243 13139 13249
rect 13081 13240 13093 13243
rect 12860 13212 13093 13240
rect 12860 13200 12866 13212
rect 13081 13209 13093 13212
rect 13127 13209 13139 13243
rect 13081 13203 13139 13209
rect 14918 13200 14924 13252
rect 14976 13240 14982 13252
rect 15105 13243 15163 13249
rect 15105 13240 15117 13243
rect 14976 13212 15117 13240
rect 14976 13200 14982 13212
rect 15105 13209 15117 13212
rect 15151 13209 15163 13243
rect 15105 13203 15163 13209
rect 8711 13144 10180 13172
rect 8711 13141 8723 13144
rect 8665 13135 8723 13141
rect 12158 13132 12164 13184
rect 12216 13172 12222 13184
rect 12437 13175 12495 13181
rect 12437 13172 12449 13175
rect 12216 13144 12449 13172
rect 12216 13132 12222 13144
rect 12437 13141 12449 13144
rect 12483 13141 12495 13175
rect 12437 13135 12495 13141
rect 1104 13082 16100 13104
rect 1104 13030 3481 13082
rect 3533 13030 3545 13082
rect 3597 13030 3609 13082
rect 3661 13030 3673 13082
rect 3725 13030 8480 13082
rect 8532 13030 8544 13082
rect 8596 13030 8608 13082
rect 8660 13030 8672 13082
rect 8724 13030 13478 13082
rect 13530 13030 13542 13082
rect 13594 13030 13606 13082
rect 13658 13030 13670 13082
rect 13722 13030 16100 13082
rect 1104 13008 16100 13030
rect 7650 12928 7656 12980
rect 7708 12968 7714 12980
rect 8018 12968 8024 12980
rect 7708 12940 8024 12968
rect 7708 12928 7714 12940
rect 8018 12928 8024 12940
rect 8076 12968 8082 12980
rect 9306 12968 9312 12980
rect 8076 12940 9312 12968
rect 8076 12928 8082 12940
rect 9306 12928 9312 12940
rect 9364 12928 9370 12980
rect 9766 12928 9772 12980
rect 9824 12968 9830 12980
rect 12802 12968 12808 12980
rect 9824 12940 12808 12968
rect 9824 12928 9830 12940
rect 12802 12928 12808 12940
rect 12860 12928 12866 12980
rect 7926 12900 7932 12912
rect 7760 12872 7932 12900
rect 7650 12832 7656 12844
rect 5828 12804 7656 12832
rect 1946 12724 1952 12776
rect 2004 12764 2010 12776
rect 2317 12767 2375 12773
rect 2317 12764 2329 12767
rect 2004 12736 2329 12764
rect 2004 12724 2010 12736
rect 2317 12733 2329 12736
rect 2363 12733 2375 12767
rect 2317 12727 2375 12733
rect 3510 12724 3516 12776
rect 3568 12764 3574 12776
rect 3697 12767 3755 12773
rect 3697 12764 3709 12767
rect 3568 12736 3709 12764
rect 3568 12724 3574 12736
rect 3697 12733 3709 12736
rect 3743 12764 3755 12767
rect 5442 12764 5448 12776
rect 3743 12736 5448 12764
rect 3743 12733 3755 12736
rect 3697 12727 3755 12733
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 5828 12773 5856 12804
rect 7650 12792 7656 12804
rect 7708 12792 7714 12844
rect 7760 12841 7788 12872
rect 7926 12860 7932 12872
rect 7984 12900 7990 12912
rect 8478 12900 8484 12912
rect 7984 12872 8484 12900
rect 7984 12860 7990 12872
rect 8478 12860 8484 12872
rect 8536 12860 8542 12912
rect 13725 12903 13783 12909
rect 13725 12869 13737 12903
rect 13771 12900 13783 12903
rect 14093 12903 14151 12909
rect 14093 12900 14105 12903
rect 13771 12872 14105 12900
rect 13771 12869 13783 12872
rect 13725 12863 13783 12869
rect 14093 12869 14105 12872
rect 14139 12869 14151 12903
rect 14093 12863 14151 12869
rect 7745 12835 7803 12841
rect 7745 12801 7757 12835
rect 7791 12801 7803 12835
rect 9398 12832 9404 12844
rect 7745 12795 7803 12801
rect 7944 12804 9404 12832
rect 5629 12767 5687 12773
rect 5629 12733 5641 12767
rect 5675 12733 5687 12767
rect 5629 12727 5687 12733
rect 5813 12767 5871 12773
rect 5813 12733 5825 12767
rect 5859 12733 5871 12767
rect 6546 12764 6552 12776
rect 6507 12736 6552 12764
rect 5813 12727 5871 12733
rect 3878 12696 3884 12708
rect 3839 12668 3884 12696
rect 3878 12656 3884 12668
rect 3936 12656 3942 12708
rect 5166 12656 5172 12708
rect 5224 12696 5230 12708
rect 5644 12696 5672 12727
rect 6546 12724 6552 12736
rect 6604 12724 6610 12776
rect 6733 12767 6791 12773
rect 6733 12733 6745 12767
rect 6779 12733 6791 12767
rect 7098 12764 7104 12776
rect 7059 12736 7104 12764
rect 6733 12727 6791 12733
rect 6270 12696 6276 12708
rect 5224 12668 6276 12696
rect 5224 12656 5230 12668
rect 6270 12656 6276 12668
rect 6328 12656 6334 12708
rect 2133 12631 2191 12637
rect 2133 12597 2145 12631
rect 2179 12628 2191 12631
rect 2222 12628 2228 12640
rect 2179 12600 2228 12628
rect 2179 12597 2191 12600
rect 2133 12591 2191 12597
rect 2222 12588 2228 12600
rect 2280 12588 2286 12640
rect 4065 12631 4123 12637
rect 4065 12597 4077 12631
rect 4111 12628 4123 12631
rect 4154 12628 4160 12640
rect 4111 12600 4160 12628
rect 4111 12597 4123 12600
rect 4065 12591 4123 12597
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 5718 12628 5724 12640
rect 5679 12600 5724 12628
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 6748 12628 6776 12727
rect 7098 12724 7104 12736
rect 7156 12724 7162 12776
rect 7377 12767 7435 12773
rect 7377 12733 7389 12767
rect 7423 12764 7435 12767
rect 7834 12764 7840 12776
rect 7423 12736 7840 12764
rect 7423 12733 7435 12736
rect 7377 12727 7435 12733
rect 7834 12724 7840 12736
rect 7892 12764 7898 12776
rect 7944 12764 7972 12804
rect 9398 12792 9404 12804
rect 9456 12792 9462 12844
rect 7892 12736 7972 12764
rect 8113 12767 8171 12773
rect 7892 12724 7898 12736
rect 8113 12733 8125 12767
rect 8159 12764 8171 12767
rect 8478 12764 8484 12776
rect 8159 12736 8484 12764
rect 8159 12733 8171 12736
rect 8113 12727 8171 12733
rect 8478 12724 8484 12736
rect 8536 12724 8542 12776
rect 9766 12724 9772 12776
rect 9824 12764 9830 12776
rect 13354 12764 13360 12776
rect 9824 12736 13360 12764
rect 9824 12724 9830 12736
rect 13354 12724 13360 12736
rect 13412 12724 13418 12776
rect 14277 12767 14335 12773
rect 14277 12733 14289 12767
rect 14323 12764 14335 12767
rect 14918 12764 14924 12776
rect 14323 12736 14924 12764
rect 14323 12733 14335 12736
rect 14277 12727 14335 12733
rect 14918 12724 14924 12736
rect 14976 12724 14982 12776
rect 7190 12696 7196 12708
rect 7151 12668 7196 12696
rect 7190 12656 7196 12668
rect 7248 12656 7254 12708
rect 7282 12656 7288 12708
rect 7340 12696 7346 12708
rect 7926 12696 7932 12708
rect 7340 12668 7932 12696
rect 7340 12656 7346 12668
rect 7926 12656 7932 12668
rect 7984 12656 7990 12708
rect 8294 12696 8300 12708
rect 8255 12668 8300 12696
rect 8294 12656 8300 12668
rect 8352 12656 8358 12708
rect 14553 12699 14611 12705
rect 14553 12665 14565 12699
rect 14599 12696 14611 12699
rect 15010 12696 15016 12708
rect 14599 12668 15016 12696
rect 14599 12665 14611 12668
rect 14553 12659 14611 12665
rect 15010 12656 15016 12668
rect 15068 12656 15074 12708
rect 7742 12628 7748 12640
rect 6748 12600 7748 12628
rect 7742 12588 7748 12600
rect 7800 12588 7806 12640
rect 13722 12628 13728 12640
rect 13683 12600 13728 12628
rect 13722 12588 13728 12600
rect 13780 12628 13786 12640
rect 14369 12631 14427 12637
rect 14369 12628 14381 12631
rect 13780 12600 14381 12628
rect 13780 12588 13786 12600
rect 14369 12597 14381 12600
rect 14415 12597 14427 12631
rect 14369 12591 14427 12597
rect 1104 12538 16100 12560
rect 1104 12486 5980 12538
rect 6032 12486 6044 12538
rect 6096 12486 6108 12538
rect 6160 12486 6172 12538
rect 6224 12486 10979 12538
rect 11031 12486 11043 12538
rect 11095 12486 11107 12538
rect 11159 12486 11171 12538
rect 11223 12486 16100 12538
rect 1104 12464 16100 12486
rect 3878 12384 3884 12436
rect 3936 12424 3942 12436
rect 4893 12427 4951 12433
rect 4893 12424 4905 12427
rect 3936 12396 4905 12424
rect 3936 12384 3942 12396
rect 4893 12393 4905 12396
rect 4939 12393 4951 12427
rect 4893 12387 4951 12393
rect 4982 12384 4988 12436
rect 5040 12424 5046 12436
rect 5350 12424 5356 12436
rect 5040 12396 5356 12424
rect 5040 12384 5046 12396
rect 5350 12384 5356 12396
rect 5408 12424 5414 12436
rect 5408 12396 6224 12424
rect 5408 12384 5414 12396
rect 2222 12316 2228 12368
rect 2280 12316 2286 12368
rect 2866 12316 2872 12368
rect 2924 12356 2930 12368
rect 4154 12356 4160 12368
rect 2924 12328 3280 12356
rect 4115 12328 4160 12356
rect 2924 12316 2930 12328
rect 3252 12300 3280 12328
rect 4154 12316 4160 12328
rect 4212 12316 4218 12368
rect 4246 12316 4252 12368
rect 4304 12356 4310 12368
rect 6086 12356 6092 12368
rect 4304 12328 4349 12356
rect 6047 12328 6092 12356
rect 4304 12316 4310 12328
rect 6086 12316 6092 12328
rect 6144 12316 6150 12368
rect 3234 12248 3240 12300
rect 3292 12288 3298 12300
rect 3510 12288 3516 12300
rect 3292 12260 3337 12288
rect 3471 12260 3516 12288
rect 3292 12248 3298 12260
rect 3510 12248 3516 12260
rect 3568 12248 3574 12300
rect 3697 12291 3755 12297
rect 3697 12257 3709 12291
rect 3743 12288 3755 12291
rect 3878 12288 3884 12300
rect 3743 12260 3884 12288
rect 3743 12257 3755 12260
rect 3697 12251 3755 12257
rect 3878 12248 3884 12260
rect 3936 12248 3942 12300
rect 4065 12291 4123 12297
rect 4065 12257 4077 12291
rect 4111 12257 4123 12291
rect 4367 12291 4425 12297
rect 4367 12288 4379 12291
rect 4065 12251 4123 12257
rect 4356 12257 4379 12288
rect 4413 12257 4425 12291
rect 4614 12288 4620 12300
rect 4575 12260 4620 12288
rect 4356 12251 4425 12257
rect 1670 12180 1676 12232
rect 1728 12220 1734 12232
rect 2866 12220 2872 12232
rect 1728 12192 2872 12220
rect 1728 12180 1734 12192
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12220 3019 12223
rect 3605 12223 3663 12229
rect 3007 12192 3464 12220
rect 3007 12189 3019 12192
rect 2961 12183 3019 12189
rect 3436 12152 3464 12192
rect 3605 12189 3617 12223
rect 3651 12220 3663 12223
rect 4080 12220 4108 12251
rect 3651 12192 4108 12220
rect 3651 12189 3663 12192
rect 3605 12183 3663 12189
rect 3881 12155 3939 12161
rect 3881 12152 3893 12155
rect 3436 12124 3893 12152
rect 3881 12121 3893 12124
rect 3927 12121 3939 12155
rect 3881 12115 3939 12121
rect 4356 12096 4384 12251
rect 4614 12248 4620 12260
rect 4672 12288 4678 12300
rect 4982 12288 4988 12300
rect 4672 12260 4988 12288
rect 4672 12248 4678 12260
rect 4982 12248 4988 12260
rect 5040 12248 5046 12300
rect 5166 12288 5172 12300
rect 5127 12260 5172 12288
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 5445 12291 5503 12297
rect 5445 12257 5457 12291
rect 5491 12288 5503 12291
rect 5718 12288 5724 12300
rect 5491 12260 5724 12288
rect 5491 12257 5503 12260
rect 5445 12251 5503 12257
rect 5718 12248 5724 12260
rect 5776 12248 5782 12300
rect 5905 12291 5963 12297
rect 5905 12257 5917 12291
rect 5951 12257 5963 12291
rect 5905 12251 5963 12257
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12220 4951 12223
rect 5074 12220 5080 12232
rect 4939 12192 5080 12220
rect 4939 12189 4951 12192
rect 4893 12183 4951 12189
rect 1489 12087 1547 12093
rect 1489 12053 1501 12087
rect 1535 12084 1547 12087
rect 4338 12084 4344 12096
rect 1535 12056 4344 12084
rect 1535 12053 1547 12056
rect 1489 12047 1547 12053
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 4430 12044 4436 12096
rect 4488 12084 4494 12096
rect 4540 12084 4568 12183
rect 5074 12180 5080 12192
rect 5132 12220 5138 12232
rect 5251 12223 5309 12229
rect 5251 12220 5263 12223
rect 5132 12192 5263 12220
rect 5132 12180 5138 12192
rect 5251 12189 5263 12192
rect 5297 12189 5309 12223
rect 5251 12183 5309 12189
rect 5629 12223 5687 12229
rect 5629 12189 5641 12223
rect 5675 12220 5687 12223
rect 5810 12220 5816 12232
rect 5675 12192 5816 12220
rect 5675 12189 5687 12192
rect 5629 12183 5687 12189
rect 5810 12180 5816 12192
rect 5868 12180 5874 12232
rect 5353 12155 5411 12161
rect 5353 12121 5365 12155
rect 5399 12152 5411 12155
rect 5442 12152 5448 12164
rect 5399 12124 5448 12152
rect 5399 12121 5411 12124
rect 5353 12115 5411 12121
rect 5442 12112 5448 12124
rect 5500 12152 5506 12164
rect 5721 12155 5779 12161
rect 5721 12152 5733 12155
rect 5500 12124 5733 12152
rect 5500 12112 5506 12124
rect 5721 12121 5733 12124
rect 5767 12121 5779 12155
rect 5721 12115 5779 12121
rect 4706 12084 4712 12096
rect 4488 12056 4568 12084
rect 4667 12056 4712 12084
rect 4488 12044 4494 12056
rect 4706 12044 4712 12056
rect 4764 12084 4770 12096
rect 5920 12084 5948 12251
rect 5994 12248 6000 12300
rect 6052 12288 6058 12300
rect 6196 12288 6224 12396
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 8386 12424 8392 12436
rect 6972 12396 8392 12424
rect 6972 12384 6978 12396
rect 8386 12384 8392 12396
rect 8444 12384 8450 12436
rect 9766 12424 9772 12436
rect 9727 12396 9772 12424
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 11330 12384 11336 12436
rect 11388 12424 11394 12436
rect 11517 12427 11575 12433
rect 11517 12424 11529 12427
rect 11388 12396 11529 12424
rect 11388 12384 11394 12396
rect 11517 12393 11529 12396
rect 11563 12393 11575 12427
rect 11517 12387 11575 12393
rect 12713 12427 12771 12433
rect 12713 12393 12725 12427
rect 12759 12424 12771 12427
rect 12759 12396 13584 12424
rect 12759 12393 12771 12396
rect 12713 12387 12771 12393
rect 7377 12359 7435 12365
rect 6472 12328 7328 12356
rect 6472 12300 6500 12328
rect 6273 12291 6331 12297
rect 6273 12288 6285 12291
rect 6052 12260 6097 12288
rect 6196 12260 6285 12288
rect 6052 12248 6058 12260
rect 6273 12257 6285 12260
rect 6319 12257 6331 12291
rect 6454 12288 6460 12300
rect 6367 12260 6460 12288
rect 6273 12251 6331 12257
rect 6454 12248 6460 12260
rect 6512 12248 6518 12300
rect 6546 12248 6552 12300
rect 6604 12288 6610 12300
rect 6733 12291 6791 12297
rect 6604 12260 6649 12288
rect 6604 12248 6610 12260
rect 6733 12257 6745 12291
rect 6779 12288 6791 12291
rect 7006 12288 7012 12300
rect 6779 12260 7012 12288
rect 6779 12257 6791 12260
rect 6733 12251 6791 12257
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 7300 12297 7328 12328
rect 7377 12325 7389 12359
rect 7423 12356 7435 12359
rect 7650 12356 7656 12368
rect 7423 12328 7656 12356
rect 7423 12325 7435 12328
rect 7377 12319 7435 12325
rect 7650 12316 7656 12328
rect 7708 12356 7714 12368
rect 8110 12356 8116 12368
rect 7708 12328 8116 12356
rect 7708 12316 7714 12328
rect 7760 12297 7788 12328
rect 8110 12316 8116 12328
rect 8168 12316 8174 12368
rect 8294 12356 8300 12368
rect 8220 12328 8300 12356
rect 7285 12291 7343 12297
rect 7285 12257 7297 12291
rect 7331 12257 7343 12291
rect 7285 12251 7343 12257
rect 7745 12291 7803 12297
rect 7745 12257 7757 12291
rect 7791 12257 7803 12291
rect 8018 12288 8024 12300
rect 7979 12260 8024 12288
rect 7745 12251 7803 12257
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 8220 12297 8248 12328
rect 8294 12316 8300 12328
rect 8352 12356 8358 12368
rect 9858 12356 9864 12368
rect 8352 12328 9076 12356
rect 8352 12316 8358 12328
rect 9048 12300 9076 12328
rect 9462 12328 9720 12356
rect 9819 12328 9864 12356
rect 8205 12291 8263 12297
rect 8205 12257 8217 12291
rect 8251 12257 8263 12291
rect 8478 12288 8484 12300
rect 8391 12260 8484 12288
rect 8205 12251 8263 12257
rect 8478 12248 8484 12260
rect 8536 12288 8542 12300
rect 8536 12260 8984 12288
rect 8536 12248 8542 12260
rect 6914 12220 6920 12232
rect 6875 12192 6920 12220
rect 6914 12180 6920 12192
rect 6972 12180 6978 12232
rect 7837 12223 7895 12229
rect 7837 12189 7849 12223
rect 7883 12220 7895 12223
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 7883 12192 8401 12220
rect 7883 12189 7895 12192
rect 7837 12183 7895 12189
rect 8389 12189 8401 12192
rect 8435 12189 8447 12223
rect 8389 12183 8447 12189
rect 6270 12112 6276 12164
rect 6328 12152 6334 12164
rect 7852 12152 7880 12183
rect 6328 12124 7880 12152
rect 6328 12112 6334 12124
rect 7926 12112 7932 12164
rect 7984 12152 7990 12164
rect 8956 12152 8984 12260
rect 9030 12248 9036 12300
rect 9088 12288 9094 12300
rect 9125 12291 9183 12297
rect 9125 12288 9137 12291
rect 9088 12260 9137 12288
rect 9088 12248 9094 12260
rect 9125 12257 9137 12260
rect 9171 12257 9183 12291
rect 9125 12251 9183 12257
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 9462 12288 9490 12328
rect 9582 12288 9588 12300
rect 9364 12260 9490 12288
rect 9543 12260 9588 12288
rect 9364 12248 9370 12260
rect 9582 12248 9588 12260
rect 9640 12248 9646 12300
rect 9692 12288 9720 12328
rect 9858 12316 9864 12328
rect 9916 12316 9922 12368
rect 10336 12328 12204 12356
rect 10336 12297 10364 12328
rect 12176 12300 12204 12328
rect 12434 12316 12440 12368
rect 12492 12356 12498 12368
rect 12957 12359 13015 12365
rect 12957 12356 12969 12359
rect 12492 12328 12969 12356
rect 12492 12316 12498 12328
rect 12957 12325 12969 12328
rect 13003 12325 13015 12359
rect 13170 12356 13176 12368
rect 13131 12328 13176 12356
rect 12957 12319 13015 12325
rect 13170 12316 13176 12328
rect 13228 12316 13234 12368
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 9692 12260 10057 12288
rect 10045 12257 10057 12260
rect 10091 12257 10103 12291
rect 10045 12251 10103 12257
rect 10321 12291 10379 12297
rect 10321 12257 10333 12291
rect 10367 12257 10379 12291
rect 10321 12251 10379 12257
rect 9214 12180 9220 12232
rect 9272 12220 9278 12232
rect 9766 12220 9772 12232
rect 9272 12192 9772 12220
rect 9272 12180 9278 12192
rect 9766 12180 9772 12192
rect 9824 12180 9830 12232
rect 10060 12220 10088 12251
rect 11054 12248 11060 12300
rect 11112 12288 11118 12300
rect 11425 12291 11483 12297
rect 11425 12288 11437 12291
rect 11112 12260 11437 12288
rect 11112 12248 11118 12260
rect 11425 12257 11437 12260
rect 11471 12257 11483 12291
rect 11425 12251 11483 12257
rect 12158 12248 12164 12300
rect 12216 12288 12222 12300
rect 12253 12291 12311 12297
rect 12253 12288 12265 12291
rect 12216 12260 12265 12288
rect 12216 12248 12222 12260
rect 12253 12257 12265 12260
rect 12299 12257 12311 12291
rect 12253 12251 12311 12257
rect 12529 12291 12587 12297
rect 12529 12257 12541 12291
rect 12575 12288 12587 12291
rect 13265 12291 13323 12297
rect 12575 12260 13032 12288
rect 12575 12257 12587 12260
rect 12529 12251 12587 12257
rect 13004 12232 13032 12260
rect 13265 12257 13277 12291
rect 13311 12288 13323 12291
rect 13354 12288 13360 12300
rect 13311 12260 13360 12288
rect 13311 12257 13323 12260
rect 13265 12251 13323 12257
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 10060 12192 12388 12220
rect 12360 12164 12388 12192
rect 12986 12180 12992 12232
rect 13044 12180 13050 12232
rect 13556 12220 13584 12396
rect 13722 12356 13728 12368
rect 13683 12328 13728 12356
rect 13722 12316 13728 12328
rect 13780 12316 13786 12368
rect 13832 12328 14596 12356
rect 13832 12297 13860 12328
rect 13817 12291 13875 12297
rect 13817 12257 13829 12291
rect 13863 12257 13875 12291
rect 13817 12251 13875 12257
rect 14369 12291 14427 12297
rect 14369 12257 14381 12291
rect 14415 12257 14427 12291
rect 14568 12288 14596 12328
rect 14918 12297 14924 12300
rect 14897 12291 14924 12297
rect 14897 12288 14909 12291
rect 14568 12260 14909 12288
rect 14369 12251 14427 12257
rect 14897 12257 14909 12260
rect 14897 12251 14924 12257
rect 14384 12220 14412 12251
rect 14918 12248 14924 12251
rect 14976 12248 14982 12300
rect 15010 12248 15016 12300
rect 15068 12288 15074 12300
rect 15068 12260 15113 12288
rect 15068 12248 15074 12260
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 13556 12192 15393 12220
rect 15381 12189 15393 12192
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 9306 12152 9312 12164
rect 7984 12124 8892 12152
rect 8956 12124 9312 12152
rect 7984 12112 7990 12124
rect 4764 12056 5948 12084
rect 7561 12087 7619 12093
rect 4764 12044 4770 12056
rect 7561 12053 7573 12087
rect 7607 12084 7619 12087
rect 8294 12084 8300 12096
rect 7607 12056 8300 12084
rect 7607 12053 7619 12056
rect 7561 12047 7619 12053
rect 8294 12044 8300 12056
rect 8352 12044 8358 12096
rect 8864 12084 8892 12124
rect 9306 12112 9312 12124
rect 9364 12112 9370 12164
rect 9401 12155 9459 12161
rect 9401 12121 9413 12155
rect 9447 12121 9459 12155
rect 9401 12115 9459 12121
rect 8938 12084 8944 12096
rect 8851 12056 8944 12084
rect 8938 12044 8944 12056
rect 8996 12084 9002 12096
rect 9416 12084 9444 12115
rect 9490 12112 9496 12164
rect 9548 12152 9554 12164
rect 9548 12124 9593 12152
rect 9548 12112 9554 12124
rect 9858 12112 9864 12164
rect 9916 12152 9922 12164
rect 10137 12155 10195 12161
rect 10137 12152 10149 12155
rect 9916 12124 10149 12152
rect 9916 12112 9922 12124
rect 10137 12121 10149 12124
rect 10183 12121 10195 12155
rect 10137 12115 10195 12121
rect 10226 12112 10232 12164
rect 10284 12152 10290 12164
rect 12342 12152 12348 12164
rect 10284 12124 10329 12152
rect 12303 12124 12348 12152
rect 10284 12112 10290 12124
rect 12342 12112 12348 12124
rect 12400 12112 12406 12164
rect 12434 12112 12440 12164
rect 12492 12152 12498 12164
rect 12492 12124 12537 12152
rect 12636 12124 13032 12152
rect 12492 12112 12498 12124
rect 12250 12084 12256 12096
rect 8996 12056 12256 12084
rect 8996 12044 9002 12056
rect 12250 12044 12256 12056
rect 12308 12084 12314 12096
rect 12636 12084 12664 12124
rect 12308 12056 12664 12084
rect 12308 12044 12314 12056
rect 12710 12044 12716 12096
rect 12768 12084 12774 12096
rect 13004 12093 13032 12124
rect 12805 12087 12863 12093
rect 12805 12084 12817 12087
rect 12768 12056 12817 12084
rect 12768 12044 12774 12056
rect 12805 12053 12817 12056
rect 12851 12053 12863 12087
rect 12805 12047 12863 12053
rect 12989 12087 13047 12093
rect 12989 12053 13001 12087
rect 13035 12053 13047 12087
rect 12989 12047 13047 12053
rect 14921 12087 14979 12093
rect 14921 12053 14933 12087
rect 14967 12084 14979 12087
rect 15010 12084 15016 12096
rect 14967 12056 15016 12084
rect 14967 12053 14979 12056
rect 14921 12047 14979 12053
rect 15010 12044 15016 12056
rect 15068 12044 15074 12096
rect 1104 11994 16100 12016
rect 1104 11942 3481 11994
rect 3533 11942 3545 11994
rect 3597 11942 3609 11994
rect 3661 11942 3673 11994
rect 3725 11942 8480 11994
rect 8532 11942 8544 11994
rect 8596 11942 8608 11994
rect 8660 11942 8672 11994
rect 8724 11942 13478 11994
rect 13530 11942 13542 11994
rect 13594 11942 13606 11994
rect 13658 11942 13670 11994
rect 13722 11942 16100 11994
rect 1104 11920 16100 11942
rect 6454 11840 6460 11892
rect 6512 11880 6518 11892
rect 6549 11883 6607 11889
rect 6549 11880 6561 11883
rect 6512 11852 6561 11880
rect 6512 11840 6518 11852
rect 6549 11849 6561 11852
rect 6595 11849 6607 11883
rect 6549 11843 6607 11849
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 9493 11883 9551 11889
rect 8352 11852 9444 11880
rect 8352 11840 8358 11852
rect 2774 11772 2780 11824
rect 2832 11812 2838 11824
rect 4062 11812 4068 11824
rect 2832 11784 4068 11812
rect 2832 11772 2838 11784
rect 4062 11772 4068 11784
rect 4120 11812 4126 11824
rect 4430 11812 4436 11824
rect 4120 11784 4436 11812
rect 4120 11772 4126 11784
rect 4430 11772 4436 11784
rect 4488 11772 4494 11824
rect 8849 11815 8907 11821
rect 8849 11781 8861 11815
rect 8895 11812 8907 11815
rect 8938 11812 8944 11824
rect 8895 11784 8944 11812
rect 8895 11781 8907 11784
rect 8849 11775 8907 11781
rect 8938 11772 8944 11784
rect 8996 11772 9002 11824
rect 9416 11812 9444 11852
rect 9493 11849 9505 11883
rect 9539 11880 9551 11883
rect 9582 11880 9588 11892
rect 9539 11852 9588 11880
rect 9539 11849 9551 11852
rect 9493 11843 9551 11849
rect 9582 11840 9588 11852
rect 9640 11880 9646 11892
rect 9858 11880 9864 11892
rect 9640 11852 9864 11880
rect 9640 11840 9646 11852
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 10505 11883 10563 11889
rect 10505 11849 10517 11883
rect 10551 11880 10563 11883
rect 11054 11880 11060 11892
rect 10551 11852 11060 11880
rect 10551 11849 10563 11852
rect 10505 11843 10563 11849
rect 11054 11840 11060 11852
rect 11112 11840 11118 11892
rect 10410 11812 10416 11824
rect 9140 11784 9352 11812
rect 9416 11784 9674 11812
rect 9140 11744 9168 11784
rect 8772 11716 9168 11744
rect 8772 11688 8800 11716
rect 4338 11636 4344 11688
rect 4396 11676 4402 11688
rect 5350 11676 5356 11688
rect 4396 11648 5356 11676
rect 4396 11636 4402 11648
rect 5350 11636 5356 11648
rect 5408 11676 5414 11688
rect 5994 11676 6000 11688
rect 5408 11648 6000 11676
rect 5408 11636 5414 11648
rect 5994 11636 6000 11648
rect 6052 11676 6058 11688
rect 6089 11679 6147 11685
rect 6089 11676 6101 11679
rect 6052 11648 6101 11676
rect 6052 11636 6058 11648
rect 6089 11645 6101 11648
rect 6135 11645 6147 11679
rect 8754 11676 8760 11688
rect 8715 11648 8760 11676
rect 6089 11639 6147 11645
rect 8754 11636 8760 11648
rect 8812 11636 8818 11688
rect 8938 11676 8944 11688
rect 8899 11648 8944 11676
rect 8938 11636 8944 11648
rect 8996 11636 9002 11688
rect 9033 11679 9091 11685
rect 9033 11645 9045 11679
rect 9079 11645 9091 11679
rect 9033 11639 9091 11645
rect 6730 11608 6736 11620
rect 6691 11580 6736 11608
rect 6730 11568 6736 11580
rect 6788 11568 6794 11620
rect 6917 11611 6975 11617
rect 6917 11577 6929 11611
rect 6963 11577 6975 11611
rect 9048 11608 9076 11639
rect 9122 11636 9128 11688
rect 9180 11676 9186 11688
rect 9324 11685 9352 11784
rect 9646 11744 9674 11784
rect 9876 11784 10416 11812
rect 9876 11744 9904 11784
rect 10410 11772 10416 11784
rect 10468 11772 10474 11824
rect 10594 11744 10600 11756
rect 9646 11716 9904 11744
rect 9968 11716 10600 11744
rect 9214 11679 9272 11685
rect 9214 11676 9226 11679
rect 9180 11648 9226 11676
rect 9180 11636 9186 11648
rect 9214 11645 9226 11648
rect 9260 11645 9272 11679
rect 9214 11639 9272 11645
rect 9309 11679 9367 11685
rect 9309 11645 9321 11679
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 9493 11679 9551 11685
rect 9493 11645 9505 11679
rect 9539 11676 9551 11679
rect 9582 11676 9588 11688
rect 9539 11648 9588 11676
rect 9539 11645 9551 11648
rect 9493 11639 9551 11645
rect 9582 11636 9588 11648
rect 9640 11636 9646 11688
rect 9674 11636 9680 11688
rect 9732 11676 9738 11688
rect 9968 11685 9996 11716
rect 10594 11704 10600 11716
rect 10652 11744 10658 11756
rect 10689 11747 10747 11753
rect 10689 11744 10701 11747
rect 10652 11716 10701 11744
rect 10652 11704 10658 11716
rect 10689 11713 10701 11716
rect 10735 11744 10747 11747
rect 12161 11747 12219 11753
rect 12161 11744 12173 11747
rect 10735 11716 12173 11744
rect 10735 11713 10747 11716
rect 10689 11707 10747 11713
rect 12161 11713 12173 11716
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 12250 11704 12256 11756
rect 12308 11744 12314 11756
rect 12345 11747 12403 11753
rect 12345 11744 12357 11747
rect 12308 11716 12357 11744
rect 12308 11704 12314 11716
rect 12345 11713 12357 11716
rect 12391 11713 12403 11747
rect 12345 11707 12403 11713
rect 9953 11679 10011 11685
rect 9953 11676 9965 11679
rect 9732 11648 9965 11676
rect 9732 11636 9738 11648
rect 9953 11645 9965 11648
rect 9999 11645 10011 11679
rect 10502 11676 10508 11688
rect 10463 11648 10508 11676
rect 9953 11639 10011 11645
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 10870 11636 10876 11688
rect 10928 11676 10934 11688
rect 11057 11679 11115 11685
rect 11057 11676 11069 11679
rect 10928 11648 11069 11676
rect 10928 11636 10934 11648
rect 11057 11645 11069 11648
rect 11103 11645 11115 11679
rect 11057 11639 11115 11645
rect 12434 11636 12440 11688
rect 12492 11676 12498 11688
rect 12529 11679 12587 11685
rect 12529 11676 12541 11679
rect 12492 11648 12541 11676
rect 12492 11636 12498 11648
rect 12529 11645 12541 11648
rect 12575 11645 12587 11679
rect 12529 11639 12587 11645
rect 12621 11679 12679 11685
rect 12621 11645 12633 11679
rect 12667 11676 12679 11679
rect 13170 11676 13176 11688
rect 12667 11648 13176 11676
rect 12667 11645 12679 11648
rect 12621 11639 12679 11645
rect 9048 11580 9720 11608
rect 6917 11571 6975 11577
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 6181 11543 6239 11549
rect 6181 11540 6193 11543
rect 5500 11512 6193 11540
rect 5500 11500 5506 11512
rect 6181 11509 6193 11512
rect 6227 11540 6239 11543
rect 6270 11540 6276 11552
rect 6227 11512 6276 11540
rect 6227 11509 6239 11512
rect 6181 11503 6239 11509
rect 6270 11500 6276 11512
rect 6328 11540 6334 11552
rect 6932 11540 6960 11571
rect 8110 11540 8116 11552
rect 6328 11512 8116 11540
rect 6328 11500 6334 11512
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 8573 11543 8631 11549
rect 8573 11540 8585 11543
rect 8352 11512 8585 11540
rect 8352 11500 8358 11512
rect 8573 11509 8585 11512
rect 8619 11509 8631 11543
rect 8573 11503 8631 11509
rect 9306 11500 9312 11552
rect 9364 11540 9370 11552
rect 9582 11540 9588 11552
rect 9364 11512 9588 11540
rect 9364 11500 9370 11512
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 9692 11549 9720 11580
rect 11882 11568 11888 11620
rect 11940 11608 11946 11620
rect 12342 11608 12348 11620
rect 11940 11580 12348 11608
rect 11940 11568 11946 11580
rect 12342 11568 12348 11580
rect 12400 11608 12406 11620
rect 12636 11608 12664 11639
rect 13170 11636 13176 11648
rect 13228 11636 13234 11688
rect 12400 11580 12664 11608
rect 12400 11568 12406 11580
rect 9677 11543 9735 11549
rect 9677 11509 9689 11543
rect 9723 11509 9735 11543
rect 9677 11503 9735 11509
rect 1104 11450 16100 11472
rect 1104 11398 5980 11450
rect 6032 11398 6044 11450
rect 6096 11398 6108 11450
rect 6160 11398 6172 11450
rect 6224 11398 10979 11450
rect 11031 11398 11043 11450
rect 11095 11398 11107 11450
rect 11159 11398 11171 11450
rect 11223 11398 16100 11450
rect 1104 11376 16100 11398
rect 5350 11336 5356 11348
rect 5311 11308 5356 11336
rect 5350 11296 5356 11308
rect 5408 11336 5414 11348
rect 7190 11336 7196 11348
rect 5408 11308 7196 11336
rect 5408 11296 5414 11308
rect 2130 11228 2136 11280
rect 2188 11228 2194 11280
rect 6914 11268 6920 11280
rect 4264 11240 6920 11268
rect 4264 11209 4292 11240
rect 6914 11228 6920 11240
rect 6972 11228 6978 11280
rect 4249 11203 4307 11209
rect 4249 11169 4261 11203
rect 4295 11169 4307 11203
rect 4430 11200 4436 11212
rect 4391 11172 4436 11200
rect 4249 11163 4307 11169
rect 4430 11160 4436 11172
rect 4488 11160 4494 11212
rect 5074 11160 5080 11212
rect 5132 11200 5138 11212
rect 5132 11172 5580 11200
rect 5132 11160 5138 11172
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 1670 11132 1676 11144
rect 1443 11104 1676 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 1670 11092 1676 11104
rect 1728 11092 1734 11144
rect 3878 11092 3884 11144
rect 3936 11132 3942 11144
rect 4706 11132 4712 11144
rect 3936 11104 4712 11132
rect 3936 11092 3942 11104
rect 4706 11092 4712 11104
rect 4764 11132 4770 11144
rect 5552 11141 5580 11172
rect 6730 11160 6736 11212
rect 6788 11200 6794 11212
rect 7024 11209 7052 11308
rect 7190 11296 7196 11308
rect 7248 11296 7254 11348
rect 7558 11336 7564 11348
rect 7519 11308 7564 11336
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 8110 11296 8116 11348
rect 8168 11336 8174 11348
rect 9398 11336 9404 11348
rect 8168 11308 9404 11336
rect 8168 11296 8174 11308
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 10965 11339 11023 11345
rect 10965 11336 10977 11339
rect 10928 11308 10977 11336
rect 10928 11296 10934 11308
rect 10965 11305 10977 11308
rect 11011 11305 11023 11339
rect 10965 11299 11023 11305
rect 7300 11240 9812 11268
rect 6825 11203 6883 11209
rect 6825 11200 6837 11203
rect 6788 11172 6837 11200
rect 6788 11160 6794 11172
rect 6825 11169 6837 11172
rect 6871 11169 6883 11203
rect 6825 11163 6883 11169
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11169 7067 11203
rect 7009 11163 7067 11169
rect 5445 11135 5503 11141
rect 5445 11132 5457 11135
rect 4764 11104 5457 11132
rect 4764 11092 4770 11104
rect 5445 11101 5457 11104
rect 5491 11101 5503 11135
rect 5445 11095 5503 11101
rect 5537 11135 5595 11141
rect 5537 11101 5549 11135
rect 5583 11101 5595 11135
rect 6840 11132 6868 11163
rect 7098 11160 7104 11212
rect 7156 11200 7162 11212
rect 7300 11209 7328 11240
rect 9784 11212 9812 11240
rect 15010 11228 15016 11280
rect 15068 11268 15074 11280
rect 15289 11271 15347 11277
rect 15289 11268 15301 11271
rect 15068 11240 15301 11268
rect 15068 11228 15074 11240
rect 15289 11237 15301 11240
rect 15335 11237 15347 11271
rect 15289 11231 15347 11237
rect 7193 11203 7251 11209
rect 7193 11200 7205 11203
rect 7156 11172 7205 11200
rect 7156 11160 7162 11172
rect 7193 11169 7205 11172
rect 7239 11169 7251 11203
rect 7193 11163 7251 11169
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 7653 11203 7711 11209
rect 7653 11169 7665 11203
rect 7699 11200 7711 11203
rect 7834 11200 7840 11212
rect 7699 11172 7840 11200
rect 7699 11169 7711 11172
rect 7653 11163 7711 11169
rect 7834 11160 7840 11172
rect 7892 11160 7898 11212
rect 8846 11160 8852 11212
rect 8904 11200 8910 11212
rect 9309 11203 9367 11209
rect 9309 11200 9321 11203
rect 8904 11172 9321 11200
rect 8904 11160 8910 11172
rect 9309 11169 9321 11172
rect 9355 11169 9367 11203
rect 9582 11200 9588 11212
rect 9543 11172 9588 11200
rect 9309 11163 9367 11169
rect 9582 11160 9588 11172
rect 9640 11160 9646 11212
rect 9766 11200 9772 11212
rect 9727 11172 9772 11200
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 10870 11200 10876 11212
rect 10831 11172 10876 11200
rect 10870 11160 10876 11172
rect 10928 11160 10934 11212
rect 7745 11135 7803 11141
rect 7745 11132 7757 11135
rect 6840 11104 7757 11132
rect 5537 11095 5595 11101
rect 7745 11101 7757 11104
rect 7791 11132 7803 11135
rect 8938 11132 8944 11144
rect 7791 11104 8944 11132
rect 7791 11101 7803 11104
rect 7745 11095 7803 11101
rect 8938 11092 8944 11104
rect 8996 11132 9002 11144
rect 9493 11135 9551 11141
rect 9493 11132 9505 11135
rect 8996 11104 9505 11132
rect 8996 11092 9002 11104
rect 9493 11101 9505 11104
rect 9539 11101 9551 11135
rect 9493 11095 9551 11101
rect 3786 11024 3792 11076
rect 3844 11064 3850 11076
rect 3844 11036 4200 11064
rect 3844 11024 3850 11036
rect 1660 10999 1718 11005
rect 1660 10965 1672 10999
rect 1706 10996 1718 10999
rect 2222 10996 2228 11008
rect 1706 10968 2228 10996
rect 1706 10965 1718 10968
rect 1660 10959 1718 10965
rect 2222 10956 2228 10968
rect 2280 10956 2286 11008
rect 3145 10999 3203 11005
rect 3145 10965 3157 10999
rect 3191 10996 3203 10999
rect 4062 10996 4068 11008
rect 3191 10968 4068 10996
rect 3191 10965 3203 10968
rect 3145 10959 3203 10965
rect 4062 10956 4068 10968
rect 4120 10956 4126 11008
rect 4172 10996 4200 11036
rect 4338 11024 4344 11076
rect 4396 11064 4402 11076
rect 7101 11067 7159 11073
rect 7101 11064 7113 11067
rect 4396 11036 7113 11064
rect 4396 11024 4402 11036
rect 7101 11033 7113 11036
rect 7147 11064 7159 11067
rect 8846 11064 8852 11076
rect 7147 11036 8852 11064
rect 7147 11033 7159 11036
rect 7101 11027 7159 11033
rect 8846 11024 8852 11036
rect 8904 11024 8910 11076
rect 9122 11024 9128 11076
rect 9180 11064 9186 11076
rect 9401 11067 9459 11073
rect 9180 11036 9225 11064
rect 9180 11024 9186 11036
rect 9401 11033 9413 11067
rect 9447 11064 9459 11067
rect 9858 11064 9864 11076
rect 9447 11036 9864 11064
rect 9447 11033 9459 11036
rect 9401 11027 9459 11033
rect 9858 11024 9864 11036
rect 9916 11024 9922 11076
rect 15102 11064 15108 11076
rect 15063 11036 15108 11064
rect 15102 11024 15108 11036
rect 15160 11024 15166 11076
rect 4249 10999 4307 11005
rect 4249 10996 4261 10999
rect 4172 10968 4261 10996
rect 4249 10965 4261 10968
rect 4295 10965 4307 10999
rect 4249 10959 4307 10965
rect 4617 10999 4675 11005
rect 4617 10965 4629 10999
rect 4663 10996 4675 10999
rect 4706 10996 4712 11008
rect 4663 10968 4712 10996
rect 4663 10965 4675 10968
rect 4617 10959 4675 10965
rect 4706 10956 4712 10968
rect 4764 10956 4770 11008
rect 4985 10999 5043 11005
rect 4985 10965 4997 10999
rect 5031 10996 5043 10999
rect 5074 10996 5080 11008
rect 5031 10968 5080 10996
rect 5031 10965 5043 10968
rect 4985 10959 5043 10965
rect 5074 10956 5080 10968
rect 5132 10956 5138 11008
rect 7006 10956 7012 11008
rect 7064 10996 7070 11008
rect 9214 10996 9220 11008
rect 7064 10968 9220 10996
rect 7064 10956 7070 10968
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 9306 10956 9312 11008
rect 9364 10996 9370 11008
rect 12986 10996 12992 11008
rect 9364 10968 12992 10996
rect 9364 10956 9370 10968
rect 12986 10956 12992 10968
rect 13044 10956 13050 11008
rect 1104 10906 16100 10928
rect 1104 10854 3481 10906
rect 3533 10854 3545 10906
rect 3597 10854 3609 10906
rect 3661 10854 3673 10906
rect 3725 10854 8480 10906
rect 8532 10854 8544 10906
rect 8596 10854 8608 10906
rect 8660 10854 8672 10906
rect 8724 10854 13478 10906
rect 13530 10854 13542 10906
rect 13594 10854 13606 10906
rect 13658 10854 13670 10906
rect 13722 10854 16100 10906
rect 1104 10832 16100 10854
rect 2130 10792 2136 10804
rect 2091 10764 2136 10792
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 2222 10752 2228 10804
rect 2280 10792 2286 10804
rect 2777 10795 2835 10801
rect 2777 10792 2789 10795
rect 2280 10764 2789 10792
rect 2280 10752 2286 10764
rect 2777 10761 2789 10764
rect 2823 10761 2835 10795
rect 2777 10755 2835 10761
rect 2869 10795 2927 10801
rect 2869 10761 2881 10795
rect 2915 10792 2927 10795
rect 2958 10792 2964 10804
rect 2915 10764 2964 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 2958 10752 2964 10764
rect 3016 10792 3022 10804
rect 4154 10792 4160 10804
rect 3016 10764 4160 10792
rect 3016 10752 3022 10764
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 4614 10752 4620 10804
rect 4672 10792 4678 10804
rect 4672 10764 4936 10792
rect 4672 10752 4678 10764
rect 3053 10727 3111 10733
rect 3053 10724 3065 10727
rect 2746 10696 3065 10724
rect 2746 10665 2774 10696
rect 3053 10693 3065 10696
rect 3099 10693 3111 10727
rect 3053 10687 3111 10693
rect 3786 10684 3792 10736
rect 3844 10724 3850 10736
rect 3844 10696 4844 10724
rect 3844 10684 3850 10696
rect 2731 10659 2789 10665
rect 2731 10625 2743 10659
rect 2777 10625 2789 10659
rect 4525 10659 4583 10665
rect 4525 10656 4537 10659
rect 2731 10619 2789 10625
rect 4356 10628 4537 10656
rect 1946 10588 1952 10600
rect 1907 10560 1952 10588
rect 1946 10548 1952 10560
rect 2004 10548 2010 10600
rect 2961 10591 3019 10597
rect 2961 10557 2973 10591
rect 3007 10588 3019 10591
rect 3050 10588 3056 10600
rect 3007 10560 3056 10588
rect 3007 10557 3019 10560
rect 2961 10551 3019 10557
rect 3050 10548 3056 10560
rect 3108 10548 3114 10600
rect 3234 10588 3240 10600
rect 3195 10560 3240 10588
rect 3234 10548 3240 10560
rect 3292 10548 3298 10600
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10557 3387 10591
rect 3329 10551 3387 10557
rect 2593 10523 2651 10529
rect 2593 10489 2605 10523
rect 2639 10520 2651 10523
rect 2774 10520 2780 10532
rect 2639 10492 2780 10520
rect 2639 10489 2651 10492
rect 2593 10483 2651 10489
rect 2774 10480 2780 10492
rect 2832 10480 2838 10532
rect 3344 10520 3372 10551
rect 3418 10548 3424 10600
rect 3476 10588 3482 10600
rect 3697 10591 3755 10597
rect 3697 10588 3709 10591
rect 3476 10560 3709 10588
rect 3476 10548 3482 10560
rect 3697 10557 3709 10560
rect 3743 10588 3755 10591
rect 3786 10588 3792 10600
rect 3743 10560 3792 10588
rect 3743 10557 3755 10560
rect 3697 10551 3755 10557
rect 3786 10548 3792 10560
rect 3844 10548 3850 10600
rect 3878 10548 3884 10600
rect 3936 10597 3942 10600
rect 3936 10591 3985 10597
rect 3936 10557 3939 10591
rect 3973 10557 3985 10591
rect 3936 10551 3985 10557
rect 3936 10548 3942 10551
rect 4062 10548 4068 10600
rect 4120 10588 4126 10600
rect 4356 10597 4384 10628
rect 4525 10625 4537 10628
rect 4571 10656 4583 10659
rect 4614 10656 4620 10668
rect 4571 10628 4620 10656
rect 4571 10625 4583 10628
rect 4525 10619 4583 10625
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 4341 10591 4399 10597
rect 4120 10560 4165 10588
rect 4120 10548 4126 10560
rect 4341 10557 4353 10591
rect 4387 10557 4399 10591
rect 4341 10551 4399 10557
rect 4430 10548 4436 10600
rect 4488 10588 4494 10600
rect 4816 10597 4844 10696
rect 4908 10656 4936 10764
rect 4982 10752 4988 10804
rect 5040 10792 5046 10804
rect 8110 10792 8116 10804
rect 5040 10764 5085 10792
rect 8071 10764 8116 10792
rect 5040 10752 5046 10764
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 8665 10795 8723 10801
rect 8665 10761 8677 10795
rect 8711 10792 8723 10795
rect 9493 10795 9551 10801
rect 8711 10764 9444 10792
rect 8711 10761 8723 10764
rect 8665 10755 8723 10761
rect 7098 10684 7104 10736
rect 7156 10724 7162 10736
rect 8205 10727 8263 10733
rect 8205 10724 8217 10727
rect 7156 10696 8217 10724
rect 7156 10684 7162 10696
rect 8205 10693 8217 10696
rect 8251 10693 8263 10727
rect 8205 10687 8263 10693
rect 9125 10727 9183 10733
rect 9125 10693 9137 10727
rect 9171 10724 9183 10727
rect 9416 10724 9444 10764
rect 9493 10761 9505 10795
rect 9539 10792 9551 10795
rect 9582 10792 9588 10804
rect 9539 10764 9588 10792
rect 9539 10761 9551 10764
rect 9493 10755 9551 10761
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 9766 10752 9772 10804
rect 9824 10792 9830 10804
rect 9824 10764 13308 10792
rect 9824 10752 9830 10764
rect 9784 10724 9812 10752
rect 9171 10696 9352 10724
rect 9416 10696 9812 10724
rect 9171 10693 9183 10696
rect 9125 10687 9183 10693
rect 8996 10659 9054 10665
rect 4908 10628 5396 10656
rect 4709 10591 4767 10597
rect 4488 10560 4533 10588
rect 4488 10548 4494 10560
rect 4709 10557 4721 10591
rect 4755 10557 4767 10591
rect 4709 10551 4767 10557
rect 4801 10591 4859 10597
rect 4801 10557 4813 10591
rect 4847 10557 4859 10591
rect 5074 10588 5080 10600
rect 5035 10560 5080 10588
rect 4801 10551 4859 10557
rect 3605 10523 3663 10529
rect 3605 10520 3617 10523
rect 3344 10492 3617 10520
rect 3605 10489 3617 10492
rect 3651 10489 3663 10523
rect 3605 10483 3663 10489
rect 4157 10523 4215 10529
rect 4157 10489 4169 10523
rect 4203 10520 4215 10523
rect 4448 10520 4476 10548
rect 4203 10492 4476 10520
rect 4203 10489 4215 10492
rect 4157 10483 4215 10489
rect 3620 10452 3648 10483
rect 3789 10455 3847 10461
rect 3789 10452 3801 10455
rect 3620 10424 3801 10452
rect 3789 10421 3801 10424
rect 3835 10452 3847 10455
rect 4724 10452 4752 10551
rect 5074 10548 5080 10560
rect 5132 10548 5138 10600
rect 5258 10588 5264 10600
rect 5219 10560 5264 10588
rect 5258 10548 5264 10560
rect 5316 10548 5322 10600
rect 5368 10597 5396 10628
rect 8996 10625 9008 10659
rect 9042 10656 9054 10659
rect 9214 10656 9220 10668
rect 9042 10625 9076 10656
rect 9175 10628 9220 10656
rect 8996 10619 9076 10625
rect 5353 10591 5411 10597
rect 5353 10557 5365 10591
rect 5399 10557 5411 10591
rect 5353 10551 5411 10557
rect 5442 10548 5448 10600
rect 5500 10588 5506 10600
rect 5500 10560 5545 10588
rect 5500 10548 5506 10560
rect 7834 10548 7840 10600
rect 7892 10588 7898 10600
rect 7929 10591 7987 10597
rect 7929 10588 7941 10591
rect 7892 10560 7941 10588
rect 7892 10548 7898 10560
rect 7929 10557 7941 10560
rect 7975 10557 7987 10591
rect 7929 10551 7987 10557
rect 8297 10591 8355 10597
rect 8297 10557 8309 10591
rect 8343 10557 8355 10591
rect 8297 10551 8355 10557
rect 8312 10520 8340 10551
rect 8386 10548 8392 10600
rect 8444 10588 8450 10600
rect 9048 10588 9076 10619
rect 9214 10616 9220 10628
rect 9272 10616 9278 10668
rect 9324 10656 9352 10696
rect 9858 10684 9864 10736
rect 9916 10724 9922 10736
rect 10965 10727 11023 10733
rect 9916 10696 10916 10724
rect 9916 10684 9922 10696
rect 9398 10656 9404 10668
rect 9324 10628 9404 10656
rect 9398 10616 9404 10628
rect 9456 10616 9462 10668
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 9968 10628 10609 10656
rect 9306 10588 9312 10600
rect 8444 10560 8984 10588
rect 9048 10560 9312 10588
rect 8444 10548 8450 10560
rect 8846 10520 8852 10532
rect 8312 10492 8852 10520
rect 8846 10480 8852 10492
rect 8904 10480 8910 10532
rect 3835 10424 4752 10452
rect 5721 10455 5779 10461
rect 3835 10421 3847 10424
rect 3789 10415 3847 10421
rect 5721 10421 5733 10455
rect 5767 10452 5779 10455
rect 5810 10452 5816 10464
rect 5767 10424 5816 10452
rect 5767 10421 5779 10424
rect 5721 10415 5779 10421
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 8956 10452 8984 10560
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 9968 10597 9996 10628
rect 10597 10625 10609 10628
rect 10643 10625 10655 10659
rect 10888 10656 10916 10696
rect 10965 10693 10977 10727
rect 11011 10724 11023 10727
rect 11057 10727 11115 10733
rect 11057 10724 11069 10727
rect 11011 10696 11069 10724
rect 11011 10693 11023 10696
rect 10965 10687 11023 10693
rect 11057 10693 11069 10696
rect 11103 10693 11115 10727
rect 12066 10724 12072 10736
rect 12027 10696 12072 10724
rect 11057 10687 11115 10693
rect 12066 10684 12072 10696
rect 12124 10684 12130 10736
rect 11977 10659 12035 10665
rect 11977 10656 11989 10659
rect 10888 10628 11989 10656
rect 10597 10619 10655 10625
rect 11977 10625 11989 10628
rect 12023 10656 12035 10659
rect 12434 10656 12440 10668
rect 12023 10628 12440 10656
rect 12023 10625 12035 10628
rect 11977 10619 12035 10625
rect 12434 10616 12440 10628
rect 12492 10616 12498 10668
rect 13280 10656 13308 10764
rect 14277 10727 14335 10733
rect 14277 10693 14289 10727
rect 14323 10724 14335 10727
rect 14369 10727 14427 10733
rect 14369 10724 14381 10727
rect 14323 10696 14381 10724
rect 14323 10693 14335 10696
rect 14277 10687 14335 10693
rect 14369 10693 14381 10696
rect 14415 10693 14427 10727
rect 14369 10687 14427 10693
rect 13909 10659 13967 10665
rect 13909 10656 13921 10659
rect 13280 10628 13921 10656
rect 9953 10591 10011 10597
rect 9953 10557 9965 10591
rect 9999 10557 10011 10591
rect 10502 10588 10508 10600
rect 10463 10560 10508 10588
rect 9953 10551 10011 10557
rect 9968 10452 9996 10551
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 11241 10591 11299 10597
rect 11241 10557 11253 10591
rect 11287 10557 11299 10591
rect 11882 10588 11888 10600
rect 11843 10560 11888 10588
rect 11241 10551 11299 10557
rect 10413 10523 10471 10529
rect 10413 10489 10425 10523
rect 10459 10489 10471 10523
rect 10520 10520 10548 10548
rect 11256 10520 11284 10551
rect 11882 10548 11888 10560
rect 11940 10548 11946 10600
rect 12161 10591 12219 10597
rect 12161 10557 12173 10591
rect 12207 10588 12219 10591
rect 12250 10588 12256 10600
rect 12207 10560 12256 10588
rect 12207 10557 12219 10560
rect 12161 10551 12219 10557
rect 12250 10548 12256 10560
rect 12308 10548 12314 10600
rect 13280 10597 13308 10628
rect 13909 10625 13921 10628
rect 13955 10625 13967 10659
rect 13909 10619 13967 10625
rect 13265 10591 13323 10597
rect 13265 10557 13277 10591
rect 13311 10557 13323 10591
rect 13265 10551 13323 10557
rect 13817 10591 13875 10597
rect 13817 10557 13829 10591
rect 13863 10588 13875 10591
rect 14553 10591 14611 10597
rect 14553 10588 14565 10591
rect 13863 10560 14565 10588
rect 13863 10557 13875 10560
rect 13817 10551 13875 10557
rect 14553 10557 14565 10560
rect 14599 10588 14611 10591
rect 15102 10588 15108 10600
rect 14599 10560 15108 10588
rect 14599 10557 14611 10560
rect 14553 10551 14611 10557
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 10520 10492 11284 10520
rect 13725 10523 13783 10529
rect 10413 10483 10471 10489
rect 13725 10489 13737 10523
rect 13771 10520 13783 10523
rect 13771 10492 14320 10520
rect 13771 10489 13783 10492
rect 13725 10483 13783 10489
rect 8956 10424 9996 10452
rect 10428 10452 10456 10483
rect 10870 10452 10876 10464
rect 10428 10424 10876 10452
rect 10870 10412 10876 10424
rect 10928 10452 10934 10464
rect 10965 10455 11023 10461
rect 10965 10452 10977 10455
rect 10928 10424 10977 10452
rect 10928 10412 10934 10424
rect 10965 10421 10977 10424
rect 11011 10421 11023 10455
rect 11698 10452 11704 10464
rect 11659 10424 11704 10452
rect 10965 10415 11023 10421
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 14292 10461 14320 10492
rect 14277 10455 14335 10461
rect 14277 10421 14289 10455
rect 14323 10452 14335 10455
rect 14645 10455 14703 10461
rect 14645 10452 14657 10455
rect 14323 10424 14657 10452
rect 14323 10421 14335 10424
rect 14277 10415 14335 10421
rect 14645 10421 14657 10424
rect 14691 10421 14703 10455
rect 14645 10415 14703 10421
rect 14737 10455 14795 10461
rect 14737 10421 14749 10455
rect 14783 10452 14795 10455
rect 15010 10452 15016 10464
rect 14783 10424 15016 10452
rect 14783 10421 14795 10424
rect 14737 10415 14795 10421
rect 15010 10412 15016 10424
rect 15068 10412 15074 10464
rect 1104 10362 16100 10384
rect 1104 10310 5980 10362
rect 6032 10310 6044 10362
rect 6096 10310 6108 10362
rect 6160 10310 6172 10362
rect 6224 10310 10979 10362
rect 11031 10310 11043 10362
rect 11095 10310 11107 10362
rect 11159 10310 11171 10362
rect 11223 10310 16100 10362
rect 1104 10288 16100 10310
rect 3050 10208 3056 10260
rect 3108 10248 3114 10260
rect 3605 10251 3663 10257
rect 3605 10248 3617 10251
rect 3108 10220 3617 10248
rect 3108 10208 3114 10220
rect 3605 10217 3617 10220
rect 3651 10248 3663 10251
rect 4430 10248 4436 10260
rect 3651 10220 4436 10248
rect 3651 10217 3663 10220
rect 3605 10211 3663 10217
rect 4430 10208 4436 10220
rect 4488 10208 4494 10260
rect 5810 10208 5816 10260
rect 5868 10248 5874 10260
rect 6181 10251 6239 10257
rect 6181 10248 6193 10251
rect 5868 10220 6193 10248
rect 5868 10208 5874 10220
rect 6181 10217 6193 10220
rect 6227 10217 6239 10251
rect 9398 10248 9404 10260
rect 6181 10211 6239 10217
rect 7576 10220 9404 10248
rect 4154 10140 4160 10192
rect 4212 10180 4218 10192
rect 5258 10180 5264 10192
rect 4212 10152 5264 10180
rect 4212 10140 4218 10152
rect 5258 10140 5264 10152
rect 5316 10180 5322 10192
rect 5353 10183 5411 10189
rect 5353 10180 5365 10183
rect 5316 10152 5365 10180
rect 5316 10140 5322 10152
rect 5353 10149 5365 10152
rect 5399 10149 5411 10183
rect 5353 10143 5411 10149
rect 6255 10152 7512 10180
rect 3697 10115 3755 10121
rect 3697 10081 3709 10115
rect 3743 10112 3755 10115
rect 4062 10112 4068 10124
rect 3743 10084 4068 10112
rect 3743 10081 3755 10084
rect 3697 10075 3755 10081
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 4338 10072 4344 10124
rect 4396 10112 4402 10124
rect 4433 10115 4491 10121
rect 4433 10112 4445 10115
rect 4396 10084 4445 10112
rect 4396 10072 4402 10084
rect 4433 10081 4445 10084
rect 4479 10081 4491 10115
rect 4706 10112 4712 10124
rect 4667 10084 4712 10112
rect 4433 10075 4491 10081
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 4798 10072 4804 10124
rect 4856 10112 4862 10124
rect 5810 10112 5816 10124
rect 4856 10084 4901 10112
rect 5771 10084 5816 10112
rect 4856 10072 4862 10084
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 6255 10121 6283 10152
rect 6240 10115 6298 10121
rect 6240 10081 6252 10115
rect 6286 10081 6298 10115
rect 6240 10075 6298 10081
rect 6549 10115 6607 10121
rect 6549 10081 6561 10115
rect 6595 10081 6607 10115
rect 6549 10075 6607 10081
rect 3878 10004 3884 10056
rect 3936 10044 3942 10056
rect 4249 10047 4307 10053
rect 4249 10044 4261 10047
rect 3936 10016 4261 10044
rect 3936 10004 3942 10016
rect 4249 10013 4261 10016
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10044 5779 10047
rect 6255 10044 6283 10075
rect 5767 10016 6283 10044
rect 5767 10013 5779 10016
rect 5721 10007 5779 10013
rect 1946 9936 1952 9988
rect 2004 9976 2010 9988
rect 6564 9976 6592 10075
rect 7484 10053 7512 10152
rect 7576 10121 7604 10220
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 10226 10208 10232 10260
rect 10284 10248 10290 10260
rect 12158 10248 12164 10260
rect 10284 10220 12164 10248
rect 10284 10208 10290 10220
rect 12158 10208 12164 10220
rect 12216 10248 12222 10260
rect 12216 10220 13676 10248
rect 12216 10208 12222 10220
rect 7742 10140 7748 10192
rect 7800 10140 7806 10192
rect 12250 10140 12256 10192
rect 12308 10180 12314 10192
rect 13648 10189 13676 10220
rect 13449 10183 13507 10189
rect 13449 10180 13461 10183
rect 12308 10152 13461 10180
rect 12308 10140 12314 10152
rect 13449 10149 13461 10152
rect 13495 10149 13507 10183
rect 13449 10143 13507 10149
rect 13633 10183 13691 10189
rect 13633 10149 13645 10183
rect 13679 10149 13691 10183
rect 15102 10180 15108 10192
rect 13633 10143 13691 10149
rect 14936 10152 15108 10180
rect 7561 10115 7619 10121
rect 7561 10081 7573 10115
rect 7607 10081 7619 10115
rect 7561 10075 7619 10081
rect 7653 10115 7711 10121
rect 7653 10081 7665 10115
rect 7699 10112 7711 10115
rect 7760 10112 7788 10140
rect 7699 10084 7788 10112
rect 7699 10081 7711 10084
rect 7653 10075 7711 10081
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 10229 10115 10287 10121
rect 10229 10112 10241 10115
rect 10008 10084 10241 10112
rect 10008 10072 10014 10084
rect 10229 10081 10241 10084
rect 10275 10081 10287 10115
rect 10229 10075 10287 10081
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10112 10563 10115
rect 10594 10112 10600 10124
rect 10551 10084 10600 10112
rect 10551 10081 10563 10084
rect 10505 10075 10563 10081
rect 10594 10072 10600 10084
rect 10652 10112 10658 10124
rect 12069 10115 12127 10121
rect 12069 10112 12081 10115
rect 10652 10084 12081 10112
rect 10652 10072 10658 10084
rect 12069 10081 12081 10084
rect 12115 10112 12127 10115
rect 12115 10084 12480 10112
rect 12115 10081 12127 10084
rect 12069 10075 12127 10081
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10044 7803 10047
rect 7791 10016 8294 10044
rect 7791 10013 7803 10016
rect 7745 10007 7803 10013
rect 2004 9948 6592 9976
rect 7484 9976 7512 10007
rect 7834 9976 7840 9988
rect 7484 9948 7840 9976
rect 2004 9936 2010 9948
rect 7834 9936 7840 9948
rect 7892 9936 7898 9988
rect 8266 9976 8294 10016
rect 9398 10004 9404 10056
rect 9456 10044 9462 10056
rect 10321 10047 10379 10053
rect 10321 10044 10333 10047
rect 9456 10016 10333 10044
rect 9456 10004 9462 10016
rect 10321 10013 10333 10016
rect 10367 10044 10379 10047
rect 11974 10044 11980 10056
rect 10367 10016 11980 10044
rect 10367 10013 10379 10016
rect 10321 10007 10379 10013
rect 11974 10004 11980 10016
rect 12032 10004 12038 10056
rect 12158 10044 12164 10056
rect 12119 10016 12164 10044
rect 12158 10004 12164 10016
rect 12216 10004 12222 10056
rect 12452 10044 12480 10084
rect 12526 10072 12532 10124
rect 12584 10112 12590 10124
rect 12621 10115 12679 10121
rect 12621 10112 12633 10115
rect 12584 10084 12633 10112
rect 12584 10072 12590 10084
rect 12621 10081 12633 10084
rect 12667 10081 12679 10115
rect 12802 10112 12808 10124
rect 12763 10084 12808 10112
rect 12621 10075 12679 10081
rect 12802 10072 12808 10084
rect 12860 10072 12866 10124
rect 12986 10112 12992 10124
rect 12947 10084 12992 10112
rect 12986 10072 12992 10084
rect 13044 10072 13050 10124
rect 14936 10121 14964 10152
rect 15102 10140 15108 10152
rect 15160 10140 15166 10192
rect 13081 10115 13139 10121
rect 13081 10081 13093 10115
rect 13127 10081 13139 10115
rect 13081 10075 13139 10081
rect 13357 10115 13415 10121
rect 13357 10081 13369 10115
rect 13403 10112 13415 10115
rect 14369 10115 14427 10121
rect 14369 10112 14381 10115
rect 13403 10084 14381 10112
rect 13403 10081 13415 10084
rect 13357 10075 13415 10081
rect 14369 10081 14381 10084
rect 14415 10081 14427 10115
rect 14369 10075 14427 10081
rect 14921 10115 14979 10121
rect 14921 10081 14933 10115
rect 14967 10081 14979 10115
rect 14921 10075 14979 10081
rect 13096 10044 13124 10075
rect 12452 10016 13124 10044
rect 14384 10044 14412 10075
rect 15010 10072 15016 10124
rect 15068 10112 15074 10124
rect 15746 10112 15752 10124
rect 15068 10084 15113 10112
rect 15707 10084 15752 10112
rect 15068 10072 15074 10084
rect 15746 10072 15752 10084
rect 15804 10072 15810 10124
rect 15381 10047 15439 10053
rect 15381 10044 15393 10047
rect 14384 10016 15393 10044
rect 15381 10013 15393 10016
rect 15427 10013 15439 10047
rect 15381 10007 15439 10013
rect 8846 9976 8852 9988
rect 8266 9948 8852 9976
rect 8846 9936 8852 9948
rect 8904 9976 8910 9988
rect 10413 9979 10471 9985
rect 10413 9976 10425 9979
rect 8904 9948 10425 9976
rect 8904 9936 8910 9948
rect 10413 9945 10425 9948
rect 10459 9976 10471 9979
rect 11882 9976 11888 9988
rect 10459 9948 11888 9976
rect 10459 9945 10471 9948
rect 10413 9939 10471 9945
rect 11882 9936 11888 9948
rect 11940 9976 11946 9988
rect 12253 9979 12311 9985
rect 12253 9976 12265 9979
rect 11940 9948 12265 9976
rect 11940 9936 11946 9948
rect 12253 9945 12265 9948
rect 12299 9976 12311 9979
rect 12299 9948 12940 9976
rect 12299 9945 12311 9948
rect 12253 9939 12311 9945
rect 12912 9920 12940 9948
rect 6362 9908 6368 9920
rect 6323 9880 6368 9908
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 6733 9911 6791 9917
rect 6733 9877 6745 9911
rect 6779 9908 6791 9911
rect 7006 9908 7012 9920
rect 6779 9880 7012 9908
rect 6779 9877 6791 9880
rect 6733 9871 6791 9877
rect 7006 9868 7012 9880
rect 7064 9868 7070 9920
rect 7282 9908 7288 9920
rect 7243 9880 7288 9908
rect 7282 9868 7288 9880
rect 7340 9868 7346 9920
rect 10042 9908 10048 9920
rect 10003 9880 10048 9908
rect 10042 9868 10048 9880
rect 10100 9868 10106 9920
rect 11790 9908 11796 9920
rect 11751 9880 11796 9908
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 11974 9868 11980 9920
rect 12032 9908 12038 9920
rect 12345 9911 12403 9917
rect 12345 9908 12357 9911
rect 12032 9880 12357 9908
rect 12032 9868 12038 9880
rect 12345 9877 12357 9880
rect 12391 9908 12403 9911
rect 12802 9908 12808 9920
rect 12391 9880 12808 9908
rect 12391 9877 12403 9880
rect 12345 9871 12403 9877
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 12894 9868 12900 9920
rect 12952 9908 12958 9920
rect 13814 9908 13820 9920
rect 12952 9880 12997 9908
rect 13775 9880 13820 9908
rect 12952 9868 12958 9880
rect 13814 9868 13820 9880
rect 13872 9868 13878 9920
rect 14921 9911 14979 9917
rect 14921 9877 14933 9911
rect 14967 9908 14979 9911
rect 15013 9911 15071 9917
rect 15013 9908 15025 9911
rect 14967 9880 15025 9908
rect 14967 9877 14979 9880
rect 14921 9871 14979 9877
rect 15013 9877 15025 9880
rect 15059 9908 15071 9911
rect 15286 9908 15292 9920
rect 15059 9880 15292 9908
rect 15059 9877 15071 9880
rect 15013 9871 15071 9877
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 15562 9908 15568 9920
rect 15523 9880 15568 9908
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 1104 9818 16100 9840
rect 1104 9766 3481 9818
rect 3533 9766 3545 9818
rect 3597 9766 3609 9818
rect 3661 9766 3673 9818
rect 3725 9766 8480 9818
rect 8532 9766 8544 9818
rect 8596 9766 8608 9818
rect 8660 9766 8672 9818
rect 8724 9766 13478 9818
rect 13530 9766 13542 9818
rect 13594 9766 13606 9818
rect 13658 9766 13670 9818
rect 13722 9766 16100 9818
rect 1104 9744 16100 9766
rect 2958 9704 2964 9716
rect 2919 9676 2964 9704
rect 2958 9664 2964 9676
rect 3016 9664 3022 9716
rect 7834 9664 7840 9716
rect 7892 9704 7898 9716
rect 8205 9707 8263 9713
rect 8205 9704 8217 9707
rect 7892 9676 8217 9704
rect 7892 9664 7898 9676
rect 8205 9673 8217 9676
rect 8251 9673 8263 9707
rect 8205 9667 8263 9673
rect 10502 9664 10508 9716
rect 10560 9704 10566 9716
rect 11057 9707 11115 9713
rect 11057 9704 11069 9707
rect 10560 9676 11069 9704
rect 10560 9664 10566 9676
rect 11057 9673 11069 9676
rect 11103 9673 11115 9707
rect 11057 9667 11115 9673
rect 3234 9636 3240 9648
rect 2746 9608 3240 9636
rect 2746 9568 2774 9608
rect 3234 9596 3240 9608
rect 3292 9596 3298 9648
rect 2700 9540 2774 9568
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 1946 9460 1952 9512
rect 2004 9500 2010 9512
rect 2700 9509 2728 9540
rect 6362 9528 6368 9580
rect 6420 9568 6426 9580
rect 6733 9571 6791 9577
rect 6733 9568 6745 9571
rect 6420 9540 6745 9568
rect 6420 9528 6426 9540
rect 6733 9537 6745 9540
rect 6779 9537 6791 9571
rect 6733 9531 6791 9537
rect 2041 9503 2099 9509
rect 2041 9500 2053 9503
rect 2004 9472 2053 9500
rect 2004 9460 2010 9472
rect 2041 9469 2053 9472
rect 2087 9469 2099 9503
rect 2041 9463 2099 9469
rect 2685 9503 2743 9509
rect 2685 9469 2697 9503
rect 2731 9469 2743 9503
rect 2685 9463 2743 9469
rect 2774 9460 2780 9512
rect 2832 9500 2838 9512
rect 3053 9503 3111 9509
rect 2832 9472 2877 9500
rect 2832 9460 2838 9472
rect 3053 9469 3065 9503
rect 3099 9500 3111 9503
rect 3326 9500 3332 9512
rect 3099 9472 3332 9500
rect 3099 9469 3111 9472
rect 3053 9463 3111 9469
rect 3326 9460 3332 9472
rect 3384 9460 3390 9512
rect 5718 9460 5724 9512
rect 5776 9500 5782 9512
rect 6457 9503 6515 9509
rect 6457 9500 6469 9503
rect 5776 9472 6469 9500
rect 5776 9460 5782 9472
rect 6457 9469 6469 9472
rect 6503 9469 6515 9503
rect 6457 9463 6515 9469
rect 8757 9503 8815 9509
rect 8757 9469 8769 9503
rect 8803 9500 8815 9503
rect 9030 9500 9036 9512
rect 8803 9472 9036 9500
rect 8803 9469 8815 9472
rect 8757 9463 8815 9469
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9585 9503 9643 9509
rect 9585 9469 9597 9503
rect 9631 9500 9643 9503
rect 9674 9500 9680 9512
rect 9631 9472 9680 9500
rect 9631 9469 9643 9472
rect 9585 9463 9643 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 15286 9500 15292 9512
rect 15247 9472 15292 9500
rect 15286 9460 15292 9472
rect 15344 9460 15350 9512
rect 5810 9432 5816 9444
rect 1596 9404 5816 9432
rect 1596 9373 1624 9404
rect 5810 9392 5816 9404
rect 5868 9392 5874 9444
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 7064 9404 7222 9432
rect 7064 9392 7070 9404
rect 8110 9392 8116 9444
rect 8168 9432 8174 9444
rect 8389 9435 8447 9441
rect 8389 9432 8401 9435
rect 8168 9404 8401 9432
rect 8168 9392 8174 9404
rect 8389 9401 8401 9404
rect 8435 9401 8447 9435
rect 8389 9395 8447 9401
rect 8573 9435 8631 9441
rect 8573 9401 8585 9435
rect 8619 9432 8631 9435
rect 8846 9432 8852 9444
rect 8619 9404 8852 9432
rect 8619 9401 8631 9404
rect 8573 9395 8631 9401
rect 8846 9392 8852 9404
rect 8904 9392 8910 9444
rect 10594 9392 10600 9444
rect 10652 9432 10658 9444
rect 10965 9435 11023 9441
rect 10965 9432 10977 9435
rect 10652 9404 10977 9432
rect 10652 9392 10658 9404
rect 10965 9401 10977 9404
rect 11011 9401 11023 9435
rect 15102 9432 15108 9444
rect 15063 9404 15108 9432
rect 10965 9395 11023 9401
rect 15102 9392 15108 9404
rect 15160 9392 15166 9444
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9333 1639 9367
rect 2222 9364 2228 9376
rect 2183 9336 2228 9364
rect 1581 9327 1639 9333
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 2498 9364 2504 9376
rect 2459 9336 2504 9364
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 9766 9364 9772 9376
rect 9727 9336 9772 9364
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 1104 9274 16100 9296
rect 1104 9222 5980 9274
rect 6032 9222 6044 9274
rect 6096 9222 6108 9274
rect 6160 9222 6172 9274
rect 6224 9222 10979 9274
rect 11031 9222 11043 9274
rect 11095 9222 11107 9274
rect 11159 9222 11171 9274
rect 11223 9222 16100 9274
rect 1104 9200 16100 9222
rect 2498 9160 2504 9172
rect 1688 9132 2504 9160
rect 1688 9101 1716 9132
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 8110 9160 8116 9172
rect 3896 9132 8116 9160
rect 1673 9095 1731 9101
rect 1673 9061 1685 9095
rect 1719 9061 1731 9095
rect 1673 9055 1731 9061
rect 2222 9052 2228 9104
rect 2280 9052 2286 9104
rect 3896 9033 3924 9132
rect 8110 9120 8116 9132
rect 8168 9120 8174 9172
rect 9674 9160 9680 9172
rect 9508 9132 9680 9160
rect 5810 9052 5816 9104
rect 5868 9092 5874 9104
rect 6181 9095 6239 9101
rect 6181 9092 6193 9095
rect 5868 9064 6193 9092
rect 5868 9052 5874 9064
rect 6181 9061 6193 9064
rect 6227 9092 6239 9095
rect 6914 9092 6920 9104
rect 6227 9064 6920 9092
rect 6227 9061 6239 9064
rect 6181 9055 6239 9061
rect 6914 9052 6920 9064
rect 6972 9052 6978 9104
rect 3881 9027 3939 9033
rect 3881 8993 3893 9027
rect 3927 8993 3939 9027
rect 4062 9024 4068 9036
rect 4023 8996 4068 9024
rect 3881 8987 3939 8993
rect 4062 8984 4068 8996
rect 4120 8984 4126 9036
rect 4430 8984 4436 9036
rect 4488 9024 4494 9036
rect 4525 9027 4583 9033
rect 4525 9024 4537 9027
rect 4488 8996 4537 9024
rect 4488 8984 4494 8996
rect 4525 8993 4537 8996
rect 4571 8993 4583 9027
rect 4706 9024 4712 9036
rect 4667 8996 4712 9024
rect 4525 8987 4583 8993
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 5169 9027 5227 9033
rect 5169 8993 5181 9027
rect 5215 9024 5227 9027
rect 5350 9024 5356 9036
rect 5215 8996 5356 9024
rect 5215 8993 5227 8996
rect 5169 8987 5227 8993
rect 5350 8984 5356 8996
rect 5408 8984 5414 9036
rect 5905 9027 5963 9033
rect 5905 8993 5917 9027
rect 5951 9024 5963 9027
rect 6365 9027 6423 9033
rect 5951 8996 6040 9024
rect 5951 8993 5963 8996
rect 5905 8987 5963 8993
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8956 1455 8959
rect 1670 8956 1676 8968
rect 1443 8928 1676 8956
rect 1443 8925 1455 8928
rect 1397 8919 1455 8925
rect 1670 8916 1676 8928
rect 1728 8956 1734 8968
rect 5718 8956 5724 8968
rect 1728 8928 5724 8956
rect 1728 8916 1734 8928
rect 5718 8916 5724 8928
rect 5776 8916 5782 8968
rect 3145 8823 3203 8829
rect 3145 8789 3157 8823
rect 3191 8820 3203 8823
rect 3326 8820 3332 8832
rect 3191 8792 3332 8820
rect 3191 8789 3203 8792
rect 3145 8783 3203 8789
rect 3326 8780 3332 8792
rect 3384 8820 3390 8832
rect 3881 8823 3939 8829
rect 3881 8820 3893 8823
rect 3384 8792 3893 8820
rect 3384 8780 3390 8792
rect 3881 8789 3893 8792
rect 3927 8789 3939 8823
rect 3881 8783 3939 8789
rect 4154 8780 4160 8832
rect 4212 8820 4218 8832
rect 4249 8823 4307 8829
rect 4249 8820 4261 8823
rect 4212 8792 4261 8820
rect 4212 8780 4218 8792
rect 4249 8789 4261 8792
rect 4295 8789 4307 8823
rect 4249 8783 4307 8789
rect 4614 8780 4620 8832
rect 4672 8820 4678 8832
rect 4801 8823 4859 8829
rect 4801 8820 4813 8823
rect 4672 8792 4813 8820
rect 4672 8780 4678 8792
rect 4801 8789 4813 8792
rect 4847 8789 4859 8823
rect 5258 8820 5264 8832
rect 5219 8792 5264 8820
rect 4801 8783 4859 8789
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 5810 8820 5816 8832
rect 5771 8792 5816 8820
rect 5810 8780 5816 8792
rect 5868 8780 5874 8832
rect 6012 8829 6040 8996
rect 6365 8993 6377 9027
rect 6411 9024 6423 9027
rect 6822 9024 6828 9036
rect 6411 8996 6828 9024
rect 6411 8993 6423 8996
rect 6365 8987 6423 8993
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 9122 9024 9128 9036
rect 9083 8996 9128 9024
rect 9122 8984 9128 8996
rect 9180 8984 9186 9036
rect 9508 9024 9536 9132
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 9769 9163 9827 9169
rect 9769 9129 9781 9163
rect 9815 9129 9827 9163
rect 10594 9160 10600 9172
rect 10555 9132 10600 9160
rect 9769 9123 9827 9129
rect 9585 9095 9643 9101
rect 9585 9061 9597 9095
rect 9631 9092 9643 9095
rect 9784 9092 9812 9123
rect 10594 9120 10600 9132
rect 10652 9120 10658 9172
rect 10689 9095 10747 9101
rect 10689 9092 10701 9095
rect 9631 9064 10701 9092
rect 9631 9061 9643 9064
rect 9585 9055 9643 9061
rect 10689 9061 10701 9064
rect 10735 9061 10747 9095
rect 10689 9055 10747 9061
rect 12894 9052 12900 9104
rect 12952 9092 12958 9104
rect 12952 9064 13584 9092
rect 12952 9052 12958 9064
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 9508 8996 9689 9024
rect 9677 8993 9689 8996
rect 9723 8993 9735 9027
rect 9677 8987 9735 8993
rect 10042 8984 10048 9036
rect 10100 9024 10106 9036
rect 10229 9027 10287 9033
rect 10229 9024 10241 9027
rect 10100 8996 10241 9024
rect 10100 8984 10106 8996
rect 10229 8993 10241 8996
rect 10275 8993 10287 9027
rect 12526 9024 12532 9036
rect 12487 8996 12532 9024
rect 10229 8987 10287 8993
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 13081 9027 13139 9033
rect 13081 8993 13093 9027
rect 13127 9024 13139 9027
rect 13170 9024 13176 9036
rect 13127 8996 13176 9024
rect 13127 8993 13139 8996
rect 13081 8987 13139 8993
rect 13170 8984 13176 8996
rect 13228 8984 13234 9036
rect 13556 9033 13584 9064
rect 13265 9027 13323 9033
rect 13265 8993 13277 9027
rect 13311 8993 13323 9027
rect 13265 8987 13323 8993
rect 13541 9027 13599 9033
rect 13541 8993 13553 9027
rect 13587 8993 13599 9027
rect 13541 8987 13599 8993
rect 9140 8956 9168 8984
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9140 8928 10149 8956
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 12989 8959 13047 8965
rect 12989 8925 13001 8959
rect 13035 8956 13047 8959
rect 13280 8956 13308 8987
rect 13354 8956 13360 8968
rect 13035 8928 13360 8956
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 9766 8888 9772 8900
rect 9727 8860 9772 8888
rect 9766 8848 9772 8860
rect 9824 8848 9830 8900
rect 10597 8891 10655 8897
rect 10597 8857 10609 8891
rect 10643 8888 10655 8891
rect 10781 8891 10839 8897
rect 10781 8888 10793 8891
rect 10643 8860 10793 8888
rect 10643 8857 10655 8860
rect 10597 8851 10655 8857
rect 10781 8857 10793 8860
rect 10827 8857 10839 8891
rect 10781 8851 10839 8857
rect 5997 8823 6055 8829
rect 5997 8789 6009 8823
rect 6043 8820 6055 8823
rect 6086 8820 6092 8832
rect 6043 8792 6092 8820
rect 6043 8789 6055 8792
rect 5997 8783 6055 8789
rect 6086 8780 6092 8792
rect 6144 8780 6150 8832
rect 13262 8820 13268 8832
rect 13223 8792 13268 8820
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 13725 8823 13783 8829
rect 13725 8789 13737 8823
rect 13771 8820 13783 8823
rect 14182 8820 14188 8832
rect 13771 8792 14188 8820
rect 13771 8789 13783 8792
rect 13725 8783 13783 8789
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 1104 8730 16100 8752
rect 1104 8678 3481 8730
rect 3533 8678 3545 8730
rect 3597 8678 3609 8730
rect 3661 8678 3673 8730
rect 3725 8678 8480 8730
rect 8532 8678 8544 8730
rect 8596 8678 8608 8730
rect 8660 8678 8672 8730
rect 8724 8678 13478 8730
rect 13530 8678 13542 8730
rect 13594 8678 13606 8730
rect 13658 8678 13670 8730
rect 13722 8678 16100 8730
rect 1104 8656 16100 8678
rect 3789 8619 3847 8625
rect 3789 8585 3801 8619
rect 3835 8616 3847 8619
rect 4706 8616 4712 8628
rect 3835 8588 4568 8616
rect 4667 8588 4712 8616
rect 3835 8585 3847 8588
rect 3789 8579 3847 8585
rect 2409 8551 2467 8557
rect 2409 8517 2421 8551
rect 2455 8548 2467 8551
rect 4338 8548 4344 8560
rect 2455 8520 4344 8548
rect 2455 8517 2467 8520
rect 2409 8511 2467 8517
rect 4338 8508 4344 8520
rect 4396 8508 4402 8560
rect 4154 8480 4160 8492
rect 4115 8452 4160 8480
rect 4154 8440 4160 8452
rect 4212 8440 4218 8492
rect 4540 8480 4568 8588
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 10318 8616 10324 8628
rect 5000 8588 10324 8616
rect 4617 8551 4675 8557
rect 4617 8517 4629 8551
rect 4663 8548 4675 8551
rect 4798 8548 4804 8560
rect 4663 8520 4804 8548
rect 4663 8517 4675 8520
rect 4617 8511 4675 8517
rect 4798 8508 4804 8520
rect 4856 8508 4862 8560
rect 5000 8480 5028 8588
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 10505 8619 10563 8625
rect 10505 8585 10517 8619
rect 10551 8616 10563 8619
rect 10594 8616 10600 8628
rect 10551 8588 10600 8616
rect 10551 8585 10563 8588
rect 10505 8579 10563 8585
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 5350 8508 5356 8560
rect 5408 8548 5414 8560
rect 5629 8551 5687 8557
rect 5629 8548 5641 8551
rect 5408 8520 5641 8548
rect 5408 8508 5414 8520
rect 5629 8517 5641 8520
rect 5675 8517 5687 8551
rect 6638 8548 6644 8560
rect 5629 8511 5687 8517
rect 5920 8520 6644 8548
rect 4540 8452 5028 8480
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8480 5135 8483
rect 5810 8480 5816 8492
rect 5123 8452 5816 8480
rect 5123 8449 5135 8452
rect 5077 8443 5135 8449
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 2222 8412 2228 8424
rect 2183 8384 2228 8412
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 2314 8372 2320 8424
rect 2372 8412 2378 8424
rect 2409 8415 2467 8421
rect 2409 8412 2421 8415
rect 2372 8384 2421 8412
rect 2372 8372 2378 8384
rect 2409 8381 2421 8384
rect 2455 8381 2467 8415
rect 2409 8375 2467 8381
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8412 3847 8415
rect 3881 8415 3939 8421
rect 3881 8412 3893 8415
rect 3835 8384 3893 8412
rect 3835 8381 3847 8384
rect 3789 8375 3847 8381
rect 3881 8381 3893 8384
rect 3927 8381 3939 8415
rect 3881 8375 3939 8381
rect 4065 8415 4123 8421
rect 4065 8381 4077 8415
rect 4111 8381 4123 8415
rect 4065 8375 4123 8381
rect 4080 8344 4108 8375
rect 4246 8372 4252 8424
rect 4304 8412 4310 8424
rect 4430 8412 4436 8424
rect 4304 8384 4349 8412
rect 4391 8384 4436 8412
rect 4304 8372 4310 8384
rect 4430 8372 4436 8384
rect 4488 8372 4494 8424
rect 4893 8415 4951 8421
rect 4893 8381 4905 8415
rect 4939 8381 4951 8415
rect 5166 8412 5172 8424
rect 5127 8384 5172 8412
rect 4893 8375 4951 8381
rect 4614 8344 4620 8356
rect 4080 8316 4620 8344
rect 4614 8304 4620 8316
rect 4672 8304 4678 8356
rect 4908 8344 4936 8375
rect 5166 8372 5172 8384
rect 5224 8372 5230 8424
rect 5258 8372 5264 8424
rect 5316 8412 5322 8424
rect 5442 8412 5448 8424
rect 5316 8384 5361 8412
rect 5403 8384 5448 8412
rect 5316 8372 5322 8384
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 5920 8421 5948 8520
rect 6638 8508 6644 8520
rect 6696 8508 6702 8560
rect 13078 8548 13084 8560
rect 13039 8520 13084 8548
rect 13078 8508 13084 8520
rect 13136 8508 13142 8560
rect 13354 8508 13360 8560
rect 13412 8548 13418 8560
rect 13541 8551 13599 8557
rect 13541 8548 13553 8551
rect 13412 8520 13553 8548
rect 13412 8508 13418 8520
rect 13541 8517 13553 8520
rect 13587 8517 13599 8551
rect 13541 8511 13599 8517
rect 15197 8551 15255 8557
rect 15197 8517 15209 8551
rect 15243 8548 15255 8551
rect 15289 8551 15347 8557
rect 15289 8548 15301 8551
rect 15243 8520 15301 8548
rect 15243 8517 15255 8520
rect 15197 8511 15255 8517
rect 15289 8517 15301 8520
rect 15335 8517 15347 8551
rect 15289 8511 15347 8517
rect 6012 8452 6592 8480
rect 6012 8421 6040 8452
rect 6564 8424 6592 8452
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 6880 8452 7144 8480
rect 6880 8440 6886 8452
rect 5905 8415 5963 8421
rect 5905 8381 5917 8415
rect 5951 8381 5963 8415
rect 5905 8375 5963 8381
rect 5997 8415 6055 8421
rect 5997 8381 6009 8415
rect 6043 8381 6055 8415
rect 5997 8375 6055 8381
rect 6086 8372 6092 8424
rect 6144 8412 6150 8424
rect 6273 8415 6331 8421
rect 6144 8384 6189 8412
rect 6144 8372 6150 8384
rect 6273 8381 6285 8415
rect 6319 8381 6331 8415
rect 6546 8412 6552 8424
rect 6507 8384 6552 8412
rect 6273 8375 6331 8381
rect 6288 8344 6316 8375
rect 6546 8372 6552 8384
rect 6604 8372 6610 8424
rect 6638 8372 6644 8424
rect 6696 8412 6702 8424
rect 6914 8412 6920 8424
rect 6696 8384 6741 8412
rect 6875 8384 6920 8412
rect 6696 8372 6702 8384
rect 6914 8372 6920 8384
rect 6972 8372 6978 8424
rect 7116 8421 7144 8452
rect 7282 8440 7288 8492
rect 7340 8480 7346 8492
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 7340 8452 7389 8480
rect 7340 8440 7346 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 9674 8440 9680 8492
rect 9732 8480 9738 8492
rect 9732 8452 10548 8480
rect 9732 8440 9738 8452
rect 7101 8415 7159 8421
rect 7101 8381 7113 8415
rect 7147 8381 7159 8415
rect 7101 8375 7159 8381
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8412 7803 8415
rect 8662 8412 8668 8424
rect 7791 8384 8668 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 9953 8415 10011 8421
rect 9953 8381 9965 8415
rect 9999 8412 10011 8415
rect 10042 8412 10048 8424
rect 9999 8384 10048 8412
rect 9999 8381 10011 8384
rect 9953 8375 10011 8381
rect 10042 8372 10048 8384
rect 10100 8372 10106 8424
rect 10520 8421 10548 8452
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 14001 8483 14059 8489
rect 14001 8480 14013 8483
rect 12584 8452 14013 8480
rect 12584 8440 12590 8452
rect 14001 8449 14013 8452
rect 14047 8449 14059 8483
rect 14829 8483 14887 8489
rect 14829 8480 14841 8483
rect 14001 8443 14059 8449
rect 14200 8452 14841 8480
rect 14200 8424 14228 8452
rect 14829 8449 14841 8452
rect 14875 8449 14887 8483
rect 14829 8443 14887 8449
rect 10505 8415 10563 8421
rect 10505 8381 10517 8415
rect 10551 8381 10563 8415
rect 11790 8412 11796 8424
rect 11751 8384 11796 8412
rect 10505 8375 10563 8381
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 13170 8372 13176 8424
rect 13228 8412 13234 8424
rect 13265 8415 13323 8421
rect 13265 8412 13277 8415
rect 13228 8384 13277 8412
rect 13228 8372 13234 8384
rect 13265 8381 13277 8384
rect 13311 8412 13323 8415
rect 13630 8412 13636 8424
rect 13311 8384 13636 8412
rect 13311 8381 13323 8384
rect 13265 8375 13323 8381
rect 13630 8372 13636 8384
rect 13688 8372 13694 8424
rect 14182 8412 14188 8424
rect 14143 8384 14188 8412
rect 14182 8372 14188 8384
rect 14240 8372 14246 8424
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 14737 8415 14795 8421
rect 14737 8412 14749 8415
rect 14608 8384 14749 8412
rect 14608 8372 14614 8384
rect 14737 8381 14749 8384
rect 14783 8412 14795 8415
rect 15102 8412 15108 8424
rect 14783 8384 15108 8412
rect 14783 8381 14795 8384
rect 14737 8375 14795 8381
rect 15102 8372 15108 8384
rect 15160 8412 15166 8424
rect 15473 8415 15531 8421
rect 15473 8412 15485 8415
rect 15160 8384 15485 8412
rect 15160 8372 15166 8384
rect 15473 8381 15485 8384
rect 15519 8381 15531 8415
rect 15473 8375 15531 8381
rect 6825 8347 6883 8353
rect 6825 8344 6837 8347
rect 4908 8316 6837 8344
rect 6825 8313 6837 8316
rect 6871 8313 6883 8347
rect 8386 8344 8392 8356
rect 8347 8316 8392 8344
rect 6825 8307 6883 8313
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 13446 8344 13452 8356
rect 13407 8316 13452 8344
rect 13446 8304 13452 8316
rect 13504 8304 13510 8356
rect 14645 8347 14703 8353
rect 14645 8313 14657 8347
rect 14691 8313 14703 8347
rect 14645 8307 14703 8313
rect 4338 8236 4344 8288
rect 4396 8276 4402 8288
rect 5442 8276 5448 8288
rect 4396 8248 5448 8276
rect 4396 8236 4402 8248
rect 5442 8236 5448 8248
rect 5500 8236 5506 8288
rect 7742 8276 7748 8288
rect 7703 8248 7748 8276
rect 7742 8236 7748 8248
rect 7800 8276 7806 8288
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 7800 8248 8217 8276
rect 7800 8236 7806 8248
rect 8205 8245 8217 8248
rect 8251 8245 8263 8279
rect 14660 8276 14688 8307
rect 14734 8276 14740 8288
rect 14647 8248 14740 8276
rect 8205 8239 8263 8245
rect 14734 8236 14740 8248
rect 14792 8276 14798 8288
rect 15197 8279 15255 8285
rect 15197 8276 15209 8279
rect 14792 8248 15209 8276
rect 14792 8236 14798 8248
rect 15197 8245 15209 8248
rect 15243 8245 15255 8279
rect 15197 8239 15255 8245
rect 1104 8186 16100 8208
rect 1104 8134 5980 8186
rect 6032 8134 6044 8186
rect 6096 8134 6108 8186
rect 6160 8134 6172 8186
rect 6224 8134 10979 8186
rect 11031 8134 11043 8186
rect 11095 8134 11107 8186
rect 11159 8134 11171 8186
rect 11223 8134 16100 8186
rect 1104 8112 16100 8134
rect 8573 8075 8631 8081
rect 8573 8041 8585 8075
rect 8619 8041 8631 8075
rect 8573 8035 8631 8041
rect 2038 8004 2044 8016
rect 1872 7976 2044 8004
rect 1872 7945 1900 7976
rect 2038 7964 2044 7976
rect 2096 8004 2102 8016
rect 2961 8007 3019 8013
rect 2961 8004 2973 8007
rect 2096 7976 2973 8004
rect 2096 7964 2102 7976
rect 2961 7973 2973 7976
rect 3007 7973 3019 8007
rect 4246 8004 4252 8016
rect 4207 7976 4252 8004
rect 2961 7967 3019 7973
rect 4246 7964 4252 7976
rect 4304 7964 4310 8016
rect 5350 8004 5356 8016
rect 4908 7976 5356 8004
rect 1857 7939 1915 7945
rect 1857 7905 1869 7939
rect 1903 7905 1915 7939
rect 2314 7936 2320 7948
rect 2275 7908 2320 7936
rect 1857 7899 1915 7905
rect 2314 7896 2320 7908
rect 2372 7896 2378 7948
rect 2682 7936 2688 7948
rect 2643 7908 2688 7936
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 3142 7936 3148 7948
rect 3103 7908 3148 7936
rect 3142 7896 3148 7908
rect 3200 7896 3206 7948
rect 3326 7936 3332 7948
rect 3287 7908 3332 7936
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 4338 7936 4344 7948
rect 4299 7908 4344 7936
rect 4338 7896 4344 7908
rect 4396 7896 4402 7948
rect 4908 7945 4936 7976
rect 5350 7964 5356 7976
rect 5408 7964 5414 8016
rect 7742 8004 7748 8016
rect 7703 7976 7748 8004
rect 7742 7964 7748 7976
rect 7800 7964 7806 8016
rect 8588 8004 8616 8035
rect 8662 8032 8668 8084
rect 8720 8072 8726 8084
rect 9674 8072 9680 8084
rect 8720 8044 8765 8072
rect 9635 8044 9680 8072
rect 8720 8032 8726 8044
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 13446 8072 13452 8084
rect 13407 8044 13452 8072
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 14734 8072 14740 8084
rect 14695 8044 14740 8072
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 8938 8004 8944 8016
rect 8588 7976 8944 8004
rect 8938 7964 8944 7976
rect 8996 8004 9002 8016
rect 9585 8007 9643 8013
rect 9585 8004 9597 8007
rect 8996 7976 9597 8004
rect 8996 7964 9002 7976
rect 9585 7973 9597 7976
rect 9631 7973 9643 8007
rect 9585 7967 9643 7973
rect 4893 7939 4951 7945
rect 4893 7905 4905 7939
rect 4939 7905 4951 7939
rect 5074 7936 5080 7948
rect 5035 7908 5080 7936
rect 4893 7899 4951 7905
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 5626 7936 5632 7948
rect 5587 7908 5632 7936
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 5810 7936 5816 7948
rect 5771 7908 5816 7936
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 7282 7936 7288 7948
rect 7243 7908 7288 7936
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 7883 7908 8340 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 2222 7868 2228 7880
rect 2183 7840 2228 7868
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 2590 7868 2596 7880
rect 2551 7840 2596 7868
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 8110 7828 8116 7880
rect 8168 7868 8174 7880
rect 8205 7871 8263 7877
rect 8205 7868 8217 7871
rect 8168 7840 8217 7868
rect 8168 7828 8174 7840
rect 8205 7837 8217 7840
rect 8251 7837 8263 7871
rect 8312 7868 8340 7908
rect 8386 7896 8392 7948
rect 8444 7936 8450 7948
rect 8573 7939 8631 7945
rect 8573 7936 8585 7939
rect 8444 7908 8585 7936
rect 8444 7896 8450 7908
rect 8573 7905 8585 7908
rect 8619 7905 8631 7939
rect 8846 7936 8852 7948
rect 8807 7908 8852 7936
rect 8573 7899 8631 7905
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 11790 7936 11796 7948
rect 11751 7908 11796 7936
rect 11790 7896 11796 7908
rect 11848 7896 11854 7948
rect 13262 7936 13268 7948
rect 13223 7908 13268 7936
rect 13262 7896 13268 7908
rect 13320 7896 13326 7948
rect 13630 7936 13636 7948
rect 13543 7908 13636 7936
rect 13630 7896 13636 7908
rect 13688 7936 13694 7948
rect 14645 7939 14703 7945
rect 13688 7908 14504 7936
rect 13688 7896 13694 7908
rect 8864 7868 8892 7896
rect 13078 7868 13084 7880
rect 8312 7840 8892 7868
rect 13039 7840 13084 7868
rect 8205 7831 8263 7837
rect 13078 7828 13084 7840
rect 13136 7828 13142 7880
rect 2501 7803 2559 7809
rect 2501 7769 2513 7803
rect 2547 7800 2559 7803
rect 4430 7800 4436 7812
rect 2547 7772 4436 7800
rect 2547 7769 2559 7772
rect 2501 7763 2559 7769
rect 4430 7760 4436 7772
rect 4488 7760 4494 7812
rect 14476 7809 14504 7908
rect 14645 7905 14657 7939
rect 14691 7936 14703 7939
rect 14734 7936 14740 7948
rect 14691 7908 14740 7936
rect 14691 7905 14703 7908
rect 14645 7899 14703 7905
rect 14734 7896 14740 7908
rect 14792 7896 14798 7948
rect 14461 7803 14519 7809
rect 14461 7769 14473 7803
rect 14507 7769 14519 7803
rect 14461 7763 14519 7769
rect 14829 7735 14887 7741
rect 14829 7701 14841 7735
rect 14875 7732 14887 7735
rect 15010 7732 15016 7744
rect 14875 7704 15016 7732
rect 14875 7701 14887 7704
rect 14829 7695 14887 7701
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 1104 7642 16100 7664
rect 1104 7590 3481 7642
rect 3533 7590 3545 7642
rect 3597 7590 3609 7642
rect 3661 7590 3673 7642
rect 3725 7590 8480 7642
rect 8532 7590 8544 7642
rect 8596 7590 8608 7642
rect 8660 7590 8672 7642
rect 8724 7590 13478 7642
rect 13530 7590 13542 7642
rect 13594 7590 13606 7642
rect 13658 7590 13670 7642
rect 13722 7590 16100 7642
rect 1104 7568 16100 7590
rect 2314 7488 2320 7540
rect 2372 7528 2378 7540
rect 2685 7531 2743 7537
rect 2685 7528 2697 7531
rect 2372 7500 2697 7528
rect 2372 7488 2378 7500
rect 2685 7497 2697 7500
rect 2731 7497 2743 7531
rect 2685 7491 2743 7497
rect 5169 7531 5227 7537
rect 5169 7497 5181 7531
rect 5215 7528 5227 7531
rect 5810 7528 5816 7540
rect 5215 7500 5816 7528
rect 5215 7497 5227 7500
rect 5169 7491 5227 7497
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 8757 7531 8815 7537
rect 8757 7497 8769 7531
rect 8803 7528 8815 7531
rect 8938 7528 8944 7540
rect 8803 7500 8944 7528
rect 8803 7497 8815 7500
rect 8757 7491 8815 7497
rect 8938 7488 8944 7500
rect 8996 7488 9002 7540
rect 3142 7460 3148 7472
rect 2424 7432 3148 7460
rect 2038 7392 2044 7404
rect 1999 7364 2044 7392
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 2424 7401 2452 7432
rect 3142 7420 3148 7432
rect 3200 7460 3206 7472
rect 3329 7463 3387 7469
rect 3329 7460 3341 7463
rect 3200 7432 3341 7460
rect 3200 7420 3206 7432
rect 3329 7429 3341 7432
rect 3375 7429 3387 7463
rect 3329 7423 3387 7429
rect 10781 7463 10839 7469
rect 10781 7429 10793 7463
rect 10827 7460 10839 7463
rect 11057 7463 11115 7469
rect 11057 7460 11069 7463
rect 10827 7432 11069 7460
rect 10827 7429 10839 7432
rect 10781 7423 10839 7429
rect 11057 7429 11069 7432
rect 11103 7429 11115 7463
rect 15010 7460 15016 7472
rect 14971 7432 15016 7460
rect 11057 7423 11115 7429
rect 15010 7420 15016 7432
rect 15068 7420 15074 7472
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7361 2467 7395
rect 2409 7355 2467 7361
rect 2682 7352 2688 7404
rect 2740 7392 2746 7404
rect 3513 7395 3571 7401
rect 3513 7392 3525 7395
rect 2740 7364 3525 7392
rect 2740 7352 2746 7364
rect 2792 7333 2820 7364
rect 3513 7361 3525 7364
rect 3559 7361 3571 7395
rect 10410 7392 10416 7404
rect 10371 7364 10416 7392
rect 3513 7355 3571 7361
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 14645 7395 14703 7401
rect 14645 7392 14657 7395
rect 14016 7364 14657 7392
rect 2501 7327 2559 7333
rect 2501 7293 2513 7327
rect 2547 7293 2559 7327
rect 2501 7287 2559 7293
rect 2777 7327 2835 7333
rect 2777 7293 2789 7327
rect 2823 7324 2835 7327
rect 3142 7324 3148 7336
rect 2823 7296 2857 7324
rect 3103 7296 3148 7324
rect 2823 7293 2835 7296
rect 2777 7287 2835 7293
rect 2516 7188 2544 7287
rect 3142 7284 3148 7296
rect 3200 7324 3206 7336
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 3200 7296 3433 7324
rect 3200 7284 3206 7296
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 4522 7284 4528 7336
rect 4580 7324 4586 7336
rect 5077 7327 5135 7333
rect 5077 7324 5089 7327
rect 4580 7296 5089 7324
rect 4580 7284 4586 7296
rect 5077 7293 5089 7296
rect 5123 7324 5135 7327
rect 5442 7324 5448 7336
rect 5123 7296 5448 7324
rect 5123 7293 5135 7296
rect 5077 7287 5135 7293
rect 5442 7284 5448 7296
rect 5500 7284 5506 7336
rect 8110 7284 8116 7336
rect 8168 7324 8174 7336
rect 8205 7327 8263 7333
rect 8205 7324 8217 7327
rect 8168 7296 8217 7324
rect 8168 7284 8174 7296
rect 8205 7293 8217 7296
rect 8251 7293 8263 7327
rect 8205 7287 8263 7293
rect 8757 7327 8815 7333
rect 8757 7293 8769 7327
rect 8803 7324 8815 7327
rect 8846 7324 8852 7336
rect 8803 7296 8852 7324
rect 8803 7293 8815 7296
rect 8757 7287 8815 7293
rect 8846 7284 8852 7296
rect 8904 7324 8910 7336
rect 9582 7324 9588 7336
rect 8904 7296 9588 7324
rect 8904 7284 8910 7296
rect 9582 7284 9588 7296
rect 9640 7284 9646 7336
rect 10870 7284 10876 7336
rect 10928 7324 10934 7336
rect 11241 7327 11299 7333
rect 11241 7324 11253 7327
rect 10928 7296 11253 7324
rect 10928 7284 10934 7296
rect 11241 7293 11253 7296
rect 11287 7324 11299 7327
rect 13078 7324 13084 7336
rect 11287 7296 13084 7324
rect 11287 7293 11299 7296
rect 11241 7287 11299 7293
rect 13078 7284 13084 7296
rect 13136 7284 13142 7336
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 14016 7333 14044 7364
rect 14645 7361 14657 7364
rect 14691 7361 14703 7395
rect 14645 7355 14703 7361
rect 14001 7327 14059 7333
rect 14001 7324 14013 7327
rect 13872 7296 14013 7324
rect 13872 7284 13878 7296
rect 14001 7293 14013 7296
rect 14047 7293 14059 7327
rect 14550 7324 14556 7336
rect 14511 7296 14556 7324
rect 14001 7287 14059 7293
rect 14550 7284 14556 7296
rect 14608 7284 14614 7336
rect 2590 7216 2596 7268
rect 2648 7256 2654 7268
rect 2961 7259 3019 7265
rect 2961 7256 2973 7259
rect 2648 7228 2973 7256
rect 2648 7216 2654 7228
rect 2961 7225 2973 7228
rect 3007 7225 3019 7259
rect 2961 7219 3019 7225
rect 3050 7216 3056 7268
rect 3108 7256 3114 7268
rect 14461 7259 14519 7265
rect 3108 7228 3153 7256
rect 3108 7216 3114 7228
rect 14461 7225 14473 7259
rect 14507 7256 14519 7259
rect 14734 7256 14740 7268
rect 14507 7228 14740 7256
rect 14507 7225 14519 7228
rect 14461 7219 14519 7225
rect 14734 7216 14740 7228
rect 14792 7256 14798 7268
rect 14792 7228 15056 7256
rect 14792 7216 14798 7228
rect 3326 7188 3332 7200
rect 2516 7160 3332 7188
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 10686 7148 10692 7200
rect 10744 7188 10750 7200
rect 10781 7191 10839 7197
rect 10781 7188 10793 7191
rect 10744 7160 10793 7188
rect 10744 7148 10750 7160
rect 10781 7157 10793 7160
rect 10827 7188 10839 7191
rect 11333 7191 11391 7197
rect 11333 7188 11345 7191
rect 10827 7160 11345 7188
rect 10827 7157 10839 7160
rect 10781 7151 10839 7157
rect 11333 7157 11345 7160
rect 11379 7157 11391 7191
rect 11333 7151 11391 7157
rect 11422 7148 11428 7200
rect 11480 7188 11486 7200
rect 15028 7197 15056 7228
rect 15013 7191 15071 7197
rect 11480 7160 11525 7188
rect 11480 7148 11486 7160
rect 15013 7157 15025 7191
rect 15059 7157 15071 7191
rect 15013 7151 15071 7157
rect 1104 7098 16100 7120
rect 1104 7046 5980 7098
rect 6032 7046 6044 7098
rect 6096 7046 6108 7098
rect 6160 7046 6172 7098
rect 6224 7046 10979 7098
rect 11031 7046 11043 7098
rect 11095 7046 11107 7098
rect 11159 7046 11171 7098
rect 11223 7046 16100 7098
rect 1104 7024 16100 7046
rect 3326 6944 3332 6996
rect 3384 6984 3390 6996
rect 3881 6987 3939 6993
rect 3881 6984 3893 6987
rect 3384 6956 3893 6984
rect 3384 6944 3390 6956
rect 3881 6953 3893 6956
rect 3927 6953 3939 6987
rect 3881 6947 3939 6953
rect 3970 6944 3976 6996
rect 4028 6984 4034 6996
rect 4065 6987 4123 6993
rect 4065 6984 4077 6987
rect 4028 6956 4077 6984
rect 4028 6944 4034 6956
rect 4065 6953 4077 6956
rect 4111 6953 4123 6987
rect 6546 6984 6552 6996
rect 6507 6956 6552 6984
rect 4065 6947 4123 6953
rect 4080 6916 4108 6947
rect 6546 6944 6552 6956
rect 6604 6944 6610 6996
rect 4080 6888 4200 6916
rect 4062 6851 4120 6857
rect 4062 6817 4074 6851
rect 4108 6817 4120 6851
rect 4172 6848 4200 6888
rect 5074 6876 5080 6928
rect 5132 6916 5138 6928
rect 5169 6919 5227 6925
rect 5169 6916 5181 6919
rect 5132 6888 5181 6916
rect 5132 6876 5138 6888
rect 5169 6885 5181 6888
rect 5215 6885 5227 6919
rect 5813 6919 5871 6925
rect 5813 6916 5825 6919
rect 5169 6879 5227 6885
rect 5644 6888 5825 6916
rect 4617 6851 4675 6857
rect 4617 6848 4629 6851
rect 4172 6820 4629 6848
rect 4062 6811 4120 6817
rect 4617 6817 4629 6820
rect 4663 6817 4675 6851
rect 4617 6811 4675 6817
rect 4709 6851 4767 6857
rect 4709 6817 4721 6851
rect 4755 6817 4767 6851
rect 4709 6811 4767 6817
rect 3878 6672 3884 6724
rect 3936 6712 3942 6724
rect 4080 6712 4108 6811
rect 4522 6780 4528 6792
rect 4483 6752 4528 6780
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 4724 6712 4752 6811
rect 4798 6808 4804 6860
rect 4856 6848 4862 6860
rect 4893 6851 4951 6857
rect 4893 6848 4905 6851
rect 4856 6820 4905 6848
rect 4856 6808 4862 6820
rect 4893 6817 4905 6820
rect 4939 6817 4951 6851
rect 4893 6811 4951 6817
rect 4982 6808 4988 6860
rect 5040 6848 5046 6860
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 5040 6820 5365 6848
rect 5040 6808 5046 6820
rect 5353 6817 5365 6820
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6848 5503 6851
rect 5534 6848 5540 6860
rect 5491 6820 5540 6848
rect 5491 6817 5503 6820
rect 5445 6811 5503 6817
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5644 6780 5672 6888
rect 5813 6885 5825 6888
rect 5859 6916 5871 6919
rect 9582 6916 9588 6928
rect 5859 6888 6316 6916
rect 5859 6885 5871 6888
rect 5813 6879 5871 6885
rect 5905 6851 5963 6857
rect 5905 6848 5917 6851
rect 5123 6752 5672 6780
rect 5736 6820 5917 6848
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 5166 6712 5172 6724
rect 3936 6684 4752 6712
rect 5127 6684 5172 6712
rect 3936 6672 3942 6684
rect 5166 6672 5172 6684
rect 5224 6672 5230 6724
rect 4433 6647 4491 6653
rect 4433 6613 4445 6647
rect 4479 6644 4491 6647
rect 5736 6644 5764 6820
rect 5905 6817 5917 6820
rect 5951 6848 5963 6851
rect 6178 6848 6184 6860
rect 5951 6820 6184 6848
rect 5951 6817 5963 6820
rect 5905 6811 5963 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 6288 6857 6316 6888
rect 6748 6888 6960 6916
rect 9543 6888 9588 6916
rect 6273 6851 6331 6857
rect 6273 6817 6285 6851
rect 6319 6817 6331 6851
rect 6273 6811 6331 6817
rect 6748 6792 6776 6888
rect 6825 6851 6883 6857
rect 6825 6817 6837 6851
rect 6871 6817 6883 6851
rect 6932 6848 6960 6888
rect 9582 6876 9588 6888
rect 9640 6876 9646 6928
rect 10686 6916 10692 6928
rect 10647 6888 10692 6916
rect 10686 6876 10692 6888
rect 10744 6876 10750 6928
rect 7193 6851 7251 6857
rect 7193 6848 7205 6851
rect 6932 6820 7205 6848
rect 6825 6811 6883 6817
rect 7193 6817 7205 6820
rect 7239 6848 7251 6851
rect 7285 6851 7343 6857
rect 7285 6848 7297 6851
rect 7239 6820 7297 6848
rect 7239 6817 7251 6820
rect 7193 6811 7251 6817
rect 7285 6817 7297 6820
rect 7331 6817 7343 6851
rect 7285 6811 7343 6817
rect 9769 6851 9827 6857
rect 9769 6817 9781 6851
rect 9815 6817 9827 6851
rect 9769 6811 9827 6817
rect 10229 6851 10287 6857
rect 10229 6817 10241 6851
rect 10275 6848 10287 6851
rect 10410 6848 10416 6860
rect 10275 6820 10416 6848
rect 10275 6817 10287 6820
rect 10229 6811 10287 6817
rect 6730 6780 6736 6792
rect 6691 6752 6736 6780
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 6840 6780 6868 6811
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 6840 6752 7113 6780
rect 7101 6749 7113 6752
rect 7147 6749 7159 6783
rect 9784 6780 9812 6811
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 10781 6851 10839 6857
rect 10781 6817 10793 6851
rect 10827 6848 10839 6851
rect 10870 6848 10876 6860
rect 10827 6820 10876 6848
rect 10827 6817 10839 6820
rect 10781 6811 10839 6817
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 11241 6851 11299 6857
rect 11241 6817 11253 6851
rect 11287 6848 11299 6851
rect 11422 6848 11428 6860
rect 11287 6820 11428 6848
rect 11287 6817 11299 6820
rect 11241 6811 11299 6817
rect 11422 6808 11428 6820
rect 11480 6808 11486 6860
rect 11698 6808 11704 6860
rect 11756 6848 11762 6860
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 11756 6820 11989 6848
rect 11756 6808 11762 6820
rect 11977 6817 11989 6820
rect 12023 6817 12035 6851
rect 13170 6848 13176 6860
rect 11977 6811 12035 6817
rect 12084 6820 12940 6848
rect 13131 6820 13176 6848
rect 11333 6783 11391 6789
rect 11333 6780 11345 6783
rect 9784 6752 11345 6780
rect 7101 6743 7159 6749
rect 11333 6749 11345 6752
rect 11379 6780 11391 6783
rect 12084 6780 12112 6820
rect 12912 6792 12940 6820
rect 13170 6808 13176 6820
rect 13228 6808 13234 6860
rect 11379 6752 12112 6780
rect 12253 6783 12311 6789
rect 11379 6749 11391 6752
rect 11333 6743 11391 6749
rect 12253 6749 12265 6783
rect 12299 6780 12311 6783
rect 12342 6780 12348 6792
rect 12299 6752 12348 6780
rect 12299 6749 12311 6752
rect 12253 6743 12311 6749
rect 6457 6715 6515 6721
rect 6457 6681 6469 6715
rect 6503 6712 6515 6715
rect 6822 6712 6828 6724
rect 6503 6684 6828 6712
rect 6503 6681 6515 6684
rect 6457 6675 6515 6681
rect 6822 6672 6828 6684
rect 6880 6672 6886 6724
rect 7116 6712 7144 6743
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 12894 6780 12900 6792
rect 12855 6752 12900 6780
rect 12894 6740 12900 6752
rect 12952 6740 12958 6792
rect 7742 6712 7748 6724
rect 7116 6684 7748 6712
rect 7742 6672 7748 6684
rect 7800 6672 7806 6724
rect 4479 6616 5764 6644
rect 7377 6647 7435 6653
rect 4479 6613 4491 6616
rect 4433 6607 4491 6613
rect 7377 6613 7389 6647
rect 7423 6644 7435 6647
rect 7558 6644 7564 6656
rect 7423 6616 7564 6644
rect 7423 6613 7435 6616
rect 7377 6607 7435 6613
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 1104 6554 16100 6576
rect 1104 6502 3481 6554
rect 3533 6502 3545 6554
rect 3597 6502 3609 6554
rect 3661 6502 3673 6554
rect 3725 6502 8480 6554
rect 8532 6502 8544 6554
rect 8596 6502 8608 6554
rect 8660 6502 8672 6554
rect 8724 6502 13478 6554
rect 13530 6502 13542 6554
rect 13594 6502 13606 6554
rect 13658 6502 13670 6554
rect 13722 6502 16100 6554
rect 1104 6480 16100 6502
rect 4065 6443 4123 6449
rect 4065 6409 4077 6443
rect 4111 6440 4123 6443
rect 4522 6440 4528 6452
rect 4111 6412 4528 6440
rect 4111 6409 4123 6412
rect 4065 6403 4123 6409
rect 4522 6400 4528 6412
rect 4580 6400 4586 6452
rect 4893 6443 4951 6449
rect 4893 6409 4905 6443
rect 4939 6440 4951 6443
rect 5074 6440 5080 6452
rect 4939 6412 5080 6440
rect 4939 6409 4951 6412
rect 4893 6403 4951 6409
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 5718 6440 5724 6452
rect 5552 6412 5724 6440
rect 5552 6372 5580 6412
rect 5718 6400 5724 6412
rect 5776 6400 5782 6452
rect 6178 6400 6184 6452
rect 6236 6440 6242 6452
rect 7009 6443 7067 6449
rect 7009 6440 7021 6443
rect 6236 6412 7021 6440
rect 6236 6400 6242 6412
rect 7009 6409 7021 6412
rect 7055 6409 7067 6443
rect 7558 6440 7564 6452
rect 7519 6412 7564 6440
rect 7009 6403 7067 6409
rect 7558 6400 7564 6412
rect 7616 6400 7622 6452
rect 7742 6440 7748 6452
rect 7703 6412 7748 6440
rect 7742 6400 7748 6412
rect 7800 6400 7806 6452
rect 5092 6344 5580 6372
rect 3050 6304 3056 6316
rect 2700 6276 3056 6304
rect 1946 6196 1952 6248
rect 2004 6236 2010 6248
rect 2133 6239 2191 6245
rect 2133 6236 2145 6239
rect 2004 6208 2145 6236
rect 2004 6196 2010 6208
rect 2133 6205 2145 6208
rect 2179 6205 2191 6239
rect 2498 6236 2504 6248
rect 2459 6208 2504 6236
rect 2133 6199 2191 6205
rect 2498 6196 2504 6208
rect 2556 6196 2562 6248
rect 2700 6245 2728 6276
rect 3050 6264 3056 6276
rect 3108 6264 3114 6316
rect 5092 6248 5120 6344
rect 5626 6332 5632 6384
rect 5684 6372 5690 6384
rect 5810 6372 5816 6384
rect 5684 6344 5816 6372
rect 5684 6332 5690 6344
rect 5810 6332 5816 6344
rect 5868 6372 5874 6384
rect 7926 6372 7932 6384
rect 5868 6344 6224 6372
rect 5868 6332 5874 6344
rect 5353 6307 5411 6313
rect 5353 6273 5365 6307
rect 5399 6304 5411 6307
rect 6089 6307 6147 6313
rect 6089 6304 6101 6307
rect 5399 6276 6101 6304
rect 5399 6273 5411 6276
rect 5353 6267 5411 6273
rect 6089 6273 6101 6276
rect 6135 6273 6147 6307
rect 6089 6267 6147 6273
rect 2685 6239 2743 6245
rect 2685 6205 2697 6239
rect 2731 6205 2743 6239
rect 2685 6199 2743 6205
rect 2869 6239 2927 6245
rect 2869 6205 2881 6239
rect 2915 6236 2927 6239
rect 3878 6236 3884 6248
rect 2915 6208 3740 6236
rect 3839 6208 3884 6236
rect 2915 6205 2927 6208
rect 2869 6199 2927 6205
rect 2774 6128 2780 6180
rect 2832 6168 2838 6180
rect 3142 6168 3148 6180
rect 2832 6140 3148 6168
rect 2832 6128 2838 6140
rect 3142 6128 3148 6140
rect 3200 6128 3206 6180
rect 3712 6168 3740 6208
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 3970 6196 3976 6248
rect 4028 6236 4034 6248
rect 4065 6239 4123 6245
rect 4065 6236 4077 6239
rect 4028 6208 4077 6236
rect 4028 6196 4034 6208
rect 4065 6205 4077 6208
rect 4111 6205 4123 6239
rect 5074 6236 5080 6248
rect 5035 6208 5080 6236
rect 4065 6199 4123 6205
rect 5074 6196 5080 6208
rect 5132 6196 5138 6248
rect 5261 6239 5319 6245
rect 5261 6205 5273 6239
rect 5307 6205 5319 6239
rect 5442 6236 5448 6248
rect 5403 6208 5448 6236
rect 5261 6199 5319 6205
rect 4246 6168 4252 6180
rect 3712 6140 4252 6168
rect 4246 6128 4252 6140
rect 4304 6128 4310 6180
rect 5276 6168 5304 6199
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 5629 6239 5687 6245
rect 5629 6205 5641 6239
rect 5675 6205 5687 6239
rect 5629 6199 5687 6205
rect 5534 6168 5540 6180
rect 5276 6140 5540 6168
rect 5534 6128 5540 6140
rect 5592 6128 5598 6180
rect 5644 6168 5672 6199
rect 5718 6196 5724 6248
rect 5776 6236 5782 6248
rect 5905 6239 5963 6245
rect 5776 6208 5821 6236
rect 5776 6196 5782 6208
rect 5905 6205 5917 6239
rect 5951 6205 5963 6239
rect 5905 6199 5963 6205
rect 5997 6239 6055 6245
rect 5997 6205 6009 6239
rect 6043 6236 6055 6239
rect 6196 6236 6224 6344
rect 7484 6344 7932 6372
rect 6043 6208 6224 6236
rect 7190 6239 7248 6245
rect 6043 6205 6055 6208
rect 5997 6199 6055 6205
rect 7190 6205 7202 6239
rect 7236 6236 7248 6239
rect 7484 6236 7512 6344
rect 7926 6332 7932 6344
rect 7984 6332 7990 6384
rect 13170 6304 13176 6316
rect 7236 6208 7512 6236
rect 7576 6276 8064 6304
rect 13131 6276 13176 6304
rect 7236 6205 7248 6208
rect 7190 6199 7248 6205
rect 5813 6171 5871 6177
rect 5813 6168 5825 6171
rect 5644 6140 5825 6168
rect 5813 6137 5825 6140
rect 5859 6137 5871 6171
rect 5813 6131 5871 6137
rect 1854 6060 1860 6112
rect 1912 6100 1918 6112
rect 1949 6103 2007 6109
rect 1949 6100 1961 6103
rect 1912 6072 1961 6100
rect 1912 6060 1918 6072
rect 1949 6069 1961 6072
rect 1995 6069 2007 6103
rect 1949 6063 2007 6069
rect 2866 6060 2872 6112
rect 2924 6100 2930 6112
rect 3053 6103 3111 6109
rect 3053 6100 3065 6103
rect 2924 6072 3065 6100
rect 2924 6060 2930 6072
rect 3053 6069 3065 6072
rect 3099 6069 3111 6103
rect 5552 6100 5580 6128
rect 5920 6100 5948 6199
rect 5552 6072 5948 6100
rect 7193 6103 7251 6109
rect 3053 6063 3111 6069
rect 7193 6069 7205 6103
rect 7239 6100 7251 6103
rect 7576 6100 7604 6276
rect 8036 6245 8064 6276
rect 13170 6264 13176 6276
rect 13228 6264 13234 6316
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6205 7711 6239
rect 7653 6199 7711 6205
rect 8021 6239 8079 6245
rect 8021 6205 8033 6239
rect 8067 6236 8079 6239
rect 8110 6236 8116 6248
rect 8067 6208 8116 6236
rect 8067 6205 8079 6208
rect 8021 6199 8079 6205
rect 7668 6168 7696 6199
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 8297 6239 8355 6245
rect 8297 6205 8309 6239
rect 8343 6205 8355 6239
rect 9582 6236 9588 6248
rect 9543 6208 9588 6236
rect 8297 6199 8355 6205
rect 7745 6171 7803 6177
rect 7745 6168 7757 6171
rect 7668 6140 7757 6168
rect 7745 6137 7757 6140
rect 7791 6168 7803 6171
rect 8205 6171 8263 6177
rect 8205 6168 8217 6171
rect 7791 6140 8217 6168
rect 7791 6137 7803 6140
rect 7745 6131 7803 6137
rect 8205 6137 8217 6140
rect 8251 6137 8263 6171
rect 8205 6131 8263 6137
rect 7926 6100 7932 6112
rect 7239 6072 7604 6100
rect 7887 6072 7932 6100
rect 7239 6069 7251 6072
rect 7193 6063 7251 6069
rect 7926 6060 7932 6072
rect 7984 6100 7990 6112
rect 8312 6100 8340 6199
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 11698 6236 11704 6248
rect 11659 6208 11704 6236
rect 11698 6196 11704 6208
rect 11756 6196 11762 6248
rect 12069 6239 12127 6245
rect 12069 6205 12081 6239
rect 12115 6236 12127 6239
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 12115 6208 12173 6236
rect 12115 6205 12127 6208
rect 12069 6199 12127 6205
rect 12161 6205 12173 6208
rect 12207 6205 12219 6239
rect 12894 6236 12900 6248
rect 12807 6208 12900 6236
rect 12161 6199 12219 6205
rect 12894 6196 12900 6208
rect 12952 6236 12958 6248
rect 13633 6239 13691 6245
rect 13633 6236 13645 6239
rect 12952 6208 13645 6236
rect 12952 6196 12958 6208
rect 13633 6205 13645 6208
rect 13679 6205 13691 6239
rect 13633 6199 13691 6205
rect 11885 6171 11943 6177
rect 11885 6137 11897 6171
rect 11931 6168 11943 6171
rect 12342 6168 12348 6180
rect 11931 6140 12348 6168
rect 11931 6137 11943 6140
rect 11885 6131 11943 6137
rect 12342 6128 12348 6140
rect 12400 6128 12406 6180
rect 13078 6168 13084 6180
rect 13039 6140 13084 6168
rect 13078 6128 13084 6140
rect 13136 6128 13142 6180
rect 7984 6072 8340 6100
rect 9769 6103 9827 6109
rect 7984 6060 7990 6072
rect 9769 6069 9781 6103
rect 9815 6100 9827 6103
rect 9858 6100 9864 6112
rect 9815 6072 9864 6100
rect 9815 6069 9827 6072
rect 9769 6063 9827 6069
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 13814 6100 13820 6112
rect 13775 6072 13820 6100
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 1104 6010 16100 6032
rect 1104 5958 5980 6010
rect 6032 5958 6044 6010
rect 6096 5958 6108 6010
rect 6160 5958 6172 6010
rect 6224 5958 10979 6010
rect 11031 5958 11043 6010
rect 11095 5958 11107 6010
rect 11159 5958 11171 6010
rect 11223 5958 16100 6010
rect 1104 5936 16100 5958
rect 1397 5899 1455 5905
rect 1397 5865 1409 5899
rect 1443 5896 1455 5899
rect 2774 5896 2780 5908
rect 1443 5868 2780 5896
rect 1443 5865 1455 5868
rect 1397 5859 1455 5865
rect 2774 5856 2780 5868
rect 2832 5856 2838 5908
rect 6730 5856 6736 5908
rect 6788 5896 6794 5908
rect 6825 5899 6883 5905
rect 6825 5896 6837 5899
rect 6788 5868 6837 5896
rect 6788 5856 6794 5868
rect 6825 5865 6837 5868
rect 6871 5865 6883 5899
rect 6825 5859 6883 5865
rect 9125 5899 9183 5905
rect 9125 5865 9137 5899
rect 9171 5865 9183 5899
rect 9125 5859 9183 5865
rect 1854 5788 1860 5840
rect 1912 5788 1918 5840
rect 2866 5828 2872 5840
rect 2827 5800 2872 5828
rect 2866 5788 2872 5800
rect 2924 5788 2930 5840
rect 3234 5788 3240 5840
rect 3292 5828 3298 5840
rect 3970 5828 3976 5840
rect 3292 5800 3976 5828
rect 3292 5788 3298 5800
rect 3970 5788 3976 5800
rect 4028 5828 4034 5840
rect 4157 5831 4215 5837
rect 4157 5828 4169 5831
rect 4028 5800 4169 5828
rect 4028 5788 4034 5800
rect 4157 5797 4169 5800
rect 4203 5797 4215 5831
rect 4157 5791 4215 5797
rect 5626 5788 5632 5840
rect 5684 5828 5690 5840
rect 6457 5831 6515 5837
rect 6457 5828 6469 5831
rect 5684 5800 6469 5828
rect 5684 5788 5690 5800
rect 6457 5797 6469 5800
rect 6503 5797 6515 5831
rect 6457 5791 6515 5797
rect 8110 5788 8116 5840
rect 8168 5828 8174 5840
rect 8573 5831 8631 5837
rect 8573 5828 8585 5831
rect 8168 5800 8585 5828
rect 8168 5788 8174 5800
rect 8573 5797 8585 5800
rect 8619 5828 8631 5831
rect 9140 5828 9168 5859
rect 8619 5800 9168 5828
rect 8619 5797 8631 5800
rect 8573 5791 8631 5797
rect 9858 5788 9864 5840
rect 9916 5788 9922 5840
rect 3786 5720 3792 5772
rect 3844 5760 3850 5772
rect 3881 5763 3939 5769
rect 3881 5760 3893 5763
rect 3844 5732 3893 5760
rect 3844 5720 3850 5732
rect 3881 5729 3893 5732
rect 3927 5729 3939 5763
rect 3881 5723 3939 5729
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5729 4123 5763
rect 4246 5760 4252 5772
rect 4207 5732 4252 5760
rect 4065 5723 4123 5729
rect 1670 5652 1676 5704
rect 1728 5692 1734 5704
rect 3145 5695 3203 5701
rect 3145 5692 3157 5695
rect 1728 5664 3157 5692
rect 1728 5652 1734 5664
rect 3145 5661 3157 5664
rect 3191 5661 3203 5695
rect 3145 5655 3203 5661
rect 3160 5624 3188 5655
rect 3970 5652 3976 5704
rect 4028 5692 4034 5704
rect 4080 5692 4108 5723
rect 4246 5720 4252 5732
rect 4304 5720 4310 5772
rect 6270 5760 6276 5772
rect 6231 5732 6276 5760
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 6549 5763 6607 5769
rect 6549 5760 6561 5763
rect 6472 5732 6561 5760
rect 6472 5704 6500 5732
rect 6549 5729 6561 5732
rect 6595 5729 6607 5763
rect 6549 5723 6607 5729
rect 6641 5763 6699 5769
rect 6641 5729 6653 5763
rect 6687 5760 6699 5763
rect 6730 5760 6736 5772
rect 6687 5732 6736 5760
rect 6687 5729 6699 5732
rect 6641 5723 6699 5729
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 8294 5760 8300 5772
rect 8255 5732 8300 5760
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 8481 5763 8539 5769
rect 8481 5729 8493 5763
rect 8527 5729 8539 5763
rect 8481 5723 8539 5729
rect 8665 5763 8723 5769
rect 8665 5729 8677 5763
rect 8711 5729 8723 5763
rect 8665 5723 8723 5729
rect 4028 5664 4108 5692
rect 4028 5652 4034 5664
rect 6454 5652 6460 5704
rect 6512 5652 6518 5704
rect 7926 5652 7932 5704
rect 7984 5692 7990 5704
rect 8202 5692 8208 5704
rect 7984 5664 8208 5692
rect 7984 5652 7990 5664
rect 8202 5652 8208 5664
rect 8260 5692 8266 5704
rect 8496 5692 8524 5723
rect 8260 5664 8524 5692
rect 8260 5652 8266 5664
rect 4982 5624 4988 5636
rect 3160 5596 4988 5624
rect 4982 5584 4988 5596
rect 5040 5584 5046 5636
rect 7006 5584 7012 5636
rect 7064 5624 7070 5636
rect 8680 5624 8708 5723
rect 11054 5720 11060 5772
rect 11112 5760 11118 5772
rect 11241 5763 11299 5769
rect 11241 5760 11253 5763
rect 11112 5732 11253 5760
rect 11112 5720 11118 5732
rect 11241 5729 11253 5732
rect 11287 5729 11299 5763
rect 12342 5760 12348 5772
rect 12303 5732 12348 5760
rect 11241 5723 11299 5729
rect 12342 5720 12348 5732
rect 12400 5720 12406 5772
rect 13814 5720 13820 5772
rect 13872 5760 13878 5772
rect 14461 5763 14519 5769
rect 14461 5760 14473 5763
rect 13872 5732 14473 5760
rect 13872 5720 13878 5732
rect 14461 5729 14473 5732
rect 14507 5729 14519 5763
rect 14461 5723 14519 5729
rect 10597 5695 10655 5701
rect 10597 5692 10609 5695
rect 8864 5664 10609 5692
rect 8864 5633 8892 5664
rect 10597 5661 10609 5664
rect 10643 5661 10655 5695
rect 10597 5655 10655 5661
rect 10873 5695 10931 5701
rect 10873 5661 10885 5695
rect 10919 5692 10931 5695
rect 11330 5692 11336 5704
rect 10919 5664 11336 5692
rect 10919 5661 10931 5664
rect 10873 5655 10931 5661
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 7064 5596 8708 5624
rect 7064 5584 7070 5596
rect 4433 5559 4491 5565
rect 4433 5525 4445 5559
rect 4479 5556 4491 5559
rect 4706 5556 4712 5568
rect 4479 5528 4712 5556
rect 4479 5525 4491 5528
rect 4433 5519 4491 5525
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 8680 5556 8708 5596
rect 8849 5627 8907 5633
rect 8849 5593 8861 5627
rect 8895 5593 8907 5627
rect 12161 5627 12219 5633
rect 12161 5624 12173 5627
rect 8849 5587 8907 5593
rect 10796 5596 12173 5624
rect 10796 5568 10824 5596
rect 12161 5593 12173 5596
rect 12207 5624 12219 5627
rect 12526 5624 12532 5636
rect 12207 5596 12532 5624
rect 12207 5593 12219 5596
rect 12161 5587 12219 5593
rect 12526 5584 12532 5596
rect 12584 5584 12590 5636
rect 9398 5556 9404 5568
rect 8680 5528 9404 5556
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 10778 5516 10784 5568
rect 10836 5516 10842 5568
rect 11238 5556 11244 5568
rect 11199 5528 11244 5556
rect 11238 5516 11244 5528
rect 11296 5516 11302 5568
rect 14458 5556 14464 5568
rect 14419 5528 14464 5556
rect 14458 5516 14464 5528
rect 14516 5516 14522 5568
rect 1104 5466 16100 5488
rect 1104 5414 3481 5466
rect 3533 5414 3545 5466
rect 3597 5414 3609 5466
rect 3661 5414 3673 5466
rect 3725 5414 8480 5466
rect 8532 5414 8544 5466
rect 8596 5414 8608 5466
rect 8660 5414 8672 5466
rect 8724 5414 13478 5466
rect 13530 5414 13542 5466
rect 13594 5414 13606 5466
rect 13658 5414 13670 5466
rect 13722 5414 16100 5466
rect 1104 5392 16100 5414
rect 3234 5352 3240 5364
rect 3195 5324 3240 5352
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 5353 5355 5411 5361
rect 5353 5321 5365 5355
rect 5399 5352 5411 5355
rect 6270 5352 6276 5364
rect 5399 5324 6276 5352
rect 5399 5321 5411 5324
rect 5353 5315 5411 5321
rect 6270 5312 6276 5324
rect 6328 5352 6334 5364
rect 6457 5355 6515 5361
rect 6457 5352 6469 5355
rect 6328 5324 6469 5352
rect 6328 5312 6334 5324
rect 6457 5321 6469 5324
rect 6503 5321 6515 5355
rect 6457 5315 6515 5321
rect 9030 5312 9036 5364
rect 9088 5352 9094 5364
rect 11238 5352 11244 5364
rect 9088 5324 11244 5352
rect 9088 5312 9094 5324
rect 5166 5244 5172 5296
rect 5224 5284 5230 5296
rect 7929 5287 7987 5293
rect 7929 5284 7941 5287
rect 5224 5256 7941 5284
rect 5224 5244 5230 5256
rect 7929 5253 7941 5256
rect 7975 5284 7987 5287
rect 8754 5284 8760 5296
rect 7975 5256 8760 5284
rect 7975 5253 7987 5256
rect 7929 5247 7987 5253
rect 8754 5244 8760 5256
rect 8812 5244 8818 5296
rect 10318 5244 10324 5296
rect 10376 5284 10382 5296
rect 10965 5287 11023 5293
rect 10965 5284 10977 5287
rect 10376 5256 10977 5284
rect 10376 5244 10382 5256
rect 10965 5253 10977 5256
rect 11011 5253 11023 5287
rect 10965 5247 11023 5253
rect 4706 5216 4712 5228
rect 4667 5188 4712 5216
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 4982 5216 4988 5228
rect 4943 5188 4988 5216
rect 4982 5176 4988 5188
rect 5040 5176 5046 5228
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 7009 5219 7067 5225
rect 7009 5216 7021 5219
rect 6788 5188 7021 5216
rect 6788 5176 6794 5188
rect 7009 5185 7021 5188
rect 7055 5216 7067 5219
rect 9306 5216 9312 5228
rect 7055 5188 9312 5216
rect 7055 5185 7067 5188
rect 7009 5179 7067 5185
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 10870 5216 10876 5228
rect 9416 5188 10876 5216
rect 9416 5160 9444 5188
rect 10870 5176 10876 5188
rect 10928 5176 10934 5228
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5117 5319 5151
rect 5261 5111 5319 5117
rect 5813 5151 5871 5157
rect 5813 5117 5825 5151
rect 5859 5117 5871 5151
rect 5813 5111 5871 5117
rect 4154 5040 4160 5092
rect 4212 5040 4218 5092
rect 5276 5080 5304 5111
rect 5626 5080 5632 5092
rect 5276 5052 5632 5080
rect 5626 5040 5632 5052
rect 5684 5080 5690 5092
rect 5828 5080 5856 5111
rect 6454 5108 6460 5160
rect 6512 5148 6518 5160
rect 6638 5151 6696 5157
rect 6638 5148 6650 5151
rect 6512 5120 6650 5148
rect 6512 5108 6518 5120
rect 6638 5117 6650 5120
rect 6684 5148 6696 5151
rect 7101 5151 7159 5157
rect 7101 5148 7113 5151
rect 6684 5120 7113 5148
rect 6684 5117 6696 5120
rect 6638 5111 6696 5117
rect 7101 5117 7113 5120
rect 7147 5117 7159 5151
rect 7101 5111 7159 5117
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5148 7987 5151
rect 8205 5151 8263 5157
rect 8205 5148 8217 5151
rect 7975 5120 8217 5148
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 8205 5117 8217 5120
rect 8251 5117 8263 5151
rect 8205 5111 8263 5117
rect 5684 5052 5856 5080
rect 7116 5080 7144 5111
rect 8294 5108 8300 5160
rect 8352 5148 8358 5160
rect 9030 5148 9036 5160
rect 8352 5120 9036 5148
rect 8352 5108 8358 5120
rect 9030 5108 9036 5120
rect 9088 5108 9094 5160
rect 9398 5148 9404 5160
rect 9359 5120 9404 5148
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 9582 5108 9588 5160
rect 9640 5148 9646 5160
rect 9858 5148 9864 5160
rect 9640 5120 9864 5148
rect 9640 5108 9646 5120
rect 9858 5108 9864 5120
rect 9916 5148 9922 5160
rect 10505 5151 10563 5157
rect 10505 5148 10517 5151
rect 9916 5120 10517 5148
rect 9916 5108 9922 5120
rect 10505 5117 10517 5120
rect 10551 5148 10563 5151
rect 10778 5148 10784 5160
rect 10551 5120 10784 5148
rect 10551 5117 10563 5120
rect 10505 5111 10563 5117
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 9122 5080 9128 5092
rect 7116 5052 9128 5080
rect 5684 5040 5690 5052
rect 9122 5040 9128 5052
rect 9180 5080 9186 5092
rect 9217 5083 9275 5089
rect 9217 5080 9229 5083
rect 9180 5052 9229 5080
rect 9180 5040 9186 5052
rect 9217 5049 9229 5052
rect 9263 5049 9275 5083
rect 9217 5043 9275 5049
rect 9306 5040 9312 5092
rect 9364 5080 9370 5092
rect 9364 5052 9409 5080
rect 9364 5040 9370 5052
rect 5534 5012 5540 5024
rect 5495 4984 5540 5012
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 5721 5015 5779 5021
rect 5721 4981 5733 5015
rect 5767 5012 5779 5015
rect 6270 5012 6276 5024
rect 5767 4984 6276 5012
rect 5767 4981 5779 4984
rect 5721 4975 5779 4981
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6641 5015 6699 5021
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 6730 5012 6736 5024
rect 6687 4984 6736 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 6730 4972 6736 4984
rect 6788 4972 6794 5024
rect 7926 4972 7932 5024
rect 7984 5012 7990 5024
rect 8021 5015 8079 5021
rect 8021 5012 8033 5015
rect 7984 4984 8033 5012
rect 7984 4972 7990 4984
rect 8021 4981 8033 4984
rect 8067 4981 8079 5015
rect 9582 5012 9588 5024
rect 9543 4984 9588 5012
rect 8021 4975 8079 4981
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 10318 5012 10324 5024
rect 10279 4984 10324 5012
rect 10318 4972 10324 4984
rect 10376 4972 10382 5024
rect 11072 5012 11100 5324
rect 11238 5312 11244 5324
rect 11296 5312 11302 5364
rect 15562 5352 15568 5364
rect 12452 5324 15568 5352
rect 12342 5216 12348 5228
rect 12303 5188 12348 5216
rect 12342 5176 12348 5188
rect 12400 5176 12406 5228
rect 11149 5151 11207 5157
rect 11149 5117 11161 5151
rect 11195 5148 11207 5151
rect 11882 5148 11888 5160
rect 11195 5120 11888 5148
rect 11195 5117 11207 5120
rect 11149 5111 11207 5117
rect 11882 5108 11888 5120
rect 11940 5108 11946 5160
rect 12158 5148 12164 5160
rect 12119 5120 12164 5148
rect 12158 5108 12164 5120
rect 12216 5108 12222 5160
rect 12452 5157 12480 5324
rect 15562 5312 15568 5324
rect 15620 5312 15626 5364
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 13817 5219 13875 5225
rect 13817 5216 13829 5219
rect 13780 5188 13829 5216
rect 13780 5176 13786 5188
rect 13817 5185 13829 5188
rect 13863 5216 13875 5219
rect 14458 5216 14464 5228
rect 13863 5188 14464 5216
rect 13863 5185 13875 5188
rect 13817 5179 13875 5185
rect 14458 5176 14464 5188
rect 14516 5176 14522 5228
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5117 12495 5151
rect 12437 5111 12495 5117
rect 12526 5108 12532 5160
rect 12584 5148 12590 5160
rect 13170 5148 13176 5160
rect 12584 5120 13176 5148
rect 12584 5108 12590 5120
rect 13170 5108 13176 5120
rect 13228 5108 13234 5160
rect 11241 5083 11299 5089
rect 11241 5049 11253 5083
rect 11287 5080 11299 5083
rect 11422 5080 11428 5092
rect 11287 5052 11428 5080
rect 11287 5049 11299 5052
rect 11241 5043 11299 5049
rect 11422 5040 11428 5052
rect 11480 5040 11486 5092
rect 11517 5083 11575 5089
rect 11517 5049 11529 5083
rect 11563 5080 11575 5083
rect 11606 5080 11612 5092
rect 11563 5052 11612 5080
rect 11563 5049 11575 5052
rect 11517 5043 11575 5049
rect 11606 5040 11612 5052
rect 11664 5040 11670 5092
rect 14090 5080 14096 5092
rect 14051 5052 14096 5080
rect 14090 5040 14096 5052
rect 14148 5040 14154 5092
rect 14182 5040 14188 5092
rect 14240 5080 14246 5092
rect 14240 5052 14582 5080
rect 14240 5040 14246 5052
rect 11333 5015 11391 5021
rect 11333 5012 11345 5015
rect 11072 4984 11345 5012
rect 11333 4981 11345 4984
rect 11379 5012 11391 5015
rect 11698 5012 11704 5024
rect 11379 4984 11704 5012
rect 11379 4981 11391 4984
rect 11333 4975 11391 4981
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 12986 5012 12992 5024
rect 12947 4984 12992 5012
rect 12986 4972 12992 4984
rect 13044 4972 13050 5024
rect 15562 5012 15568 5024
rect 15523 4984 15568 5012
rect 15562 4972 15568 4984
rect 15620 4972 15626 5024
rect 1104 4922 16100 4944
rect 1104 4870 5980 4922
rect 6032 4870 6044 4922
rect 6096 4870 6108 4922
rect 6160 4870 6172 4922
rect 6224 4870 10979 4922
rect 11031 4870 11043 4922
rect 11095 4870 11107 4922
rect 11159 4870 11171 4922
rect 11223 4870 16100 4922
rect 1104 4848 16100 4870
rect 2590 4808 2596 4820
rect 2551 4780 2596 4808
rect 2590 4768 2596 4780
rect 2648 4808 2654 4820
rect 2869 4811 2927 4817
rect 2869 4808 2881 4811
rect 2648 4780 2881 4808
rect 2648 4768 2654 4780
rect 2869 4777 2881 4780
rect 2915 4777 2927 4811
rect 4154 4808 4160 4820
rect 4115 4780 4160 4808
rect 2869 4771 2927 4777
rect 4154 4768 4160 4780
rect 4212 4768 4218 4820
rect 5810 4768 5816 4820
rect 5868 4808 5874 4820
rect 6089 4811 6147 4817
rect 6089 4808 6101 4811
rect 5868 4780 6101 4808
rect 5868 4768 5874 4780
rect 6089 4777 6101 4780
rect 6135 4777 6147 4811
rect 6089 4771 6147 4777
rect 9306 4768 9312 4820
rect 9364 4808 9370 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9364 4780 9413 4808
rect 9364 4768 9370 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 9401 4771 9459 4777
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 11977 4811 12035 4817
rect 9640 4780 10916 4808
rect 9640 4768 9646 4780
rect 2409 4743 2467 4749
rect 2409 4709 2421 4743
rect 2455 4740 2467 4743
rect 2498 4740 2504 4752
rect 2455 4712 2504 4740
rect 2455 4709 2467 4712
rect 2409 4703 2467 4709
rect 2498 4700 2504 4712
rect 2556 4740 2562 4752
rect 3786 4740 3792 4752
rect 2556 4712 3792 4740
rect 2556 4700 2562 4712
rect 3786 4700 3792 4712
rect 3844 4740 3850 4752
rect 4522 4740 4528 4752
rect 3844 4712 4528 4740
rect 3844 4700 3850 4712
rect 4522 4700 4528 4712
rect 4580 4700 4586 4752
rect 4982 4700 4988 4752
rect 5040 4740 5046 4752
rect 5040 4712 6960 4740
rect 5040 4700 5046 4712
rect 6932 4684 6960 4712
rect 7926 4700 7932 4752
rect 7984 4700 7990 4752
rect 10318 4700 10324 4752
rect 10376 4700 10382 4752
rect 10888 4749 10916 4780
rect 11977 4777 11989 4811
rect 12023 4777 12035 4811
rect 14182 4808 14188 4820
rect 14143 4780 14188 4808
rect 11977 4771 12035 4777
rect 10873 4743 10931 4749
rect 10873 4709 10885 4743
rect 10919 4709 10931 4743
rect 10873 4703 10931 4709
rect 10962 4700 10968 4752
rect 11020 4740 11026 4752
rect 11020 4712 11376 4740
rect 11020 4700 11026 4712
rect 1946 4632 1952 4684
rect 2004 4672 2010 4684
rect 2041 4675 2099 4681
rect 2041 4672 2053 4675
rect 2004 4644 2053 4672
rect 2004 4632 2010 4644
rect 2041 4641 2053 4644
rect 2087 4641 2099 4675
rect 2041 4635 2099 4641
rect 2685 4675 2743 4681
rect 2685 4641 2697 4675
rect 2731 4672 2743 4675
rect 2774 4672 2780 4684
rect 2731 4644 2780 4672
rect 2731 4641 2743 4644
rect 2685 4635 2743 4641
rect 2056 4604 2084 4635
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 2961 4675 3019 4681
rect 2961 4641 2973 4675
rect 3007 4672 3019 4675
rect 3050 4672 3056 4684
rect 3007 4644 3056 4672
rect 3007 4641 3019 4644
rect 2961 4635 3019 4641
rect 3050 4632 3056 4644
rect 3108 4632 3114 4684
rect 4341 4675 4399 4681
rect 4341 4641 4353 4675
rect 4387 4641 4399 4675
rect 5442 4672 5448 4684
rect 5403 4644 5448 4672
rect 4341 4635 4399 4641
rect 4356 4604 4384 4635
rect 5442 4632 5448 4644
rect 5500 4632 5506 4684
rect 5626 4632 5632 4684
rect 5684 4672 5690 4684
rect 5997 4675 6055 4681
rect 5997 4672 6009 4675
rect 5684 4644 6009 4672
rect 5684 4632 5690 4644
rect 5997 4641 6009 4644
rect 6043 4641 6055 4675
rect 6914 4672 6920 4684
rect 6827 4644 6920 4672
rect 5997 4635 6055 4641
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 11348 4681 11376 4712
rect 11422 4700 11428 4752
rect 11480 4740 11486 4752
rect 11517 4743 11575 4749
rect 11517 4740 11529 4743
rect 11480 4712 11529 4740
rect 11480 4700 11486 4712
rect 11517 4709 11529 4712
rect 11563 4740 11575 4743
rect 11992 4740 12020 4771
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 11563 4712 12020 4740
rect 11563 4709 11575 4712
rect 11517 4703 11575 4709
rect 12986 4700 12992 4752
rect 13044 4700 13050 4752
rect 13170 4700 13176 4752
rect 13228 4740 13234 4752
rect 13228 4712 14044 4740
rect 13228 4700 13234 4712
rect 11333 4675 11391 4681
rect 11333 4641 11345 4675
rect 11379 4641 11391 4675
rect 11606 4672 11612 4684
rect 11567 4644 11612 4672
rect 11333 4635 11391 4641
rect 5166 4604 5172 4616
rect 2056 4576 5172 4604
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 5350 4604 5356 4616
rect 5311 4576 5356 4604
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 7190 4604 7196 4616
rect 7151 4576 7196 4604
rect 7190 4564 7196 4576
rect 7248 4564 7254 4616
rect 7282 4564 7288 4616
rect 7340 4604 7346 4616
rect 8202 4604 8208 4616
rect 7340 4576 8208 4604
rect 7340 4564 7346 4576
rect 8202 4564 8208 4576
rect 8260 4604 8266 4616
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 8260 4576 8953 4604
rect 8260 4564 8266 4576
rect 8941 4573 8953 4576
rect 8987 4573 8999 4607
rect 11146 4604 11152 4616
rect 11107 4576 11152 4604
rect 8941 4567 8999 4573
rect 11146 4564 11152 4576
rect 11204 4564 11210 4616
rect 11348 4604 11376 4635
rect 11606 4632 11612 4644
rect 11664 4632 11670 4684
rect 11698 4632 11704 4684
rect 11756 4672 11762 4684
rect 11756 4644 11801 4672
rect 11756 4632 11762 4644
rect 13722 4632 13728 4684
rect 13780 4672 13786 4684
rect 14016 4681 14044 4712
rect 15028 4712 15608 4740
rect 14001 4675 14059 4681
rect 13780 4644 13825 4672
rect 13780 4632 13786 4644
rect 14001 4641 14013 4675
rect 14047 4641 14059 4675
rect 14001 4635 14059 4641
rect 14090 4632 14096 4684
rect 14148 4672 14154 4684
rect 15028 4681 15056 4712
rect 15580 4684 15608 4712
rect 14829 4675 14887 4681
rect 14829 4672 14841 4675
rect 14148 4644 14841 4672
rect 14148 4632 14154 4644
rect 12066 4604 12072 4616
rect 11348 4576 12072 4604
rect 12066 4564 12072 4576
rect 12124 4564 12130 4616
rect 13449 4607 13507 4613
rect 13449 4604 13461 4607
rect 12406 4576 13461 4604
rect 8754 4496 8760 4548
rect 8812 4536 8818 4548
rect 9858 4536 9864 4548
rect 8812 4508 9864 4536
rect 8812 4496 8818 4508
rect 9858 4496 9864 4508
rect 9916 4496 9922 4548
rect 11885 4539 11943 4545
rect 11885 4505 11897 4539
rect 11931 4536 11943 4539
rect 12406 4536 12434 4576
rect 13449 4573 13461 4576
rect 13495 4573 13507 4607
rect 13449 4567 13507 4573
rect 11931 4508 12434 4536
rect 14660 4536 14688 4644
rect 14829 4641 14841 4644
rect 14875 4641 14887 4675
rect 14829 4635 14887 4641
rect 15013 4675 15071 4681
rect 15013 4641 15025 4675
rect 15059 4641 15071 4675
rect 15013 4635 15071 4641
rect 15562 4632 15568 4684
rect 15620 4672 15626 4684
rect 15620 4644 15665 4672
rect 15620 4632 15626 4644
rect 15657 4607 15715 4613
rect 15657 4573 15669 4607
rect 15703 4573 15715 4607
rect 15657 4567 15715 4573
rect 15672 4536 15700 4567
rect 15746 4536 15752 4548
rect 14660 4508 15752 4536
rect 11931 4505 11943 4508
rect 11885 4499 11943 4505
rect 15746 4496 15752 4508
rect 15804 4496 15810 4548
rect 2222 4468 2228 4480
rect 2183 4440 2228 4468
rect 2222 4428 2228 4440
rect 2280 4428 2286 4480
rect 2406 4468 2412 4480
rect 2367 4440 2412 4468
rect 2406 4428 2412 4440
rect 2464 4428 2470 4480
rect 4522 4428 4528 4480
rect 4580 4468 4586 4480
rect 8294 4468 8300 4480
rect 4580 4440 8300 4468
rect 4580 4428 4586 4440
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 12066 4428 12072 4480
rect 12124 4468 12130 4480
rect 14553 4471 14611 4477
rect 14553 4468 14565 4471
rect 12124 4440 14565 4468
rect 12124 4428 12130 4440
rect 14553 4437 14565 4440
rect 14599 4437 14611 4471
rect 14553 4431 14611 4437
rect 1104 4378 16100 4400
rect 1104 4326 3481 4378
rect 3533 4326 3545 4378
rect 3597 4326 3609 4378
rect 3661 4326 3673 4378
rect 3725 4326 8480 4378
rect 8532 4326 8544 4378
rect 8596 4326 8608 4378
rect 8660 4326 8672 4378
rect 8724 4326 13478 4378
rect 13530 4326 13542 4378
rect 13594 4326 13606 4378
rect 13658 4326 13670 4378
rect 13722 4326 16100 4378
rect 1104 4304 16100 4326
rect 1660 4267 1718 4273
rect 1660 4233 1672 4267
rect 1706 4264 1718 4267
rect 2406 4264 2412 4276
rect 1706 4236 2412 4264
rect 1706 4233 1718 4236
rect 1660 4227 1718 4233
rect 2406 4224 2412 4236
rect 2464 4224 2470 4276
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 3145 4267 3203 4273
rect 3145 4264 3157 4267
rect 3108 4236 3157 4264
rect 3108 4224 3114 4236
rect 3145 4233 3157 4236
rect 3191 4264 3203 4267
rect 3234 4264 3240 4276
rect 3191 4236 3240 4264
rect 3191 4233 3203 4236
rect 3145 4227 3203 4233
rect 3234 4224 3240 4236
rect 3292 4224 3298 4276
rect 11146 4224 11152 4276
rect 11204 4264 11210 4276
rect 12434 4264 12440 4276
rect 11204 4236 12440 4264
rect 11204 4224 11210 4236
rect 12434 4224 12440 4236
rect 12492 4264 12498 4276
rect 13814 4264 13820 4276
rect 12492 4236 13820 4264
rect 12492 4224 12498 4236
rect 13814 4224 13820 4236
rect 13872 4224 13878 4276
rect 15746 4264 15752 4276
rect 15707 4236 15752 4264
rect 15746 4224 15752 4236
rect 15804 4224 15810 4276
rect 5442 4156 5448 4208
rect 5500 4196 5506 4208
rect 5500 4168 6132 4196
rect 5500 4156 5506 4168
rect 1394 4128 1400 4140
rect 1307 4100 1400 4128
rect 1394 4088 1400 4100
rect 1452 4128 1458 4140
rect 1670 4128 1676 4140
rect 1452 4100 1676 4128
rect 1452 4088 1458 4100
rect 1670 4088 1676 4100
rect 1728 4088 1734 4140
rect 5626 4128 5632 4140
rect 5587 4100 5632 4128
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 5350 4020 5356 4072
rect 5408 4060 5414 4072
rect 6104 4069 6132 4168
rect 11606 4088 11612 4140
rect 11664 4128 11670 4140
rect 11664 4100 12020 4128
rect 11664 4088 11670 4100
rect 11992 4072 12020 4100
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13872 4100 14013 4128
rect 13872 4088 13878 4100
rect 14001 4097 14013 4100
rect 14047 4097 14059 4131
rect 14001 4091 14059 4097
rect 5537 4063 5595 4069
rect 5537 4060 5549 4063
rect 5408 4032 5549 4060
rect 5408 4020 5414 4032
rect 5537 4029 5549 4032
rect 5583 4029 5595 4063
rect 5537 4023 5595 4029
rect 6089 4063 6147 4069
rect 6089 4029 6101 4063
rect 6135 4060 6147 4063
rect 6638 4060 6644 4072
rect 6135 4032 6644 4060
rect 6135 4029 6147 4032
rect 6089 4023 6147 4029
rect 2222 3952 2228 4004
rect 2280 3952 2286 4004
rect 5552 3992 5580 4023
rect 6638 4020 6644 4032
rect 6696 4020 6702 4072
rect 7282 4060 7288 4072
rect 7243 4032 7288 4060
rect 7282 4020 7288 4032
rect 7340 4020 7346 4072
rect 11698 4060 11704 4072
rect 11659 4032 11704 4060
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 11974 4060 11980 4072
rect 11887 4032 11980 4060
rect 11974 4020 11980 4032
rect 12032 4020 12038 4072
rect 12066 4020 12072 4072
rect 12124 4060 12130 4072
rect 12124 4032 12169 4060
rect 12124 4020 12130 4032
rect 6362 3992 6368 4004
rect 5552 3964 6368 3992
rect 6362 3952 6368 3964
rect 6420 3952 6426 4004
rect 9306 3992 9312 4004
rect 6472 3964 9312 3992
rect 6270 3884 6276 3936
rect 6328 3924 6334 3936
rect 6472 3924 6500 3964
rect 9306 3952 9312 3964
rect 9364 3952 9370 4004
rect 11882 3992 11888 4004
rect 11843 3964 11888 3992
rect 11882 3952 11888 3964
rect 11940 3952 11946 4004
rect 14274 3992 14280 4004
rect 14235 3964 14280 3992
rect 14274 3952 14280 3964
rect 14332 3952 14338 4004
rect 14918 3952 14924 4004
rect 14976 3952 14982 4004
rect 6328 3896 6500 3924
rect 6328 3884 6334 3896
rect 6546 3884 6552 3936
rect 6604 3924 6610 3936
rect 7193 3927 7251 3933
rect 7193 3924 7205 3927
rect 6604 3896 7205 3924
rect 6604 3884 6610 3896
rect 7193 3893 7205 3896
rect 7239 3893 7251 3927
rect 7193 3887 7251 3893
rect 12253 3927 12311 3933
rect 12253 3893 12265 3927
rect 12299 3924 12311 3927
rect 13538 3924 13544 3936
rect 12299 3896 13544 3924
rect 12299 3893 12311 3896
rect 12253 3887 12311 3893
rect 13538 3884 13544 3896
rect 13596 3884 13602 3936
rect 1104 3834 16100 3856
rect 1104 3782 5980 3834
rect 6032 3782 6044 3834
rect 6096 3782 6108 3834
rect 6160 3782 6172 3834
rect 6224 3782 10979 3834
rect 11031 3782 11043 3834
rect 11095 3782 11107 3834
rect 11159 3782 11171 3834
rect 11223 3782 16100 3834
rect 1104 3760 16100 3782
rect 3234 3680 3240 3732
rect 3292 3720 3298 3732
rect 4249 3723 4307 3729
rect 4249 3720 4261 3723
rect 3292 3692 4261 3720
rect 3292 3680 3298 3692
rect 4249 3689 4261 3692
rect 4295 3689 4307 3723
rect 7006 3720 7012 3732
rect 4249 3683 4307 3689
rect 6288 3692 7012 3720
rect 3970 3652 3976 3664
rect 3931 3624 3976 3652
rect 3970 3612 3976 3624
rect 4028 3612 4034 3664
rect 4077 3624 4292 3652
rect 3326 3544 3332 3596
rect 3384 3584 3390 3596
rect 4077 3584 4105 3624
rect 4264 3596 4292 3624
rect 3384 3556 4105 3584
rect 4157 3587 4215 3593
rect 3384 3544 3390 3556
rect 4157 3553 4169 3587
rect 4203 3553 4215 3587
rect 4157 3547 4215 3553
rect 4172 3516 4200 3547
rect 4246 3544 4252 3596
rect 4304 3584 4310 3596
rect 6288 3593 6316 3692
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 8573 3723 8631 3729
rect 8573 3720 8585 3723
rect 7116 3692 8585 3720
rect 6362 3612 6368 3664
rect 6420 3652 6426 3664
rect 7116 3652 7144 3692
rect 8573 3689 8585 3692
rect 8619 3689 8631 3723
rect 8573 3683 8631 3689
rect 11974 3680 11980 3732
rect 12032 3720 12038 3732
rect 12069 3723 12127 3729
rect 12069 3720 12081 3723
rect 12032 3692 12081 3720
rect 12032 3680 12038 3692
rect 12069 3689 12081 3692
rect 12115 3689 12127 3723
rect 12069 3683 12127 3689
rect 9214 3652 9220 3664
rect 6420 3624 7144 3652
rect 8680 3624 9220 3652
rect 6420 3612 6426 3624
rect 4341 3587 4399 3593
rect 4341 3584 4353 3587
rect 4304 3556 4353 3584
rect 4304 3544 4310 3556
rect 4341 3553 4353 3556
rect 4387 3584 4399 3587
rect 6273 3587 6331 3593
rect 6273 3584 6285 3587
rect 4387 3556 6285 3584
rect 4387 3553 4399 3556
rect 4341 3547 4399 3553
rect 6273 3553 6285 3556
rect 6319 3553 6331 3587
rect 6454 3584 6460 3596
rect 6415 3556 6460 3584
rect 6273 3547 6331 3553
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 6822 3584 6828 3596
rect 6783 3556 6828 3584
rect 6822 3544 6828 3556
rect 6880 3544 6886 3596
rect 7006 3544 7012 3596
rect 7064 3584 7070 3596
rect 8680 3593 8708 3624
rect 9214 3612 9220 3624
rect 9272 3652 9278 3664
rect 9401 3655 9459 3661
rect 9401 3652 9413 3655
rect 9272 3624 9413 3652
rect 9272 3612 9278 3624
rect 9401 3621 9413 3624
rect 9447 3621 9459 3655
rect 9401 3615 9459 3621
rect 11514 3612 11520 3664
rect 11572 3612 11578 3664
rect 12526 3612 12532 3664
rect 12584 3612 12590 3664
rect 13538 3652 13544 3664
rect 13499 3624 13544 3652
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 7469 3587 7527 3593
rect 7469 3584 7481 3587
rect 7064 3556 7481 3584
rect 7064 3544 7070 3556
rect 7469 3553 7481 3556
rect 7515 3553 7527 3587
rect 7469 3547 7527 3553
rect 8665 3587 8723 3593
rect 8665 3553 8677 3587
rect 8711 3553 8723 3587
rect 8665 3547 8723 3553
rect 9030 3544 9036 3596
rect 9088 3584 9094 3596
rect 9125 3587 9183 3593
rect 9125 3584 9137 3587
rect 9088 3556 9137 3584
rect 9088 3544 9094 3556
rect 9125 3553 9137 3556
rect 9171 3553 9183 3587
rect 9306 3584 9312 3596
rect 9267 3556 9312 3584
rect 9125 3547 9183 3553
rect 9306 3544 9312 3556
rect 9364 3544 9370 3596
rect 9490 3584 9496 3596
rect 9451 3556 9496 3584
rect 9490 3544 9496 3556
rect 9548 3544 9554 3596
rect 9858 3544 9864 3596
rect 9916 3584 9922 3596
rect 10042 3584 10048 3596
rect 9916 3556 10048 3584
rect 9916 3544 9922 3556
rect 10042 3544 10048 3556
rect 10100 3544 10106 3596
rect 13814 3544 13820 3596
rect 13872 3584 13878 3596
rect 13872 3556 13917 3584
rect 13872 3544 13878 3556
rect 4172 3488 4292 3516
rect 4264 3460 4292 3488
rect 6362 3476 6368 3528
rect 6420 3516 6426 3528
rect 6549 3519 6607 3525
rect 6549 3516 6561 3519
rect 6420 3488 6561 3516
rect 6420 3476 6426 3488
rect 6549 3485 6561 3488
rect 6595 3485 6607 3519
rect 6549 3479 6607 3485
rect 6638 3476 6644 3528
rect 6696 3516 6702 3528
rect 6696 3488 6741 3516
rect 6696 3476 6702 3488
rect 7098 3476 7104 3528
rect 7156 3516 7162 3528
rect 7281 3519 7339 3525
rect 7281 3516 7293 3519
rect 7156 3488 7293 3516
rect 7156 3476 7162 3488
rect 7281 3485 7293 3488
rect 7327 3485 7339 3519
rect 7281 3479 7339 3485
rect 7374 3476 7380 3528
rect 7432 3516 7438 3528
rect 7561 3519 7619 3525
rect 7432 3488 7477 3516
rect 7432 3476 7438 3488
rect 7561 3485 7573 3519
rect 7607 3485 7619 3519
rect 7561 3479 7619 3485
rect 4246 3408 4252 3460
rect 4304 3408 4310 3460
rect 7190 3448 7196 3460
rect 6840 3420 7196 3448
rect 4525 3383 4583 3389
rect 4525 3349 4537 3383
rect 4571 3380 4583 3383
rect 6840 3380 6868 3420
rect 7190 3408 7196 3420
rect 7248 3448 7254 3460
rect 7576 3448 7604 3479
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 10229 3519 10287 3525
rect 10229 3516 10241 3519
rect 7708 3488 10241 3516
rect 7708 3476 7714 3488
rect 10229 3485 10241 3488
rect 10275 3485 10287 3519
rect 10229 3479 10287 3485
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3516 10563 3519
rect 11146 3516 11152 3528
rect 10551 3488 11152 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 7248 3420 7604 3448
rect 7248 3408 7254 3420
rect 7006 3380 7012 3392
rect 4571 3352 6868 3380
rect 6967 3352 7012 3380
rect 4571 3349 4583 3352
rect 4525 3343 4583 3349
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 7101 3383 7159 3389
rect 7101 3349 7113 3383
rect 7147 3380 7159 3383
rect 7282 3380 7288 3392
rect 7147 3352 7288 3380
rect 7147 3349 7159 3352
rect 7101 3343 7159 3349
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 9674 3380 9680 3392
rect 9635 3352 9680 3380
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 9766 3340 9772 3392
rect 9824 3380 9830 3392
rect 9861 3383 9919 3389
rect 9861 3380 9873 3383
rect 9824 3352 9873 3380
rect 9824 3340 9830 3352
rect 9861 3349 9873 3352
rect 9907 3349 9919 3383
rect 10244 3380 10272 3479
rect 11146 3476 11152 3488
rect 11204 3476 11210 3528
rect 11882 3476 11888 3528
rect 11940 3516 11946 3528
rect 11977 3519 12035 3525
rect 11977 3516 11989 3519
rect 11940 3488 11989 3516
rect 11940 3476 11946 3488
rect 11977 3485 11989 3488
rect 12023 3485 12035 3519
rect 11977 3479 12035 3485
rect 11054 3380 11060 3392
rect 10244 3352 11060 3380
rect 9861 3343 9919 3349
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 1104 3290 16100 3312
rect 1104 3238 3481 3290
rect 3533 3238 3545 3290
rect 3597 3238 3609 3290
rect 3661 3238 3673 3290
rect 3725 3238 8480 3290
rect 8532 3238 8544 3290
rect 8596 3238 8608 3290
rect 8660 3238 8672 3290
rect 8724 3238 13478 3290
rect 13530 3238 13542 3290
rect 13594 3238 13606 3290
rect 13658 3238 13670 3290
rect 13722 3238 16100 3290
rect 1104 3216 16100 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3176 1639 3179
rect 5074 3176 5080 3188
rect 1627 3148 5080 3176
rect 1627 3145 1639 3148
rect 1581 3139 1639 3145
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 6181 3179 6239 3185
rect 6181 3145 6193 3179
rect 6227 3176 6239 3179
rect 7098 3176 7104 3188
rect 6227 3148 7104 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 7098 3136 7104 3148
rect 7156 3136 7162 3188
rect 9122 3176 9128 3188
rect 9083 3148 9128 3176
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 9214 3136 9220 3188
rect 9272 3176 9278 3188
rect 9309 3179 9367 3185
rect 9309 3176 9321 3179
rect 9272 3148 9321 3176
rect 9272 3136 9278 3148
rect 9309 3145 9321 3148
rect 9355 3145 9367 3179
rect 11146 3176 11152 3188
rect 11107 3148 11152 3176
rect 9309 3139 9367 3145
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 14274 3136 14280 3188
rect 14332 3176 14338 3188
rect 14553 3179 14611 3185
rect 14553 3176 14565 3179
rect 14332 3148 14565 3176
rect 14332 3136 14338 3148
rect 14553 3145 14565 3148
rect 14599 3145 14611 3179
rect 14918 3176 14924 3188
rect 14879 3148 14924 3176
rect 14553 3139 14611 3145
rect 14918 3136 14924 3148
rect 14976 3136 14982 3188
rect 3234 3068 3240 3120
rect 3292 3108 3298 3120
rect 3881 3111 3939 3117
rect 3292 3080 3832 3108
rect 3292 3068 3298 3080
rect 2774 3000 2780 3052
rect 2832 3040 2838 3052
rect 3145 3043 3203 3049
rect 3145 3040 3157 3043
rect 2832 3012 3157 3040
rect 2832 3000 2838 3012
rect 3145 3009 3157 3012
rect 3191 3040 3203 3043
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 3191 3012 3617 3040
rect 3191 3009 3203 3012
rect 3145 3003 3203 3009
rect 3605 3009 3617 3012
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 474 2932 480 2984
rect 532 2972 538 2984
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 532 2944 1409 2972
rect 532 2932 538 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 1946 2932 1952 2984
rect 2004 2972 2010 2984
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 2004 2944 2237 2972
rect 2004 2932 2010 2944
rect 2225 2941 2237 2944
rect 2271 2941 2283 2975
rect 2225 2935 2283 2941
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2972 2927 2975
rect 2958 2972 2964 2984
rect 2915 2944 2964 2972
rect 2915 2941 2927 2944
rect 2869 2935 2927 2941
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 3053 2975 3111 2981
rect 3053 2941 3065 2975
rect 3099 2941 3111 2975
rect 3234 2972 3240 2984
rect 3195 2944 3240 2972
rect 3053 2935 3111 2941
rect 1670 2864 1676 2916
rect 1728 2904 1734 2916
rect 2685 2907 2743 2913
rect 2685 2904 2697 2907
rect 1728 2876 2697 2904
rect 1728 2864 1734 2876
rect 2685 2873 2697 2876
rect 2731 2873 2743 2907
rect 3068 2904 3096 2935
rect 3234 2932 3240 2944
rect 3292 2932 3298 2984
rect 3326 2932 3332 2984
rect 3384 2972 3390 2984
rect 3421 2975 3479 2981
rect 3421 2972 3433 2975
rect 3384 2944 3433 2972
rect 3384 2932 3390 2944
rect 3421 2941 3433 2944
rect 3467 2941 3479 2975
rect 3421 2935 3479 2941
rect 3510 2932 3516 2984
rect 3568 2972 3574 2984
rect 3697 2975 3755 2981
rect 3568 2944 3613 2972
rect 3568 2932 3574 2944
rect 3697 2941 3709 2975
rect 3743 2941 3755 2975
rect 3804 2972 3832 3080
rect 3881 3077 3893 3111
rect 3927 3108 3939 3111
rect 4154 3108 4160 3120
rect 3927 3080 4160 3108
rect 3927 3077 3939 3080
rect 3881 3071 3939 3077
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 4430 3068 4436 3120
rect 4488 3108 4494 3120
rect 5813 3111 5871 3117
rect 5813 3108 5825 3111
rect 4488 3080 5825 3108
rect 4488 3068 4494 3080
rect 5813 3077 5825 3080
rect 5859 3108 5871 3111
rect 6089 3111 6147 3117
rect 6089 3108 6101 3111
rect 5859 3080 6101 3108
rect 5859 3077 5871 3080
rect 5813 3071 5871 3077
rect 6089 3077 6101 3080
rect 6135 3108 6147 3111
rect 6638 3108 6644 3120
rect 6135 3080 6644 3108
rect 6135 3077 6147 3080
rect 6089 3071 6147 3077
rect 6638 3068 6644 3080
rect 6696 3068 6702 3120
rect 9674 3068 9680 3120
rect 9732 3068 9738 3120
rect 4246 3040 4252 3052
rect 4159 3012 4252 3040
rect 4065 2975 4123 2981
rect 4065 2972 4077 2975
rect 3804 2944 4077 2972
rect 3697 2935 3755 2941
rect 4065 2941 4077 2944
rect 4111 2941 4123 2975
rect 4065 2935 4123 2941
rect 3712 2904 3740 2935
rect 4172 2913 4200 3012
rect 4246 3000 4252 3012
rect 4304 3040 4310 3052
rect 4801 3043 4859 3049
rect 4801 3040 4813 3043
rect 4304 3012 4813 3040
rect 4304 3000 4310 3012
rect 4801 3009 4813 3012
rect 4847 3009 4859 3043
rect 6178 3040 6184 3052
rect 4801 3003 4859 3009
rect 5736 3012 6184 3040
rect 4430 2972 4436 2984
rect 4391 2944 4436 2972
rect 4430 2932 4436 2944
rect 4488 2932 4494 2984
rect 4522 2932 4528 2984
rect 4580 2972 4586 2984
rect 4893 2975 4951 2981
rect 4580 2944 4625 2972
rect 4580 2932 4586 2944
rect 4893 2941 4905 2975
rect 4939 2941 4951 2975
rect 5166 2972 5172 2984
rect 5127 2944 5172 2972
rect 4893 2935 4951 2941
rect 4157 2907 4215 2913
rect 4157 2904 4169 2907
rect 3068 2876 4169 2904
rect 2685 2867 2743 2873
rect 4157 2873 4169 2876
rect 4203 2873 4215 2907
rect 4157 2867 4215 2873
rect 4249 2907 4307 2913
rect 4249 2873 4261 2907
rect 4295 2873 4307 2907
rect 4908 2904 4936 2935
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 5626 2932 5632 2984
rect 5684 2972 5690 2984
rect 5736 2981 5764 3012
rect 6178 3000 6184 3012
rect 6236 3000 6242 3052
rect 6273 3043 6331 3049
rect 6273 3009 6285 3043
rect 6319 3009 6331 3043
rect 6273 3003 6331 3009
rect 5721 2975 5779 2981
rect 5721 2972 5733 2975
rect 5684 2944 5733 2972
rect 5684 2932 5690 2944
rect 5721 2941 5733 2944
rect 5767 2941 5779 2975
rect 5721 2935 5779 2941
rect 5997 2975 6055 2981
rect 5997 2941 6009 2975
rect 6043 2941 6055 2975
rect 6288 2972 6316 3003
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 7377 3043 7435 3049
rect 7377 3040 7389 3043
rect 6972 3012 7389 3040
rect 6972 3000 6978 3012
rect 7377 3009 7389 3012
rect 7423 3040 7435 3043
rect 7650 3040 7656 3052
rect 7423 3012 7656 3040
rect 7423 3009 7435 3012
rect 7377 3003 7435 3009
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 9692 3040 9720 3068
rect 10781 3043 10839 3049
rect 10781 3040 10793 3043
rect 9692 3012 10793 3040
rect 10781 3009 10793 3012
rect 10827 3009 10839 3043
rect 11054 3040 11060 3052
rect 11015 3012 11060 3040
rect 10781 3003 10839 3009
rect 11054 3000 11060 3012
rect 11112 3040 11118 3052
rect 12434 3040 12440 3052
rect 11112 3012 12440 3040
rect 11112 3000 11118 3012
rect 12434 3000 12440 3012
rect 12492 3040 12498 3052
rect 12805 3043 12863 3049
rect 12805 3040 12817 3043
rect 12492 3012 12817 3040
rect 12492 3000 12498 3012
rect 12805 3009 12817 3012
rect 12851 3009 12863 3043
rect 12805 3003 12863 3009
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 15562 3040 15568 3052
rect 13127 3012 15568 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 15562 3000 15568 3012
rect 15620 3000 15626 3052
rect 6546 2972 6552 2984
rect 6288 2944 6552 2972
rect 5997 2935 6055 2941
rect 6012 2904 6040 2935
rect 6546 2932 6552 2944
rect 6604 2932 6610 2984
rect 6822 2972 6828 2984
rect 6783 2944 6828 2972
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 11333 2975 11391 2981
rect 11333 2941 11345 2975
rect 11379 2972 11391 2975
rect 11882 2972 11888 2984
rect 11379 2944 11888 2972
rect 11379 2941 11391 2944
rect 11333 2935 11391 2941
rect 11882 2932 11888 2944
rect 11940 2932 11946 2984
rect 14737 2975 14795 2981
rect 14737 2941 14749 2975
rect 14783 2941 14795 2975
rect 14737 2935 14795 2941
rect 6840 2904 6868 2932
rect 7650 2904 7656 2916
rect 4908 2876 5948 2904
rect 6012 2876 6868 2904
rect 7611 2876 7656 2904
rect 4249 2867 4307 2873
rect 2406 2836 2412 2848
rect 2367 2808 2412 2836
rect 2406 2796 2412 2808
rect 2464 2796 2470 2848
rect 3510 2796 3516 2848
rect 3568 2836 3574 2848
rect 3970 2836 3976 2848
rect 3568 2808 3976 2836
rect 3568 2796 3574 2808
rect 3970 2796 3976 2808
rect 4028 2836 4034 2848
rect 4264 2836 4292 2867
rect 4028 2808 4292 2836
rect 4028 2796 4034 2808
rect 4890 2796 4896 2848
rect 4948 2836 4954 2848
rect 4985 2839 5043 2845
rect 4985 2836 4997 2839
rect 4948 2808 4997 2836
rect 4948 2796 4954 2808
rect 4985 2805 4997 2808
rect 5031 2805 5043 2839
rect 5920 2836 5948 2876
rect 7650 2864 7656 2876
rect 7708 2864 7714 2916
rect 8662 2864 8668 2916
rect 8720 2864 8726 2916
rect 9766 2864 9772 2916
rect 9824 2864 9830 2916
rect 11517 2907 11575 2913
rect 11517 2873 11529 2907
rect 11563 2904 11575 2907
rect 11698 2904 11704 2916
rect 11563 2876 11704 2904
rect 11563 2873 11575 2876
rect 11517 2867 11575 2873
rect 11698 2864 11704 2876
rect 11756 2864 11762 2916
rect 13814 2864 13820 2916
rect 13872 2864 13878 2916
rect 7009 2839 7067 2845
rect 7009 2836 7021 2839
rect 5920 2808 7021 2836
rect 4985 2799 5043 2805
rect 7009 2805 7021 2808
rect 7055 2836 7067 2839
rect 7374 2836 7380 2848
rect 7055 2808 7380 2836
rect 7055 2805 7067 2808
rect 7009 2799 7067 2805
rect 7374 2796 7380 2808
rect 7432 2796 7438 2848
rect 13722 2796 13728 2848
rect 13780 2836 13786 2848
rect 14752 2836 14780 2935
rect 13780 2808 14780 2836
rect 13780 2796 13786 2808
rect 1104 2746 16100 2768
rect 1104 2694 5980 2746
rect 6032 2694 6044 2746
rect 6096 2694 6108 2746
rect 6160 2694 6172 2746
rect 6224 2694 10979 2746
rect 11031 2694 11043 2746
rect 11095 2694 11107 2746
rect 11159 2694 11171 2746
rect 11223 2694 16100 2746
rect 1104 2672 16100 2694
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3145 2635 3203 2641
rect 3145 2632 3157 2635
rect 3016 2604 3157 2632
rect 3016 2592 3022 2604
rect 3145 2601 3157 2604
rect 3191 2632 3203 2635
rect 3970 2632 3976 2644
rect 3191 2604 3976 2632
rect 3191 2601 3203 2604
rect 3145 2595 3203 2601
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 5626 2632 5632 2644
rect 5587 2604 5632 2632
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 5905 2635 5963 2641
rect 5905 2601 5917 2635
rect 5951 2632 5963 2635
rect 6733 2635 6791 2641
rect 5951 2604 6224 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 1670 2564 1676 2576
rect 1631 2536 1676 2564
rect 1670 2524 1676 2536
rect 1728 2524 1734 2576
rect 2406 2524 2412 2576
rect 2464 2524 2470 2576
rect 4154 2564 4160 2576
rect 4115 2536 4160 2564
rect 4154 2524 4160 2536
rect 4212 2524 4218 2576
rect 4890 2524 4896 2576
rect 4948 2524 4954 2576
rect 6196 2573 6224 2604
rect 6733 2601 6745 2635
rect 6779 2632 6791 2635
rect 6822 2632 6828 2644
rect 6779 2604 6828 2632
rect 6779 2601 6791 2604
rect 6733 2595 6791 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 7469 2635 7527 2641
rect 7469 2601 7481 2635
rect 7515 2632 7527 2635
rect 7650 2632 7656 2644
rect 7515 2604 7656 2632
rect 7515 2601 7527 2604
rect 7469 2595 7527 2601
rect 7650 2592 7656 2604
rect 7708 2592 7714 2644
rect 8573 2635 8631 2641
rect 8573 2601 8585 2635
rect 8619 2632 8631 2635
rect 8662 2632 8668 2644
rect 8619 2604 8668 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 11241 2635 11299 2641
rect 11241 2601 11253 2635
rect 11287 2632 11299 2635
rect 11514 2632 11520 2644
rect 11287 2604 11520 2632
rect 11287 2601 11299 2604
rect 11241 2595 11299 2601
rect 11514 2592 11520 2604
rect 11572 2592 11578 2644
rect 12158 2632 12164 2644
rect 12119 2604 12164 2632
rect 12158 2592 12164 2604
rect 12216 2592 12222 2644
rect 13814 2592 13820 2644
rect 13872 2632 13878 2644
rect 13909 2635 13967 2641
rect 13909 2632 13921 2635
rect 13872 2604 13921 2632
rect 13872 2592 13878 2604
rect 13909 2601 13921 2604
rect 13955 2601 13967 2635
rect 15562 2632 15568 2644
rect 15523 2604 15568 2632
rect 13909 2595 13967 2601
rect 15562 2592 15568 2604
rect 15620 2592 15626 2644
rect 6181 2567 6239 2573
rect 6181 2533 6193 2567
rect 6227 2533 6239 2567
rect 6181 2527 6239 2533
rect 7006 2524 7012 2576
rect 7064 2564 7070 2576
rect 7101 2567 7159 2573
rect 7101 2564 7113 2567
rect 7064 2536 7113 2564
rect 7064 2524 7070 2536
rect 7101 2533 7113 2536
rect 7147 2533 7159 2567
rect 7101 2527 7159 2533
rect 7190 2524 7196 2576
rect 7248 2564 7254 2576
rect 7285 2567 7343 2573
rect 7285 2564 7297 2567
rect 7248 2536 7297 2564
rect 7248 2524 7254 2536
rect 7285 2533 7297 2536
rect 7331 2533 7343 2567
rect 7285 2527 7343 2533
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2456 1458 2508
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2465 5779 2499
rect 5721 2459 5779 2465
rect 1412 2428 1440 2456
rect 3881 2431 3939 2437
rect 3881 2428 3893 2431
rect 1412 2400 3893 2428
rect 3881 2397 3893 2400
rect 3927 2428 3939 2431
rect 5736 2428 5764 2459
rect 6454 2456 6460 2508
rect 6512 2496 6518 2508
rect 6825 2499 6883 2505
rect 6825 2496 6837 2499
rect 6512 2468 6837 2496
rect 6512 2456 6518 2468
rect 6825 2465 6837 2468
rect 6871 2465 6883 2499
rect 6825 2459 6883 2465
rect 8389 2499 8447 2505
rect 8389 2465 8401 2499
rect 8435 2496 8447 2499
rect 10042 2496 10048 2508
rect 8435 2468 10048 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 10042 2456 10048 2468
rect 10100 2496 10106 2508
rect 11057 2499 11115 2505
rect 11057 2496 11069 2499
rect 10100 2468 11069 2496
rect 10100 2456 10106 2468
rect 11057 2465 11069 2468
rect 11103 2465 11115 2499
rect 11974 2496 11980 2508
rect 11935 2468 11980 2496
rect 11057 2459 11115 2465
rect 11974 2456 11980 2468
rect 12032 2456 12038 2508
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 13722 2496 13728 2508
rect 12492 2468 13728 2496
rect 12492 2456 12498 2468
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 15746 2496 15752 2508
rect 15707 2468 15752 2496
rect 15746 2456 15752 2468
rect 15804 2456 15810 2508
rect 3927 2400 5764 2428
rect 3927 2397 3939 2400
rect 3881 2391 3939 2397
rect 5994 2360 6000 2372
rect 5955 2332 6000 2360
rect 5994 2320 6000 2332
rect 6052 2320 6058 2372
rect 1104 2202 16100 2224
rect 1104 2150 3481 2202
rect 3533 2150 3545 2202
rect 3597 2150 3609 2202
rect 3661 2150 3673 2202
rect 3725 2150 8480 2202
rect 8532 2150 8544 2202
rect 8596 2150 8608 2202
rect 8660 2150 8672 2202
rect 8724 2150 13478 2202
rect 13530 2150 13542 2202
rect 13594 2150 13606 2202
rect 13658 2150 13670 2202
rect 13722 2150 16100 2202
rect 1104 2128 16100 2150
<< via1 >>
rect 5980 16838 6032 16890
rect 6044 16838 6096 16890
rect 6108 16838 6160 16890
rect 6172 16838 6224 16890
rect 10979 16838 11031 16890
rect 11043 16838 11095 16890
rect 11107 16838 11159 16890
rect 11171 16838 11223 16890
rect 2320 16736 2372 16788
rect 4528 16736 4580 16788
rect 11336 16736 11388 16788
rect 6736 16668 6788 16720
rect 16580 16668 16632 16720
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 5080 16600 5132 16652
rect 11244 16643 11296 16652
rect 11244 16609 11253 16643
rect 11253 16609 11287 16643
rect 11287 16609 11296 16643
rect 11244 16600 11296 16609
rect 3481 16294 3533 16346
rect 3545 16294 3597 16346
rect 3609 16294 3661 16346
rect 3673 16294 3725 16346
rect 8480 16294 8532 16346
rect 8544 16294 8596 16346
rect 8608 16294 8660 16346
rect 8672 16294 8724 16346
rect 13478 16294 13530 16346
rect 13542 16294 13594 16346
rect 13606 16294 13658 16346
rect 13670 16294 13722 16346
rect 3792 16192 3844 16244
rect 11244 16192 11296 16244
rect 3424 16124 3476 16176
rect 4436 16124 4488 16176
rect 3148 16056 3200 16108
rect 4712 16099 4764 16108
rect 4712 16065 4721 16099
rect 4721 16065 4755 16099
rect 4755 16065 4764 16099
rect 4712 16056 4764 16065
rect 3516 15988 3568 16040
rect 6552 16056 6604 16108
rect 5080 15988 5132 16040
rect 5356 16031 5408 16040
rect 5356 15997 5365 16031
rect 5365 15997 5399 16031
rect 5399 15997 5408 16031
rect 5356 15988 5408 15997
rect 6644 16031 6696 16040
rect 6644 15997 6653 16031
rect 6653 15997 6687 16031
rect 6687 15997 6696 16031
rect 6644 15988 6696 15997
rect 7012 15988 7064 16040
rect 2412 15963 2464 15972
rect 2412 15929 2421 15963
rect 2421 15929 2455 15963
rect 2455 15929 2464 15963
rect 2412 15920 2464 15929
rect 4252 15920 4304 15972
rect 9864 15988 9916 16040
rect 13268 16031 13320 16040
rect 9220 15963 9272 15972
rect 4620 15852 4672 15904
rect 5080 15852 5132 15904
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 5816 15852 5868 15904
rect 6552 15895 6604 15904
rect 6552 15861 6561 15895
rect 6561 15861 6595 15895
rect 6595 15861 6604 15895
rect 6552 15852 6604 15861
rect 9220 15929 9229 15963
rect 9229 15929 9263 15963
rect 9263 15929 9272 15963
rect 9220 15920 9272 15929
rect 13268 15997 13277 16031
rect 13277 15997 13311 16031
rect 13311 15997 13320 16031
rect 13268 15988 13320 15997
rect 13544 15852 13596 15904
rect 13728 15895 13780 15904
rect 13728 15861 13737 15895
rect 13737 15861 13771 15895
rect 13771 15861 13780 15895
rect 13728 15852 13780 15861
rect 13820 15895 13872 15904
rect 13820 15861 13829 15895
rect 13829 15861 13863 15895
rect 13863 15861 13872 15895
rect 13820 15852 13872 15861
rect 5980 15750 6032 15802
rect 6044 15750 6096 15802
rect 6108 15750 6160 15802
rect 6172 15750 6224 15802
rect 10979 15750 11031 15802
rect 11043 15750 11095 15802
rect 11107 15750 11159 15802
rect 11171 15750 11223 15802
rect 2412 15648 2464 15700
rect 3516 15691 3568 15700
rect 3516 15657 3525 15691
rect 3525 15657 3559 15691
rect 3559 15657 3568 15691
rect 3516 15648 3568 15657
rect 4160 15648 4212 15700
rect 4712 15691 4764 15700
rect 4712 15657 4721 15691
rect 4721 15657 4755 15691
rect 4755 15657 4764 15691
rect 4712 15648 4764 15657
rect 5172 15648 5224 15700
rect 7012 15691 7064 15700
rect 7012 15657 7021 15691
rect 7021 15657 7055 15691
rect 7055 15657 7064 15691
rect 7012 15648 7064 15657
rect 9220 15648 9272 15700
rect 5080 15623 5132 15632
rect 5080 15589 5089 15623
rect 5089 15589 5123 15623
rect 5123 15589 5132 15623
rect 5080 15580 5132 15589
rect 5816 15580 5868 15632
rect 13728 15648 13780 15700
rect 2872 15487 2924 15496
rect 2872 15453 2881 15487
rect 2881 15453 2915 15487
rect 2915 15453 2924 15487
rect 2872 15444 2924 15453
rect 3424 15512 3476 15564
rect 3792 15512 3844 15564
rect 4252 15555 4304 15564
rect 4252 15521 4259 15555
rect 4259 15521 4304 15555
rect 4252 15512 4304 15521
rect 4344 15555 4396 15564
rect 4344 15521 4353 15555
rect 4353 15521 4387 15555
rect 4387 15521 4396 15555
rect 4344 15512 4396 15521
rect 4712 15512 4764 15564
rect 6460 15512 6512 15564
rect 7012 15555 7064 15564
rect 7012 15521 7021 15555
rect 7021 15521 7055 15555
rect 7055 15521 7064 15555
rect 7012 15512 7064 15521
rect 9588 15555 9640 15564
rect 9588 15521 9597 15555
rect 9597 15521 9631 15555
rect 9631 15521 9640 15555
rect 9588 15512 9640 15521
rect 12440 15512 12492 15564
rect 13268 15580 13320 15632
rect 13544 15555 13596 15564
rect 4252 15376 4304 15428
rect 3240 15308 3292 15360
rect 13544 15521 13553 15555
rect 13553 15521 13587 15555
rect 13587 15521 13596 15555
rect 13544 15512 13596 15521
rect 13820 15555 13872 15564
rect 13820 15521 13829 15555
rect 13829 15521 13863 15555
rect 13863 15521 13872 15555
rect 13820 15512 13872 15521
rect 14188 15487 14240 15496
rect 14188 15453 14197 15487
rect 14197 15453 14231 15487
rect 14231 15453 14240 15487
rect 14188 15444 14240 15453
rect 4712 15308 4764 15360
rect 5264 15308 5316 15360
rect 5816 15308 5868 15360
rect 6644 15308 6696 15360
rect 15016 15419 15068 15428
rect 15016 15385 15025 15419
rect 15025 15385 15059 15419
rect 15059 15385 15068 15419
rect 15016 15376 15068 15385
rect 3481 15206 3533 15258
rect 3545 15206 3597 15258
rect 3609 15206 3661 15258
rect 3673 15206 3725 15258
rect 8480 15206 8532 15258
rect 8544 15206 8596 15258
rect 8608 15206 8660 15258
rect 8672 15206 8724 15258
rect 13478 15206 13530 15258
rect 13542 15206 13594 15258
rect 13606 15206 13658 15258
rect 13670 15206 13722 15258
rect 4344 15104 4396 15156
rect 4988 15104 5040 15156
rect 9588 15104 9640 15156
rect 4620 14900 4672 14952
rect 7656 14900 7708 14952
rect 8208 14900 8260 14952
rect 9036 14943 9088 14952
rect 9036 14909 9045 14943
rect 9045 14909 9079 14943
rect 9079 14909 9088 14943
rect 9036 14900 9088 14909
rect 9128 14943 9180 14952
rect 9128 14909 9137 14943
rect 9137 14909 9171 14943
rect 9171 14909 9180 14943
rect 9128 14900 9180 14909
rect 4160 14832 4212 14884
rect 6460 14875 6512 14884
rect 6460 14841 6469 14875
rect 6469 14841 6503 14875
rect 6503 14841 6512 14875
rect 6460 14832 6512 14841
rect 8852 14832 8904 14884
rect 11612 14832 11664 14884
rect 5980 14662 6032 14714
rect 6044 14662 6096 14714
rect 6108 14662 6160 14714
rect 6172 14662 6224 14714
rect 10979 14662 11031 14714
rect 11043 14662 11095 14714
rect 11107 14662 11159 14714
rect 11171 14662 11223 14714
rect 1952 14467 2004 14476
rect 1952 14433 1961 14467
rect 1961 14433 1995 14467
rect 1995 14433 2004 14467
rect 3792 14492 3844 14544
rect 4436 14492 4488 14544
rect 5356 14560 5408 14612
rect 9128 14560 9180 14612
rect 11612 14603 11664 14612
rect 11612 14569 11621 14603
rect 11621 14569 11655 14603
rect 11655 14569 11664 14603
rect 11612 14560 11664 14569
rect 13820 14560 13872 14612
rect 1952 14424 2004 14433
rect 3976 14424 4028 14476
rect 4068 14288 4120 14340
rect 2228 14220 2280 14272
rect 3332 14263 3384 14272
rect 3332 14229 3341 14263
rect 3341 14229 3375 14263
rect 3375 14229 3384 14263
rect 3332 14220 3384 14229
rect 3792 14220 3844 14272
rect 3884 14263 3936 14272
rect 3884 14229 3893 14263
rect 3893 14229 3927 14263
rect 3927 14229 3936 14263
rect 4344 14356 4396 14408
rect 4252 14288 4304 14340
rect 4896 14356 4948 14408
rect 14188 14492 14240 14544
rect 5724 14424 5776 14476
rect 8208 14467 8260 14476
rect 5356 14356 5408 14408
rect 8208 14433 8217 14467
rect 8217 14433 8251 14467
rect 8251 14433 8260 14467
rect 8208 14424 8260 14433
rect 7564 14399 7616 14408
rect 7564 14365 7573 14399
rect 7573 14365 7607 14399
rect 7607 14365 7616 14399
rect 7564 14356 7616 14365
rect 11336 14424 11388 14476
rect 12164 14424 12216 14476
rect 12992 14467 13044 14476
rect 12992 14433 13001 14467
rect 13001 14433 13035 14467
rect 13035 14433 13044 14467
rect 12992 14424 13044 14433
rect 13360 14356 13412 14408
rect 5540 14288 5592 14340
rect 11796 14288 11848 14340
rect 13912 14288 13964 14340
rect 3884 14220 3936 14229
rect 5632 14220 5684 14272
rect 14832 14220 14884 14272
rect 3481 14118 3533 14170
rect 3545 14118 3597 14170
rect 3609 14118 3661 14170
rect 3673 14118 3725 14170
rect 8480 14118 8532 14170
rect 8544 14118 8596 14170
rect 8608 14118 8660 14170
rect 8672 14118 8724 14170
rect 13478 14118 13530 14170
rect 13542 14118 13594 14170
rect 13606 14118 13658 14170
rect 13670 14118 13722 14170
rect 3884 13948 3936 14000
rect 3332 13880 3384 13932
rect 4068 13948 4120 14000
rect 4988 13991 5040 14000
rect 4988 13957 4997 13991
rect 4997 13957 5031 13991
rect 5031 13957 5040 13991
rect 4988 13948 5040 13957
rect 3240 13855 3292 13864
rect 3240 13821 3249 13855
rect 3249 13821 3283 13855
rect 3283 13821 3292 13855
rect 4160 13880 4212 13932
rect 7012 14016 7064 14068
rect 9036 14016 9088 14068
rect 9404 14016 9456 14068
rect 11796 14059 11848 14068
rect 9772 13991 9824 14000
rect 9772 13957 9781 13991
rect 9781 13957 9815 13991
rect 9815 13957 9824 13991
rect 9772 13948 9824 13957
rect 11796 14025 11805 14059
rect 11805 14025 11839 14059
rect 11839 14025 11848 14059
rect 11796 14016 11848 14025
rect 13912 14059 13964 14068
rect 13912 14025 13921 14059
rect 13921 14025 13955 14059
rect 13955 14025 13964 14059
rect 13912 14016 13964 14025
rect 12072 13948 12124 14000
rect 12992 13948 13044 14000
rect 13820 13948 13872 14000
rect 14832 13991 14884 14000
rect 14832 13957 14841 13991
rect 14841 13957 14875 13991
rect 14875 13957 14884 13991
rect 14832 13948 14884 13957
rect 3240 13812 3292 13821
rect 2228 13744 2280 13796
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 2872 13676 2924 13728
rect 3792 13855 3844 13864
rect 3792 13821 3837 13855
rect 3837 13821 3844 13855
rect 3792 13812 3844 13821
rect 4068 13812 4120 13864
rect 4620 13855 4672 13864
rect 4620 13821 4629 13855
rect 4629 13821 4663 13855
rect 4663 13821 4672 13855
rect 4620 13812 4672 13821
rect 4712 13812 4764 13864
rect 4896 13855 4948 13864
rect 4896 13821 4905 13855
rect 4905 13821 4939 13855
rect 4939 13821 4948 13855
rect 4896 13812 4948 13821
rect 5540 13880 5592 13932
rect 5356 13855 5408 13864
rect 5356 13821 5365 13855
rect 5365 13821 5399 13855
rect 5399 13821 5408 13855
rect 5816 13880 5868 13932
rect 9220 13880 9272 13932
rect 9312 13880 9364 13932
rect 5356 13812 5408 13821
rect 6552 13812 6604 13864
rect 7012 13812 7064 13864
rect 7196 13855 7248 13864
rect 7196 13821 7205 13855
rect 7205 13821 7239 13855
rect 7239 13821 7248 13855
rect 7196 13812 7248 13821
rect 9496 13855 9548 13864
rect 9496 13821 9505 13855
rect 9505 13821 9539 13855
rect 9539 13821 9548 13855
rect 9496 13812 9548 13821
rect 9956 13855 10008 13864
rect 9956 13821 9965 13855
rect 9965 13821 9999 13855
rect 9999 13821 10008 13855
rect 9956 13812 10008 13821
rect 13084 13812 13136 13864
rect 13360 13812 13412 13864
rect 14648 13855 14700 13864
rect 10140 13744 10192 13796
rect 14648 13821 14657 13855
rect 14657 13821 14691 13855
rect 14691 13821 14700 13855
rect 14648 13812 14700 13821
rect 15016 13812 15068 13864
rect 3976 13676 4028 13728
rect 4988 13676 5040 13728
rect 11704 13719 11756 13728
rect 11704 13685 11713 13719
rect 11713 13685 11747 13719
rect 11747 13685 11756 13719
rect 11704 13676 11756 13685
rect 14648 13676 14700 13728
rect 5980 13574 6032 13626
rect 6044 13574 6096 13626
rect 6108 13574 6160 13626
rect 6172 13574 6224 13626
rect 10979 13574 11031 13626
rect 11043 13574 11095 13626
rect 11107 13574 11159 13626
rect 11171 13574 11223 13626
rect 4896 13472 4948 13524
rect 5632 13515 5684 13524
rect 5632 13481 5641 13515
rect 5641 13481 5675 13515
rect 5675 13481 5684 13515
rect 5632 13472 5684 13481
rect 5816 13472 5868 13524
rect 4712 13336 4764 13388
rect 5356 13379 5408 13388
rect 1492 13268 1544 13320
rect 4436 13268 4488 13320
rect 5356 13345 5365 13379
rect 5365 13345 5399 13379
rect 5399 13345 5408 13379
rect 5356 13336 5408 13345
rect 5540 13336 5592 13388
rect 6276 13379 6328 13388
rect 6276 13345 6285 13379
rect 6285 13345 6319 13379
rect 6319 13345 6328 13379
rect 7748 13472 7800 13524
rect 6276 13336 6328 13345
rect 5724 13268 5776 13320
rect 6552 13268 6604 13320
rect 6276 13200 6328 13252
rect 7656 13311 7708 13320
rect 7656 13277 7665 13311
rect 7665 13277 7699 13311
rect 7699 13277 7708 13311
rect 7656 13268 7708 13277
rect 9772 13472 9824 13524
rect 8300 13336 8352 13388
rect 11704 13472 11756 13524
rect 13360 13515 13412 13524
rect 13360 13481 13369 13515
rect 13369 13481 13403 13515
rect 13403 13481 13412 13515
rect 13360 13472 13412 13481
rect 12256 13404 12308 13456
rect 14648 13404 14700 13456
rect 8852 13379 8904 13388
rect 8852 13345 8861 13379
rect 8861 13345 8895 13379
rect 8895 13345 8904 13379
rect 8852 13336 8904 13345
rect 9036 13336 9088 13388
rect 7932 13311 7984 13320
rect 7932 13277 7941 13311
rect 7941 13277 7975 13311
rect 7975 13277 7984 13311
rect 9312 13311 9364 13320
rect 7932 13268 7984 13277
rect 9312 13277 9321 13311
rect 9321 13277 9355 13311
rect 9355 13277 9364 13311
rect 9312 13268 9364 13277
rect 10048 13336 10100 13388
rect 11336 13336 11388 13388
rect 12348 13379 12400 13388
rect 12348 13345 12357 13379
rect 12357 13345 12391 13379
rect 12391 13345 12400 13379
rect 12348 13336 12400 13345
rect 12716 13336 12768 13388
rect 12992 13379 13044 13388
rect 12992 13345 13001 13379
rect 13001 13345 13035 13379
rect 13035 13345 13044 13379
rect 12992 13336 13044 13345
rect 13084 13336 13136 13388
rect 12440 13268 12492 13320
rect 7196 13175 7248 13184
rect 7196 13141 7205 13175
rect 7205 13141 7239 13175
rect 7239 13141 7248 13175
rect 7196 13132 7248 13141
rect 12808 13200 12860 13252
rect 14924 13200 14976 13252
rect 12164 13132 12216 13184
rect 3481 13030 3533 13082
rect 3545 13030 3597 13082
rect 3609 13030 3661 13082
rect 3673 13030 3725 13082
rect 8480 13030 8532 13082
rect 8544 13030 8596 13082
rect 8608 13030 8660 13082
rect 8672 13030 8724 13082
rect 13478 13030 13530 13082
rect 13542 13030 13594 13082
rect 13606 13030 13658 13082
rect 13670 13030 13722 13082
rect 7656 12928 7708 12980
rect 8024 12928 8076 12980
rect 9312 12928 9364 12980
rect 9772 12928 9824 12980
rect 12808 12928 12860 12980
rect 1952 12724 2004 12776
rect 3516 12724 3568 12776
rect 5448 12724 5500 12776
rect 7656 12792 7708 12844
rect 7932 12860 7984 12912
rect 8484 12860 8536 12912
rect 6552 12767 6604 12776
rect 3884 12699 3936 12708
rect 3884 12665 3893 12699
rect 3893 12665 3927 12699
rect 3927 12665 3936 12699
rect 3884 12656 3936 12665
rect 5172 12656 5224 12708
rect 6552 12733 6561 12767
rect 6561 12733 6595 12767
rect 6595 12733 6604 12767
rect 6552 12724 6604 12733
rect 7104 12767 7156 12776
rect 6276 12656 6328 12708
rect 2228 12588 2280 12640
rect 4160 12588 4212 12640
rect 5724 12631 5776 12640
rect 5724 12597 5733 12631
rect 5733 12597 5767 12631
rect 5767 12597 5776 12631
rect 5724 12588 5776 12597
rect 7104 12733 7113 12767
rect 7113 12733 7147 12767
rect 7147 12733 7156 12767
rect 7104 12724 7156 12733
rect 7840 12724 7892 12776
rect 9404 12792 9456 12844
rect 8484 12724 8536 12776
rect 9772 12724 9824 12776
rect 13360 12767 13412 12776
rect 13360 12733 13369 12767
rect 13369 12733 13403 12767
rect 13403 12733 13412 12767
rect 13360 12724 13412 12733
rect 14924 12724 14976 12776
rect 7196 12699 7248 12708
rect 7196 12665 7205 12699
rect 7205 12665 7239 12699
rect 7239 12665 7248 12699
rect 7196 12656 7248 12665
rect 7288 12656 7340 12708
rect 7932 12699 7984 12708
rect 7932 12665 7941 12699
rect 7941 12665 7975 12699
rect 7975 12665 7984 12699
rect 7932 12656 7984 12665
rect 8300 12699 8352 12708
rect 8300 12665 8309 12699
rect 8309 12665 8343 12699
rect 8343 12665 8352 12699
rect 8300 12656 8352 12665
rect 15016 12656 15068 12708
rect 7748 12588 7800 12640
rect 13728 12631 13780 12640
rect 13728 12597 13737 12631
rect 13737 12597 13771 12631
rect 13771 12597 13780 12631
rect 13728 12588 13780 12597
rect 5980 12486 6032 12538
rect 6044 12486 6096 12538
rect 6108 12486 6160 12538
rect 6172 12486 6224 12538
rect 10979 12486 11031 12538
rect 11043 12486 11095 12538
rect 11107 12486 11159 12538
rect 11171 12486 11223 12538
rect 3884 12384 3936 12436
rect 4988 12384 5040 12436
rect 5356 12384 5408 12436
rect 2228 12316 2280 12368
rect 2872 12316 2924 12368
rect 4160 12359 4212 12368
rect 4160 12325 4169 12359
rect 4169 12325 4203 12359
rect 4203 12325 4212 12359
rect 4160 12316 4212 12325
rect 4252 12359 4304 12368
rect 4252 12325 4261 12359
rect 4261 12325 4295 12359
rect 4295 12325 4304 12359
rect 6092 12359 6144 12368
rect 4252 12316 4304 12325
rect 6092 12325 6101 12359
rect 6101 12325 6135 12359
rect 6135 12325 6144 12359
rect 6092 12316 6144 12325
rect 3240 12291 3292 12300
rect 3240 12257 3249 12291
rect 3249 12257 3283 12291
rect 3283 12257 3292 12291
rect 3516 12291 3568 12300
rect 3240 12248 3292 12257
rect 3516 12257 3525 12291
rect 3525 12257 3559 12291
rect 3559 12257 3568 12291
rect 3516 12248 3568 12257
rect 3884 12248 3936 12300
rect 4620 12291 4672 12300
rect 1676 12180 1728 12232
rect 2872 12180 2924 12232
rect 4620 12257 4629 12291
rect 4629 12257 4663 12291
rect 4663 12257 4672 12291
rect 4988 12291 5040 12300
rect 4620 12248 4672 12257
rect 4988 12257 4997 12291
rect 4997 12257 5031 12291
rect 5031 12257 5040 12291
rect 4988 12248 5040 12257
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5172 12248 5224 12257
rect 5724 12248 5776 12300
rect 4344 12044 4396 12096
rect 4436 12044 4488 12096
rect 5080 12180 5132 12232
rect 5816 12180 5868 12232
rect 5448 12112 5500 12164
rect 4712 12087 4764 12096
rect 4712 12053 4721 12087
rect 4721 12053 4755 12087
rect 4755 12053 4764 12087
rect 6000 12291 6052 12300
rect 6000 12257 6009 12291
rect 6009 12257 6043 12291
rect 6043 12257 6052 12291
rect 6920 12384 6972 12436
rect 8392 12384 8444 12436
rect 9772 12427 9824 12436
rect 9772 12393 9781 12427
rect 9781 12393 9815 12427
rect 9815 12393 9824 12427
rect 9772 12384 9824 12393
rect 11336 12384 11388 12436
rect 6000 12248 6052 12257
rect 6460 12291 6512 12300
rect 6460 12257 6469 12291
rect 6469 12257 6503 12291
rect 6503 12257 6512 12291
rect 6460 12248 6512 12257
rect 6552 12291 6604 12300
rect 6552 12257 6561 12291
rect 6561 12257 6595 12291
rect 6595 12257 6604 12291
rect 6552 12248 6604 12257
rect 7012 12248 7064 12300
rect 7656 12316 7708 12368
rect 8116 12316 8168 12368
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 8300 12316 8352 12368
rect 9864 12359 9916 12368
rect 8484 12291 8536 12300
rect 8484 12257 8493 12291
rect 8493 12257 8527 12291
rect 8527 12257 8536 12291
rect 8484 12248 8536 12257
rect 6920 12223 6972 12232
rect 6920 12189 6929 12223
rect 6929 12189 6963 12223
rect 6963 12189 6972 12223
rect 6920 12180 6972 12189
rect 6276 12112 6328 12164
rect 7932 12155 7984 12164
rect 7932 12121 7941 12155
rect 7941 12121 7975 12155
rect 7975 12121 7984 12155
rect 9036 12248 9088 12300
rect 9312 12291 9364 12300
rect 9312 12257 9322 12291
rect 9322 12257 9356 12291
rect 9356 12257 9364 12291
rect 9588 12291 9640 12300
rect 9312 12248 9364 12257
rect 9588 12257 9597 12291
rect 9597 12257 9631 12291
rect 9631 12257 9640 12291
rect 9588 12248 9640 12257
rect 9864 12325 9873 12359
rect 9873 12325 9907 12359
rect 9907 12325 9916 12359
rect 9864 12316 9916 12325
rect 12440 12316 12492 12368
rect 13176 12359 13228 12368
rect 13176 12325 13185 12359
rect 13185 12325 13219 12359
rect 13219 12325 13228 12359
rect 13176 12316 13228 12325
rect 9220 12180 9272 12232
rect 9772 12180 9824 12232
rect 11060 12248 11112 12300
rect 12164 12248 12216 12300
rect 13360 12248 13412 12300
rect 12992 12180 13044 12232
rect 13728 12359 13780 12368
rect 13728 12325 13737 12359
rect 13737 12325 13771 12359
rect 13771 12325 13780 12359
rect 13728 12316 13780 12325
rect 14924 12291 14976 12300
rect 14924 12257 14943 12291
rect 14943 12257 14976 12291
rect 14924 12248 14976 12257
rect 15016 12291 15068 12300
rect 15016 12257 15025 12291
rect 15025 12257 15059 12291
rect 15059 12257 15068 12291
rect 15016 12248 15068 12257
rect 7932 12112 7984 12121
rect 4712 12044 4764 12053
rect 8300 12044 8352 12096
rect 9312 12112 9364 12164
rect 8944 12044 8996 12096
rect 9496 12155 9548 12164
rect 9496 12121 9505 12155
rect 9505 12121 9539 12155
rect 9539 12121 9548 12155
rect 9496 12112 9548 12121
rect 9864 12112 9916 12164
rect 10232 12155 10284 12164
rect 10232 12121 10241 12155
rect 10241 12121 10275 12155
rect 10275 12121 10284 12155
rect 12348 12155 12400 12164
rect 10232 12112 10284 12121
rect 12348 12121 12357 12155
rect 12357 12121 12391 12155
rect 12391 12121 12400 12155
rect 12348 12112 12400 12121
rect 12440 12155 12492 12164
rect 12440 12121 12449 12155
rect 12449 12121 12483 12155
rect 12483 12121 12492 12155
rect 12440 12112 12492 12121
rect 12256 12044 12308 12096
rect 12716 12044 12768 12096
rect 15016 12087 15068 12096
rect 15016 12053 15025 12087
rect 15025 12053 15059 12087
rect 15059 12053 15068 12087
rect 15016 12044 15068 12053
rect 3481 11942 3533 11994
rect 3545 11942 3597 11994
rect 3609 11942 3661 11994
rect 3673 11942 3725 11994
rect 8480 11942 8532 11994
rect 8544 11942 8596 11994
rect 8608 11942 8660 11994
rect 8672 11942 8724 11994
rect 13478 11942 13530 11994
rect 13542 11942 13594 11994
rect 13606 11942 13658 11994
rect 13670 11942 13722 11994
rect 6460 11840 6512 11892
rect 8300 11840 8352 11892
rect 2780 11772 2832 11824
rect 4068 11772 4120 11824
rect 4436 11772 4488 11824
rect 8944 11772 8996 11824
rect 9588 11840 9640 11892
rect 9864 11840 9916 11892
rect 11060 11883 11112 11892
rect 11060 11849 11069 11883
rect 11069 11849 11103 11883
rect 11103 11849 11112 11883
rect 11060 11840 11112 11849
rect 4344 11636 4396 11688
rect 5356 11636 5408 11688
rect 6000 11636 6052 11688
rect 8760 11679 8812 11688
rect 8760 11645 8769 11679
rect 8769 11645 8803 11679
rect 8803 11645 8812 11679
rect 8760 11636 8812 11645
rect 8944 11679 8996 11688
rect 8944 11645 8953 11679
rect 8953 11645 8987 11679
rect 8987 11645 8996 11679
rect 8944 11636 8996 11645
rect 6736 11611 6788 11620
rect 6736 11577 6745 11611
rect 6745 11577 6779 11611
rect 6779 11577 6788 11611
rect 6736 11568 6788 11577
rect 9128 11636 9180 11688
rect 10416 11772 10468 11824
rect 9588 11636 9640 11688
rect 9680 11636 9732 11688
rect 10600 11704 10652 11756
rect 12256 11704 12308 11756
rect 10508 11679 10560 11688
rect 10508 11645 10517 11679
rect 10517 11645 10551 11679
rect 10551 11645 10560 11679
rect 10508 11636 10560 11645
rect 10876 11636 10928 11688
rect 12440 11636 12492 11688
rect 5448 11500 5500 11552
rect 6276 11500 6328 11552
rect 8116 11500 8168 11552
rect 8300 11500 8352 11552
rect 9312 11500 9364 11552
rect 9588 11500 9640 11552
rect 11888 11568 11940 11620
rect 12348 11568 12400 11620
rect 13176 11636 13228 11688
rect 5980 11398 6032 11450
rect 6044 11398 6096 11450
rect 6108 11398 6160 11450
rect 6172 11398 6224 11450
rect 10979 11398 11031 11450
rect 11043 11398 11095 11450
rect 11107 11398 11159 11450
rect 11171 11398 11223 11450
rect 5356 11339 5408 11348
rect 5356 11305 5365 11339
rect 5365 11305 5399 11339
rect 5399 11305 5408 11339
rect 5356 11296 5408 11305
rect 2136 11228 2188 11280
rect 6920 11228 6972 11280
rect 4436 11203 4488 11212
rect 4436 11169 4445 11203
rect 4445 11169 4479 11203
rect 4479 11169 4488 11203
rect 4436 11160 4488 11169
rect 5080 11160 5132 11212
rect 1676 11092 1728 11144
rect 3884 11092 3936 11144
rect 4712 11092 4764 11144
rect 6736 11160 6788 11212
rect 7196 11296 7248 11348
rect 7564 11339 7616 11348
rect 7564 11305 7573 11339
rect 7573 11305 7607 11339
rect 7607 11305 7616 11339
rect 7564 11296 7616 11305
rect 8116 11296 8168 11348
rect 9404 11296 9456 11348
rect 10876 11296 10928 11348
rect 7104 11160 7156 11212
rect 15016 11228 15068 11280
rect 7840 11160 7892 11212
rect 8852 11160 8904 11212
rect 9588 11203 9640 11212
rect 9588 11169 9597 11203
rect 9597 11169 9631 11203
rect 9631 11169 9640 11203
rect 9588 11160 9640 11169
rect 9772 11203 9824 11212
rect 9772 11169 9781 11203
rect 9781 11169 9815 11203
rect 9815 11169 9824 11203
rect 9772 11160 9824 11169
rect 10876 11203 10928 11212
rect 10876 11169 10885 11203
rect 10885 11169 10919 11203
rect 10919 11169 10928 11203
rect 10876 11160 10928 11169
rect 8944 11092 8996 11144
rect 3792 11024 3844 11076
rect 2228 10956 2280 11008
rect 4068 10956 4120 11008
rect 4344 11024 4396 11076
rect 8852 11024 8904 11076
rect 9128 11067 9180 11076
rect 9128 11033 9137 11067
rect 9137 11033 9171 11067
rect 9171 11033 9180 11067
rect 9128 11024 9180 11033
rect 9864 11024 9916 11076
rect 15108 11067 15160 11076
rect 15108 11033 15117 11067
rect 15117 11033 15151 11067
rect 15151 11033 15160 11067
rect 15108 11024 15160 11033
rect 4712 10956 4764 11008
rect 5080 10956 5132 11008
rect 7012 10956 7064 11008
rect 9220 10956 9272 11008
rect 9312 10956 9364 11008
rect 12992 10956 13044 11008
rect 3481 10854 3533 10906
rect 3545 10854 3597 10906
rect 3609 10854 3661 10906
rect 3673 10854 3725 10906
rect 8480 10854 8532 10906
rect 8544 10854 8596 10906
rect 8608 10854 8660 10906
rect 8672 10854 8724 10906
rect 13478 10854 13530 10906
rect 13542 10854 13594 10906
rect 13606 10854 13658 10906
rect 13670 10854 13722 10906
rect 2136 10795 2188 10804
rect 2136 10761 2145 10795
rect 2145 10761 2179 10795
rect 2179 10761 2188 10795
rect 2136 10752 2188 10761
rect 2228 10752 2280 10804
rect 2964 10752 3016 10804
rect 4160 10752 4212 10804
rect 4620 10752 4672 10804
rect 3792 10684 3844 10736
rect 1952 10591 2004 10600
rect 1952 10557 1961 10591
rect 1961 10557 1995 10591
rect 1995 10557 2004 10591
rect 1952 10548 2004 10557
rect 3056 10548 3108 10600
rect 3240 10591 3292 10600
rect 3240 10557 3249 10591
rect 3249 10557 3283 10591
rect 3283 10557 3292 10591
rect 3240 10548 3292 10557
rect 2780 10480 2832 10532
rect 3424 10548 3476 10600
rect 3792 10548 3844 10600
rect 3884 10548 3936 10600
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4620 10616 4672 10668
rect 4068 10548 4120 10557
rect 4436 10591 4488 10600
rect 4436 10557 4445 10591
rect 4445 10557 4479 10591
rect 4479 10557 4488 10591
rect 4988 10795 5040 10804
rect 4988 10761 4997 10795
rect 4997 10761 5031 10795
rect 5031 10761 5040 10795
rect 8116 10795 8168 10804
rect 4988 10752 5040 10761
rect 8116 10761 8125 10795
rect 8125 10761 8159 10795
rect 8159 10761 8168 10795
rect 8116 10752 8168 10761
rect 7104 10684 7156 10736
rect 9588 10752 9640 10804
rect 9772 10752 9824 10804
rect 4436 10548 4488 10557
rect 5080 10591 5132 10600
rect 5080 10557 5089 10591
rect 5089 10557 5123 10591
rect 5123 10557 5132 10591
rect 5080 10548 5132 10557
rect 5264 10591 5316 10600
rect 5264 10557 5273 10591
rect 5273 10557 5307 10591
rect 5307 10557 5316 10591
rect 5264 10548 5316 10557
rect 9220 10659 9272 10668
rect 5448 10591 5500 10600
rect 5448 10557 5457 10591
rect 5457 10557 5491 10591
rect 5491 10557 5500 10591
rect 5448 10548 5500 10557
rect 7840 10548 7892 10600
rect 8392 10591 8444 10600
rect 8392 10557 8401 10591
rect 8401 10557 8435 10591
rect 8435 10557 8444 10591
rect 9220 10625 9229 10659
rect 9229 10625 9263 10659
rect 9263 10625 9272 10659
rect 9220 10616 9272 10625
rect 9864 10684 9916 10736
rect 9404 10616 9456 10668
rect 8392 10548 8444 10557
rect 8852 10523 8904 10532
rect 8852 10489 8861 10523
rect 8861 10489 8895 10523
rect 8895 10489 8904 10523
rect 8852 10480 8904 10489
rect 5816 10412 5868 10464
rect 9312 10548 9364 10600
rect 12072 10727 12124 10736
rect 12072 10693 12081 10727
rect 12081 10693 12115 10727
rect 12115 10693 12124 10727
rect 12072 10684 12124 10693
rect 12440 10616 12492 10668
rect 10508 10591 10560 10600
rect 10508 10557 10517 10591
rect 10517 10557 10551 10591
rect 10551 10557 10560 10591
rect 10508 10548 10560 10557
rect 11888 10591 11940 10600
rect 11888 10557 11897 10591
rect 11897 10557 11931 10591
rect 11931 10557 11940 10591
rect 11888 10548 11940 10557
rect 12256 10548 12308 10600
rect 15108 10548 15160 10600
rect 10876 10412 10928 10464
rect 11704 10455 11756 10464
rect 11704 10421 11713 10455
rect 11713 10421 11747 10455
rect 11747 10421 11756 10455
rect 11704 10412 11756 10421
rect 15016 10412 15068 10464
rect 5980 10310 6032 10362
rect 6044 10310 6096 10362
rect 6108 10310 6160 10362
rect 6172 10310 6224 10362
rect 10979 10310 11031 10362
rect 11043 10310 11095 10362
rect 11107 10310 11159 10362
rect 11171 10310 11223 10362
rect 3056 10208 3108 10260
rect 4436 10208 4488 10260
rect 5816 10208 5868 10260
rect 4160 10140 4212 10192
rect 5264 10140 5316 10192
rect 4068 10072 4120 10124
rect 4344 10072 4396 10124
rect 4712 10115 4764 10124
rect 4712 10081 4721 10115
rect 4721 10081 4755 10115
rect 4755 10081 4764 10115
rect 4712 10072 4764 10081
rect 4804 10115 4856 10124
rect 4804 10081 4813 10115
rect 4813 10081 4847 10115
rect 4847 10081 4856 10115
rect 5816 10115 5868 10124
rect 4804 10072 4856 10081
rect 5816 10081 5825 10115
rect 5825 10081 5859 10115
rect 5859 10081 5868 10115
rect 5816 10072 5868 10081
rect 3884 10004 3936 10056
rect 1952 9936 2004 9988
rect 9404 10208 9456 10260
rect 10232 10208 10284 10260
rect 12164 10208 12216 10260
rect 7748 10140 7800 10192
rect 12256 10140 12308 10192
rect 9956 10072 10008 10124
rect 10600 10072 10652 10124
rect 7840 9936 7892 9988
rect 9404 10004 9456 10056
rect 11980 10004 12032 10056
rect 12164 10047 12216 10056
rect 12164 10013 12173 10047
rect 12173 10013 12207 10047
rect 12207 10013 12216 10047
rect 12164 10004 12216 10013
rect 12532 10115 12584 10124
rect 12532 10081 12541 10115
rect 12541 10081 12575 10115
rect 12575 10081 12584 10115
rect 12532 10072 12584 10081
rect 12808 10115 12860 10124
rect 12808 10081 12817 10115
rect 12817 10081 12851 10115
rect 12851 10081 12860 10115
rect 12808 10072 12860 10081
rect 12992 10115 13044 10124
rect 12992 10081 13001 10115
rect 13001 10081 13035 10115
rect 13035 10081 13044 10115
rect 12992 10072 13044 10081
rect 15108 10140 15160 10192
rect 15016 10115 15068 10124
rect 15016 10081 15025 10115
rect 15025 10081 15059 10115
rect 15059 10081 15068 10115
rect 15752 10115 15804 10124
rect 15016 10072 15068 10081
rect 15752 10081 15761 10115
rect 15761 10081 15795 10115
rect 15795 10081 15804 10115
rect 15752 10072 15804 10081
rect 8852 9936 8904 9988
rect 11888 9936 11940 9988
rect 6368 9911 6420 9920
rect 6368 9877 6377 9911
rect 6377 9877 6411 9911
rect 6411 9877 6420 9911
rect 6368 9868 6420 9877
rect 7012 9868 7064 9920
rect 7288 9911 7340 9920
rect 7288 9877 7297 9911
rect 7297 9877 7331 9911
rect 7331 9877 7340 9911
rect 7288 9868 7340 9877
rect 10048 9911 10100 9920
rect 10048 9877 10057 9911
rect 10057 9877 10091 9911
rect 10091 9877 10100 9911
rect 10048 9868 10100 9877
rect 11796 9911 11848 9920
rect 11796 9877 11805 9911
rect 11805 9877 11839 9911
rect 11839 9877 11848 9911
rect 11796 9868 11848 9877
rect 11980 9868 12032 9920
rect 12808 9868 12860 9920
rect 12900 9911 12952 9920
rect 12900 9877 12909 9911
rect 12909 9877 12943 9911
rect 12943 9877 12952 9911
rect 13820 9911 13872 9920
rect 12900 9868 12952 9877
rect 13820 9877 13829 9911
rect 13829 9877 13863 9911
rect 13863 9877 13872 9911
rect 13820 9868 13872 9877
rect 15292 9868 15344 9920
rect 15568 9911 15620 9920
rect 15568 9877 15577 9911
rect 15577 9877 15611 9911
rect 15611 9877 15620 9911
rect 15568 9868 15620 9877
rect 3481 9766 3533 9818
rect 3545 9766 3597 9818
rect 3609 9766 3661 9818
rect 3673 9766 3725 9818
rect 8480 9766 8532 9818
rect 8544 9766 8596 9818
rect 8608 9766 8660 9818
rect 8672 9766 8724 9818
rect 13478 9766 13530 9818
rect 13542 9766 13594 9818
rect 13606 9766 13658 9818
rect 13670 9766 13722 9818
rect 2964 9707 3016 9716
rect 2964 9673 2973 9707
rect 2973 9673 3007 9707
rect 3007 9673 3016 9707
rect 2964 9664 3016 9673
rect 7840 9664 7892 9716
rect 10508 9664 10560 9716
rect 3240 9639 3292 9648
rect 3240 9605 3249 9639
rect 3249 9605 3283 9639
rect 3283 9605 3292 9639
rect 3240 9596 3292 9605
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 1952 9460 2004 9512
rect 6368 9528 6420 9580
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 3332 9503 3384 9512
rect 3332 9469 3341 9503
rect 3341 9469 3375 9503
rect 3375 9469 3384 9503
rect 3332 9460 3384 9469
rect 5724 9460 5776 9512
rect 9036 9460 9088 9512
rect 9680 9460 9732 9512
rect 15292 9503 15344 9512
rect 15292 9469 15301 9503
rect 15301 9469 15335 9503
rect 15335 9469 15344 9503
rect 15292 9460 15344 9469
rect 5816 9392 5868 9444
rect 7012 9392 7064 9444
rect 8116 9392 8168 9444
rect 8852 9392 8904 9444
rect 10600 9392 10652 9444
rect 15108 9435 15160 9444
rect 15108 9401 15117 9435
rect 15117 9401 15151 9435
rect 15151 9401 15160 9435
rect 15108 9392 15160 9401
rect 2228 9367 2280 9376
rect 2228 9333 2237 9367
rect 2237 9333 2271 9367
rect 2271 9333 2280 9367
rect 2228 9324 2280 9333
rect 2504 9367 2556 9376
rect 2504 9333 2513 9367
rect 2513 9333 2547 9367
rect 2547 9333 2556 9367
rect 2504 9324 2556 9333
rect 9772 9367 9824 9376
rect 9772 9333 9781 9367
rect 9781 9333 9815 9367
rect 9815 9333 9824 9367
rect 9772 9324 9824 9333
rect 5980 9222 6032 9274
rect 6044 9222 6096 9274
rect 6108 9222 6160 9274
rect 6172 9222 6224 9274
rect 10979 9222 11031 9274
rect 11043 9222 11095 9274
rect 11107 9222 11159 9274
rect 11171 9222 11223 9274
rect 2504 9120 2556 9172
rect 2228 9052 2280 9104
rect 8116 9120 8168 9172
rect 5816 9052 5868 9104
rect 6920 9052 6972 9104
rect 4068 9027 4120 9036
rect 4068 8993 4077 9027
rect 4077 8993 4111 9027
rect 4111 8993 4120 9027
rect 4068 8984 4120 8993
rect 4436 8984 4488 9036
rect 4712 9027 4764 9036
rect 4712 8993 4721 9027
rect 4721 8993 4755 9027
rect 4755 8993 4764 9027
rect 4712 8984 4764 8993
rect 5356 8984 5408 9036
rect 1676 8916 1728 8968
rect 5724 8916 5776 8968
rect 3332 8780 3384 8832
rect 4160 8780 4212 8832
rect 4620 8780 4672 8832
rect 5264 8823 5316 8832
rect 5264 8789 5273 8823
rect 5273 8789 5307 8823
rect 5307 8789 5316 8823
rect 5264 8780 5316 8789
rect 5816 8823 5868 8832
rect 5816 8789 5825 8823
rect 5825 8789 5859 8823
rect 5859 8789 5868 8823
rect 5816 8780 5868 8789
rect 6828 8984 6880 9036
rect 9128 9027 9180 9036
rect 9128 8993 9137 9027
rect 9137 8993 9171 9027
rect 9171 8993 9180 9027
rect 9128 8984 9180 8993
rect 9680 9120 9732 9172
rect 10600 9163 10652 9172
rect 10600 9129 10609 9163
rect 10609 9129 10643 9163
rect 10643 9129 10652 9163
rect 10600 9120 10652 9129
rect 12900 9052 12952 9104
rect 10048 8984 10100 9036
rect 12532 9027 12584 9036
rect 12532 8993 12541 9027
rect 12541 8993 12575 9027
rect 12575 8993 12584 9027
rect 12532 8984 12584 8993
rect 13176 8984 13228 9036
rect 13360 8916 13412 8968
rect 9772 8891 9824 8900
rect 9772 8857 9781 8891
rect 9781 8857 9815 8891
rect 9815 8857 9824 8891
rect 9772 8848 9824 8857
rect 6092 8780 6144 8832
rect 13268 8823 13320 8832
rect 13268 8789 13277 8823
rect 13277 8789 13311 8823
rect 13311 8789 13320 8823
rect 13268 8780 13320 8789
rect 14188 8780 14240 8832
rect 3481 8678 3533 8730
rect 3545 8678 3597 8730
rect 3609 8678 3661 8730
rect 3673 8678 3725 8730
rect 8480 8678 8532 8730
rect 8544 8678 8596 8730
rect 8608 8678 8660 8730
rect 8672 8678 8724 8730
rect 13478 8678 13530 8730
rect 13542 8678 13594 8730
rect 13606 8678 13658 8730
rect 13670 8678 13722 8730
rect 4712 8619 4764 8628
rect 4344 8508 4396 8560
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 4712 8585 4721 8619
rect 4721 8585 4755 8619
rect 4755 8585 4764 8619
rect 4712 8576 4764 8585
rect 4804 8508 4856 8560
rect 10324 8576 10376 8628
rect 10600 8576 10652 8628
rect 5356 8508 5408 8560
rect 5816 8440 5868 8492
rect 2228 8415 2280 8424
rect 2228 8381 2237 8415
rect 2237 8381 2271 8415
rect 2271 8381 2280 8415
rect 2228 8372 2280 8381
rect 2320 8372 2372 8424
rect 4252 8415 4304 8424
rect 4252 8381 4261 8415
rect 4261 8381 4295 8415
rect 4295 8381 4304 8415
rect 4436 8415 4488 8424
rect 4252 8372 4304 8381
rect 4436 8381 4445 8415
rect 4445 8381 4479 8415
rect 4479 8381 4488 8415
rect 4436 8372 4488 8381
rect 5172 8415 5224 8424
rect 4620 8304 4672 8356
rect 5172 8381 5181 8415
rect 5181 8381 5215 8415
rect 5215 8381 5224 8415
rect 5172 8372 5224 8381
rect 5264 8415 5316 8424
rect 5264 8381 5273 8415
rect 5273 8381 5307 8415
rect 5307 8381 5316 8415
rect 5448 8415 5500 8424
rect 5264 8372 5316 8381
rect 5448 8381 5457 8415
rect 5457 8381 5491 8415
rect 5491 8381 5500 8415
rect 5448 8372 5500 8381
rect 6644 8508 6696 8560
rect 13084 8551 13136 8560
rect 13084 8517 13093 8551
rect 13093 8517 13127 8551
rect 13127 8517 13136 8551
rect 13084 8508 13136 8517
rect 13360 8508 13412 8560
rect 6828 8440 6880 8492
rect 6092 8415 6144 8424
rect 6092 8381 6101 8415
rect 6101 8381 6135 8415
rect 6135 8381 6144 8415
rect 6092 8372 6144 8381
rect 6552 8415 6604 8424
rect 6552 8381 6561 8415
rect 6561 8381 6595 8415
rect 6595 8381 6604 8415
rect 6552 8372 6604 8381
rect 6644 8415 6696 8424
rect 6644 8381 6653 8415
rect 6653 8381 6687 8415
rect 6687 8381 6696 8415
rect 6920 8415 6972 8424
rect 6644 8372 6696 8381
rect 6920 8381 6929 8415
rect 6929 8381 6963 8415
rect 6963 8381 6972 8415
rect 6920 8372 6972 8381
rect 7288 8440 7340 8492
rect 9680 8440 9732 8492
rect 8668 8372 8720 8424
rect 10048 8372 10100 8424
rect 12532 8440 12584 8492
rect 11796 8415 11848 8424
rect 11796 8381 11805 8415
rect 11805 8381 11839 8415
rect 11839 8381 11848 8415
rect 11796 8372 11848 8381
rect 13176 8372 13228 8424
rect 13636 8372 13688 8424
rect 14188 8415 14240 8424
rect 14188 8381 14197 8415
rect 14197 8381 14231 8415
rect 14231 8381 14240 8415
rect 14188 8372 14240 8381
rect 14556 8372 14608 8424
rect 15108 8372 15160 8424
rect 8392 8347 8444 8356
rect 8392 8313 8401 8347
rect 8401 8313 8435 8347
rect 8435 8313 8444 8347
rect 8392 8304 8444 8313
rect 13452 8347 13504 8356
rect 13452 8313 13461 8347
rect 13461 8313 13495 8347
rect 13495 8313 13504 8347
rect 13452 8304 13504 8313
rect 4344 8236 4396 8288
rect 5448 8236 5500 8288
rect 7748 8279 7800 8288
rect 7748 8245 7757 8279
rect 7757 8245 7791 8279
rect 7791 8245 7800 8279
rect 7748 8236 7800 8245
rect 14740 8236 14792 8288
rect 5980 8134 6032 8186
rect 6044 8134 6096 8186
rect 6108 8134 6160 8186
rect 6172 8134 6224 8186
rect 10979 8134 11031 8186
rect 11043 8134 11095 8186
rect 11107 8134 11159 8186
rect 11171 8134 11223 8186
rect 2044 7964 2096 8016
rect 4252 8007 4304 8016
rect 4252 7973 4261 8007
rect 4261 7973 4295 8007
rect 4295 7973 4304 8007
rect 4252 7964 4304 7973
rect 2320 7939 2372 7948
rect 2320 7905 2329 7939
rect 2329 7905 2363 7939
rect 2363 7905 2372 7939
rect 2320 7896 2372 7905
rect 2688 7939 2740 7948
rect 2688 7905 2697 7939
rect 2697 7905 2731 7939
rect 2731 7905 2740 7939
rect 2688 7896 2740 7905
rect 3148 7939 3200 7948
rect 3148 7905 3157 7939
rect 3157 7905 3191 7939
rect 3191 7905 3200 7939
rect 3148 7896 3200 7905
rect 3332 7939 3384 7948
rect 3332 7905 3341 7939
rect 3341 7905 3375 7939
rect 3375 7905 3384 7939
rect 3332 7896 3384 7905
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 5356 7964 5408 8016
rect 7748 8007 7800 8016
rect 7748 7973 7757 8007
rect 7757 7973 7791 8007
rect 7791 7973 7800 8007
rect 7748 7964 7800 7973
rect 8668 8075 8720 8084
rect 8668 8041 8677 8075
rect 8677 8041 8711 8075
rect 8711 8041 8720 8075
rect 9680 8075 9732 8084
rect 8668 8032 8720 8041
rect 9680 8041 9689 8075
rect 9689 8041 9723 8075
rect 9723 8041 9732 8075
rect 9680 8032 9732 8041
rect 13452 8075 13504 8084
rect 13452 8041 13461 8075
rect 13461 8041 13495 8075
rect 13495 8041 13504 8075
rect 13452 8032 13504 8041
rect 14740 8075 14792 8084
rect 14740 8041 14749 8075
rect 14749 8041 14783 8075
rect 14783 8041 14792 8075
rect 14740 8032 14792 8041
rect 8944 7964 8996 8016
rect 5080 7939 5132 7948
rect 5080 7905 5089 7939
rect 5089 7905 5123 7939
rect 5123 7905 5132 7939
rect 5080 7896 5132 7905
rect 5632 7939 5684 7948
rect 5632 7905 5641 7939
rect 5641 7905 5675 7939
rect 5675 7905 5684 7939
rect 5632 7896 5684 7905
rect 5816 7939 5868 7948
rect 5816 7905 5825 7939
rect 5825 7905 5859 7939
rect 5859 7905 5868 7939
rect 5816 7896 5868 7905
rect 7288 7939 7340 7948
rect 7288 7905 7297 7939
rect 7297 7905 7331 7939
rect 7331 7905 7340 7939
rect 7288 7896 7340 7905
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 2596 7871 2648 7880
rect 2596 7837 2605 7871
rect 2605 7837 2639 7871
rect 2639 7837 2648 7871
rect 2596 7828 2648 7837
rect 8116 7828 8168 7880
rect 8392 7896 8444 7948
rect 8852 7939 8904 7948
rect 8852 7905 8861 7939
rect 8861 7905 8895 7939
rect 8895 7905 8904 7939
rect 8852 7896 8904 7905
rect 11796 7939 11848 7948
rect 11796 7905 11805 7939
rect 11805 7905 11839 7939
rect 11839 7905 11848 7939
rect 11796 7896 11848 7905
rect 13268 7939 13320 7948
rect 13268 7905 13277 7939
rect 13277 7905 13311 7939
rect 13311 7905 13320 7939
rect 13268 7896 13320 7905
rect 13636 7939 13688 7948
rect 13636 7905 13645 7939
rect 13645 7905 13679 7939
rect 13679 7905 13688 7939
rect 13636 7896 13688 7905
rect 13084 7871 13136 7880
rect 13084 7837 13093 7871
rect 13093 7837 13127 7871
rect 13127 7837 13136 7871
rect 13084 7828 13136 7837
rect 4436 7760 4488 7812
rect 14740 7896 14792 7948
rect 15016 7692 15068 7744
rect 3481 7590 3533 7642
rect 3545 7590 3597 7642
rect 3609 7590 3661 7642
rect 3673 7590 3725 7642
rect 8480 7590 8532 7642
rect 8544 7590 8596 7642
rect 8608 7590 8660 7642
rect 8672 7590 8724 7642
rect 13478 7590 13530 7642
rect 13542 7590 13594 7642
rect 13606 7590 13658 7642
rect 13670 7590 13722 7642
rect 2320 7488 2372 7540
rect 5816 7488 5868 7540
rect 8944 7488 8996 7540
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 3148 7420 3200 7472
rect 15016 7463 15068 7472
rect 15016 7429 15025 7463
rect 15025 7429 15059 7463
rect 15059 7429 15068 7463
rect 15016 7420 15068 7429
rect 2688 7352 2740 7404
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 3148 7327 3200 7336
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3148 7284 3200 7293
rect 4528 7284 4580 7336
rect 5448 7284 5500 7336
rect 8116 7284 8168 7336
rect 8852 7284 8904 7336
rect 9588 7284 9640 7336
rect 10876 7284 10928 7336
rect 13084 7284 13136 7336
rect 13820 7284 13872 7336
rect 14556 7327 14608 7336
rect 14556 7293 14565 7327
rect 14565 7293 14599 7327
rect 14599 7293 14608 7327
rect 14556 7284 14608 7293
rect 2596 7216 2648 7268
rect 3056 7259 3108 7268
rect 3056 7225 3065 7259
rect 3065 7225 3099 7259
rect 3099 7225 3108 7259
rect 3056 7216 3108 7225
rect 14740 7216 14792 7268
rect 3332 7148 3384 7200
rect 10692 7148 10744 7200
rect 11428 7191 11480 7200
rect 11428 7157 11437 7191
rect 11437 7157 11471 7191
rect 11471 7157 11480 7191
rect 11428 7148 11480 7157
rect 5980 7046 6032 7098
rect 6044 7046 6096 7098
rect 6108 7046 6160 7098
rect 6172 7046 6224 7098
rect 10979 7046 11031 7098
rect 11043 7046 11095 7098
rect 11107 7046 11159 7098
rect 11171 7046 11223 7098
rect 3332 6944 3384 6996
rect 3976 6944 4028 6996
rect 6552 6987 6604 6996
rect 6552 6953 6561 6987
rect 6561 6953 6595 6987
rect 6595 6953 6604 6987
rect 6552 6944 6604 6953
rect 5080 6876 5132 6928
rect 3884 6672 3936 6724
rect 4528 6783 4580 6792
rect 4528 6749 4537 6783
rect 4537 6749 4571 6783
rect 4571 6749 4580 6783
rect 4528 6740 4580 6749
rect 4804 6808 4856 6860
rect 4988 6808 5040 6860
rect 5540 6808 5592 6860
rect 9588 6919 9640 6928
rect 5172 6715 5224 6724
rect 5172 6681 5181 6715
rect 5181 6681 5215 6715
rect 5215 6681 5224 6715
rect 5172 6672 5224 6681
rect 6184 6851 6236 6860
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 9588 6885 9597 6919
rect 9597 6885 9631 6919
rect 9631 6885 9640 6919
rect 9588 6876 9640 6885
rect 10692 6919 10744 6928
rect 10692 6885 10701 6919
rect 10701 6885 10735 6919
rect 10735 6885 10744 6919
rect 10692 6876 10744 6885
rect 6736 6783 6788 6792
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 10416 6808 10468 6860
rect 10876 6808 10928 6860
rect 11428 6808 11480 6860
rect 11704 6808 11756 6860
rect 13176 6851 13228 6860
rect 13176 6817 13185 6851
rect 13185 6817 13219 6851
rect 13219 6817 13228 6851
rect 13176 6808 13228 6817
rect 6828 6672 6880 6724
rect 12348 6740 12400 6792
rect 12900 6783 12952 6792
rect 12900 6749 12909 6783
rect 12909 6749 12943 6783
rect 12943 6749 12952 6783
rect 12900 6740 12952 6749
rect 7748 6672 7800 6724
rect 7564 6604 7616 6656
rect 3481 6502 3533 6554
rect 3545 6502 3597 6554
rect 3609 6502 3661 6554
rect 3673 6502 3725 6554
rect 8480 6502 8532 6554
rect 8544 6502 8596 6554
rect 8608 6502 8660 6554
rect 8672 6502 8724 6554
rect 13478 6502 13530 6554
rect 13542 6502 13594 6554
rect 13606 6502 13658 6554
rect 13670 6502 13722 6554
rect 4528 6400 4580 6452
rect 5080 6400 5132 6452
rect 5724 6400 5776 6452
rect 6184 6400 6236 6452
rect 7564 6443 7616 6452
rect 7564 6409 7573 6443
rect 7573 6409 7607 6443
rect 7607 6409 7616 6443
rect 7564 6400 7616 6409
rect 7748 6443 7800 6452
rect 7748 6409 7757 6443
rect 7757 6409 7791 6443
rect 7791 6409 7800 6443
rect 7748 6400 7800 6409
rect 1952 6196 2004 6248
rect 2504 6239 2556 6248
rect 2504 6205 2513 6239
rect 2513 6205 2547 6239
rect 2547 6205 2556 6239
rect 2504 6196 2556 6205
rect 3056 6264 3108 6316
rect 5632 6332 5684 6384
rect 5816 6332 5868 6384
rect 3884 6239 3936 6248
rect 2780 6171 2832 6180
rect 2780 6137 2789 6171
rect 2789 6137 2823 6171
rect 2823 6137 2832 6171
rect 2780 6128 2832 6137
rect 3148 6128 3200 6180
rect 3884 6205 3893 6239
rect 3893 6205 3927 6239
rect 3927 6205 3936 6239
rect 3884 6196 3936 6205
rect 3976 6196 4028 6248
rect 5080 6239 5132 6248
rect 5080 6205 5089 6239
rect 5089 6205 5123 6239
rect 5123 6205 5132 6239
rect 5080 6196 5132 6205
rect 5448 6239 5500 6248
rect 4252 6128 4304 6180
rect 5448 6205 5457 6239
rect 5457 6205 5491 6239
rect 5491 6205 5500 6239
rect 5448 6196 5500 6205
rect 5540 6128 5592 6180
rect 5724 6239 5776 6248
rect 5724 6205 5733 6239
rect 5733 6205 5767 6239
rect 5767 6205 5776 6239
rect 5724 6196 5776 6205
rect 7932 6332 7984 6384
rect 13176 6307 13228 6316
rect 1860 6060 1912 6112
rect 2872 6060 2924 6112
rect 13176 6273 13185 6307
rect 13185 6273 13219 6307
rect 13219 6273 13228 6307
rect 13176 6264 13228 6273
rect 8116 6239 8168 6248
rect 8116 6205 8125 6239
rect 8125 6205 8159 6239
rect 8159 6205 8168 6239
rect 8116 6196 8168 6205
rect 9588 6239 9640 6248
rect 7932 6103 7984 6112
rect 7932 6069 7941 6103
rect 7941 6069 7975 6103
rect 7975 6069 7984 6103
rect 9588 6205 9597 6239
rect 9597 6205 9631 6239
rect 9631 6205 9640 6239
rect 9588 6196 9640 6205
rect 11704 6239 11756 6248
rect 11704 6205 11713 6239
rect 11713 6205 11747 6239
rect 11747 6205 11756 6239
rect 11704 6196 11756 6205
rect 12900 6239 12952 6248
rect 12900 6205 12909 6239
rect 12909 6205 12943 6239
rect 12943 6205 12952 6239
rect 12900 6196 12952 6205
rect 12348 6128 12400 6180
rect 13084 6171 13136 6180
rect 13084 6137 13093 6171
rect 13093 6137 13127 6171
rect 13127 6137 13136 6171
rect 13084 6128 13136 6137
rect 7932 6060 7984 6069
rect 9864 6060 9916 6112
rect 13820 6103 13872 6112
rect 13820 6069 13829 6103
rect 13829 6069 13863 6103
rect 13863 6069 13872 6103
rect 13820 6060 13872 6069
rect 5980 5958 6032 6010
rect 6044 5958 6096 6010
rect 6108 5958 6160 6010
rect 6172 5958 6224 6010
rect 10979 5958 11031 6010
rect 11043 5958 11095 6010
rect 11107 5958 11159 6010
rect 11171 5958 11223 6010
rect 2780 5856 2832 5908
rect 6736 5856 6788 5908
rect 1860 5788 1912 5840
rect 2872 5831 2924 5840
rect 2872 5797 2881 5831
rect 2881 5797 2915 5831
rect 2915 5797 2924 5831
rect 2872 5788 2924 5797
rect 3240 5788 3292 5840
rect 3976 5788 4028 5840
rect 5632 5788 5684 5840
rect 8116 5788 8168 5840
rect 9864 5788 9916 5840
rect 3792 5720 3844 5772
rect 4252 5763 4304 5772
rect 1676 5652 1728 5704
rect 3976 5652 4028 5704
rect 4252 5729 4261 5763
rect 4261 5729 4295 5763
rect 4295 5729 4304 5763
rect 4252 5720 4304 5729
rect 6276 5763 6328 5772
rect 6276 5729 6285 5763
rect 6285 5729 6319 5763
rect 6319 5729 6328 5763
rect 6276 5720 6328 5729
rect 6736 5720 6788 5772
rect 8300 5763 8352 5772
rect 8300 5729 8309 5763
rect 8309 5729 8343 5763
rect 8343 5729 8352 5763
rect 8300 5720 8352 5729
rect 6460 5652 6512 5704
rect 7932 5652 7984 5704
rect 8208 5652 8260 5704
rect 4988 5584 5040 5636
rect 7012 5584 7064 5636
rect 11060 5720 11112 5772
rect 12348 5763 12400 5772
rect 12348 5729 12357 5763
rect 12357 5729 12391 5763
rect 12391 5729 12400 5763
rect 12348 5720 12400 5729
rect 13820 5720 13872 5772
rect 11336 5652 11388 5704
rect 4712 5516 4764 5568
rect 12532 5584 12584 5636
rect 9404 5516 9456 5568
rect 10784 5516 10836 5568
rect 11244 5559 11296 5568
rect 11244 5525 11253 5559
rect 11253 5525 11287 5559
rect 11287 5525 11296 5559
rect 11244 5516 11296 5525
rect 14464 5559 14516 5568
rect 14464 5525 14473 5559
rect 14473 5525 14507 5559
rect 14507 5525 14516 5559
rect 14464 5516 14516 5525
rect 3481 5414 3533 5466
rect 3545 5414 3597 5466
rect 3609 5414 3661 5466
rect 3673 5414 3725 5466
rect 8480 5414 8532 5466
rect 8544 5414 8596 5466
rect 8608 5414 8660 5466
rect 8672 5414 8724 5466
rect 13478 5414 13530 5466
rect 13542 5414 13594 5466
rect 13606 5414 13658 5466
rect 13670 5414 13722 5466
rect 3240 5355 3292 5364
rect 3240 5321 3249 5355
rect 3249 5321 3283 5355
rect 3283 5321 3292 5355
rect 3240 5312 3292 5321
rect 6276 5312 6328 5364
rect 9036 5312 9088 5364
rect 5172 5244 5224 5296
rect 8760 5244 8812 5296
rect 10324 5244 10376 5296
rect 4712 5219 4764 5228
rect 4712 5185 4721 5219
rect 4721 5185 4755 5219
rect 4755 5185 4764 5219
rect 4712 5176 4764 5185
rect 4988 5219 5040 5228
rect 4988 5185 4997 5219
rect 4997 5185 5031 5219
rect 5031 5185 5040 5219
rect 4988 5176 5040 5185
rect 6736 5176 6788 5228
rect 9312 5176 9364 5228
rect 10876 5176 10928 5228
rect 4160 5040 4212 5092
rect 5632 5040 5684 5092
rect 6460 5108 6512 5160
rect 8300 5108 8352 5160
rect 9036 5151 9088 5160
rect 9036 5117 9045 5151
rect 9045 5117 9079 5151
rect 9079 5117 9088 5151
rect 9036 5108 9088 5117
rect 9404 5151 9456 5160
rect 9404 5117 9413 5151
rect 9413 5117 9447 5151
rect 9447 5117 9456 5151
rect 9404 5108 9456 5117
rect 9588 5108 9640 5160
rect 9864 5108 9916 5160
rect 10784 5108 10836 5160
rect 9128 5040 9180 5092
rect 9312 5083 9364 5092
rect 9312 5049 9321 5083
rect 9321 5049 9355 5083
rect 9355 5049 9364 5083
rect 9312 5040 9364 5049
rect 5540 5015 5592 5024
rect 5540 4981 5549 5015
rect 5549 4981 5583 5015
rect 5583 4981 5592 5015
rect 5540 4972 5592 4981
rect 6276 4972 6328 5024
rect 6736 4972 6788 5024
rect 7932 4972 7984 5024
rect 9588 5015 9640 5024
rect 9588 4981 9597 5015
rect 9597 4981 9631 5015
rect 9631 4981 9640 5015
rect 9588 4972 9640 4981
rect 10324 5015 10376 5024
rect 10324 4981 10333 5015
rect 10333 4981 10367 5015
rect 10367 4981 10376 5015
rect 10324 4972 10376 4981
rect 11244 5312 11296 5364
rect 12348 5219 12400 5228
rect 12348 5185 12357 5219
rect 12357 5185 12391 5219
rect 12391 5185 12400 5219
rect 12348 5176 12400 5185
rect 11888 5108 11940 5160
rect 12164 5151 12216 5160
rect 12164 5117 12173 5151
rect 12173 5117 12207 5151
rect 12207 5117 12216 5151
rect 12164 5108 12216 5117
rect 15568 5312 15620 5364
rect 13728 5176 13780 5228
rect 14464 5176 14516 5228
rect 12532 5108 12584 5160
rect 13176 5151 13228 5160
rect 13176 5117 13185 5151
rect 13185 5117 13219 5151
rect 13219 5117 13228 5151
rect 13176 5108 13228 5117
rect 11428 5040 11480 5092
rect 11612 5040 11664 5092
rect 14096 5083 14148 5092
rect 14096 5049 14105 5083
rect 14105 5049 14139 5083
rect 14139 5049 14148 5083
rect 14096 5040 14148 5049
rect 14188 5040 14240 5092
rect 11704 4972 11756 5024
rect 12992 5015 13044 5024
rect 12992 4981 13001 5015
rect 13001 4981 13035 5015
rect 13035 4981 13044 5015
rect 12992 4972 13044 4981
rect 15568 5015 15620 5024
rect 15568 4981 15577 5015
rect 15577 4981 15611 5015
rect 15611 4981 15620 5015
rect 15568 4972 15620 4981
rect 5980 4870 6032 4922
rect 6044 4870 6096 4922
rect 6108 4870 6160 4922
rect 6172 4870 6224 4922
rect 10979 4870 11031 4922
rect 11043 4870 11095 4922
rect 11107 4870 11159 4922
rect 11171 4870 11223 4922
rect 2596 4811 2648 4820
rect 2596 4777 2605 4811
rect 2605 4777 2639 4811
rect 2639 4777 2648 4811
rect 2596 4768 2648 4777
rect 4160 4811 4212 4820
rect 4160 4777 4169 4811
rect 4169 4777 4203 4811
rect 4203 4777 4212 4811
rect 4160 4768 4212 4777
rect 5816 4768 5868 4820
rect 9312 4768 9364 4820
rect 9588 4768 9640 4820
rect 2504 4700 2556 4752
rect 3792 4700 3844 4752
rect 4528 4700 4580 4752
rect 4988 4700 5040 4752
rect 7932 4700 7984 4752
rect 10324 4700 10376 4752
rect 14188 4811 14240 4820
rect 10968 4700 11020 4752
rect 1952 4632 2004 4684
rect 2780 4632 2832 4684
rect 3056 4632 3108 4684
rect 5448 4675 5500 4684
rect 5448 4641 5457 4675
rect 5457 4641 5491 4675
rect 5491 4641 5500 4675
rect 5448 4632 5500 4641
rect 5632 4632 5684 4684
rect 6920 4675 6972 4684
rect 6920 4641 6929 4675
rect 6929 4641 6963 4675
rect 6963 4641 6972 4675
rect 6920 4632 6972 4641
rect 11428 4700 11480 4752
rect 14188 4777 14197 4811
rect 14197 4777 14231 4811
rect 14231 4777 14240 4811
rect 14188 4768 14240 4777
rect 12992 4700 13044 4752
rect 13176 4700 13228 4752
rect 11612 4675 11664 4684
rect 5172 4564 5224 4616
rect 5356 4607 5408 4616
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 7196 4607 7248 4616
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7196 4564 7248 4573
rect 7288 4564 7340 4616
rect 8208 4564 8260 4616
rect 11152 4607 11204 4616
rect 11152 4573 11161 4607
rect 11161 4573 11195 4607
rect 11195 4573 11204 4607
rect 11152 4564 11204 4573
rect 11612 4641 11621 4675
rect 11621 4641 11655 4675
rect 11655 4641 11664 4675
rect 11612 4632 11664 4641
rect 11704 4675 11756 4684
rect 11704 4641 11713 4675
rect 11713 4641 11747 4675
rect 11747 4641 11756 4675
rect 11704 4632 11756 4641
rect 13728 4675 13780 4684
rect 13728 4641 13737 4675
rect 13737 4641 13771 4675
rect 13771 4641 13780 4675
rect 13728 4632 13780 4641
rect 14096 4632 14148 4684
rect 12072 4564 12124 4616
rect 8760 4496 8812 4548
rect 9864 4496 9916 4548
rect 15568 4675 15620 4684
rect 15568 4641 15577 4675
rect 15577 4641 15611 4675
rect 15611 4641 15620 4675
rect 15568 4632 15620 4641
rect 15752 4496 15804 4548
rect 2228 4471 2280 4480
rect 2228 4437 2237 4471
rect 2237 4437 2271 4471
rect 2271 4437 2280 4471
rect 2228 4428 2280 4437
rect 2412 4471 2464 4480
rect 2412 4437 2421 4471
rect 2421 4437 2455 4471
rect 2455 4437 2464 4471
rect 2412 4428 2464 4437
rect 4528 4428 4580 4480
rect 8300 4428 8352 4480
rect 12072 4428 12124 4480
rect 3481 4326 3533 4378
rect 3545 4326 3597 4378
rect 3609 4326 3661 4378
rect 3673 4326 3725 4378
rect 8480 4326 8532 4378
rect 8544 4326 8596 4378
rect 8608 4326 8660 4378
rect 8672 4326 8724 4378
rect 13478 4326 13530 4378
rect 13542 4326 13594 4378
rect 13606 4326 13658 4378
rect 13670 4326 13722 4378
rect 2412 4224 2464 4276
rect 3056 4224 3108 4276
rect 3240 4224 3292 4276
rect 11152 4224 11204 4276
rect 12440 4224 12492 4276
rect 13820 4224 13872 4276
rect 15752 4267 15804 4276
rect 15752 4233 15761 4267
rect 15761 4233 15795 4267
rect 15795 4233 15804 4267
rect 15752 4224 15804 4233
rect 5448 4156 5500 4208
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 1676 4088 1728 4140
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 5356 4020 5408 4072
rect 11612 4088 11664 4140
rect 13820 4088 13872 4140
rect 2228 3952 2280 4004
rect 6644 4020 6696 4072
rect 7288 4063 7340 4072
rect 7288 4029 7297 4063
rect 7297 4029 7331 4063
rect 7331 4029 7340 4063
rect 7288 4020 7340 4029
rect 11704 4063 11756 4072
rect 11704 4029 11713 4063
rect 11713 4029 11747 4063
rect 11747 4029 11756 4063
rect 11704 4020 11756 4029
rect 11980 4063 12032 4072
rect 11980 4029 11989 4063
rect 11989 4029 12023 4063
rect 12023 4029 12032 4063
rect 11980 4020 12032 4029
rect 12072 4063 12124 4072
rect 12072 4029 12081 4063
rect 12081 4029 12115 4063
rect 12115 4029 12124 4063
rect 12072 4020 12124 4029
rect 6368 3952 6420 4004
rect 6276 3884 6328 3936
rect 9312 3952 9364 4004
rect 11888 3995 11940 4004
rect 11888 3961 11897 3995
rect 11897 3961 11931 3995
rect 11931 3961 11940 3995
rect 11888 3952 11940 3961
rect 14280 3995 14332 4004
rect 14280 3961 14289 3995
rect 14289 3961 14323 3995
rect 14323 3961 14332 3995
rect 14280 3952 14332 3961
rect 14924 3952 14976 4004
rect 6552 3884 6604 3936
rect 13544 3884 13596 3936
rect 5980 3782 6032 3834
rect 6044 3782 6096 3834
rect 6108 3782 6160 3834
rect 6172 3782 6224 3834
rect 10979 3782 11031 3834
rect 11043 3782 11095 3834
rect 11107 3782 11159 3834
rect 11171 3782 11223 3834
rect 3240 3680 3292 3732
rect 3976 3655 4028 3664
rect 3976 3621 3985 3655
rect 3985 3621 4019 3655
rect 4019 3621 4028 3655
rect 3976 3612 4028 3621
rect 3332 3544 3384 3596
rect 4252 3544 4304 3596
rect 7012 3680 7064 3732
rect 6368 3612 6420 3664
rect 11980 3680 12032 3732
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 6828 3587 6880 3596
rect 6828 3553 6837 3587
rect 6837 3553 6871 3587
rect 6871 3553 6880 3587
rect 6828 3544 6880 3553
rect 7012 3544 7064 3596
rect 9220 3612 9272 3664
rect 11520 3612 11572 3664
rect 12532 3612 12584 3664
rect 13544 3655 13596 3664
rect 13544 3621 13553 3655
rect 13553 3621 13587 3655
rect 13587 3621 13596 3655
rect 13544 3612 13596 3621
rect 9036 3544 9088 3596
rect 9312 3587 9364 3596
rect 9312 3553 9321 3587
rect 9321 3553 9355 3587
rect 9355 3553 9364 3587
rect 9312 3544 9364 3553
rect 9496 3587 9548 3596
rect 9496 3553 9505 3587
rect 9505 3553 9539 3587
rect 9539 3553 9548 3587
rect 9496 3544 9548 3553
rect 9864 3544 9916 3596
rect 10048 3587 10100 3596
rect 10048 3553 10057 3587
rect 10057 3553 10091 3587
rect 10091 3553 10100 3587
rect 10048 3544 10100 3553
rect 13820 3587 13872 3596
rect 13820 3553 13829 3587
rect 13829 3553 13863 3587
rect 13863 3553 13872 3587
rect 13820 3544 13872 3553
rect 6368 3476 6420 3528
rect 6644 3519 6696 3528
rect 6644 3485 6653 3519
rect 6653 3485 6687 3519
rect 6687 3485 6696 3519
rect 6644 3476 6696 3485
rect 7104 3476 7156 3528
rect 7380 3519 7432 3528
rect 7380 3485 7389 3519
rect 7389 3485 7423 3519
rect 7423 3485 7432 3519
rect 7380 3476 7432 3485
rect 4252 3408 4304 3460
rect 7196 3408 7248 3460
rect 7656 3476 7708 3528
rect 7012 3383 7064 3392
rect 7012 3349 7021 3383
rect 7021 3349 7055 3383
rect 7055 3349 7064 3383
rect 7012 3340 7064 3349
rect 7288 3340 7340 3392
rect 9680 3383 9732 3392
rect 9680 3349 9689 3383
rect 9689 3349 9723 3383
rect 9723 3349 9732 3383
rect 9680 3340 9732 3349
rect 9772 3340 9824 3392
rect 11152 3476 11204 3528
rect 11888 3476 11940 3528
rect 11060 3340 11112 3392
rect 3481 3238 3533 3290
rect 3545 3238 3597 3290
rect 3609 3238 3661 3290
rect 3673 3238 3725 3290
rect 8480 3238 8532 3290
rect 8544 3238 8596 3290
rect 8608 3238 8660 3290
rect 8672 3238 8724 3290
rect 13478 3238 13530 3290
rect 13542 3238 13594 3290
rect 13606 3238 13658 3290
rect 13670 3238 13722 3290
rect 5080 3136 5132 3188
rect 7104 3136 7156 3188
rect 9128 3179 9180 3188
rect 9128 3145 9137 3179
rect 9137 3145 9171 3179
rect 9171 3145 9180 3179
rect 9128 3136 9180 3145
rect 9220 3136 9272 3188
rect 11152 3179 11204 3188
rect 11152 3145 11161 3179
rect 11161 3145 11195 3179
rect 11195 3145 11204 3179
rect 11152 3136 11204 3145
rect 14280 3136 14332 3188
rect 14924 3179 14976 3188
rect 14924 3145 14933 3179
rect 14933 3145 14967 3179
rect 14967 3145 14976 3179
rect 14924 3136 14976 3145
rect 3240 3068 3292 3120
rect 2780 3000 2832 3052
rect 480 2932 532 2984
rect 1952 2932 2004 2984
rect 2964 2932 3016 2984
rect 3240 2975 3292 2984
rect 1676 2864 1728 2916
rect 3240 2941 3249 2975
rect 3249 2941 3283 2975
rect 3283 2941 3292 2975
rect 3240 2932 3292 2941
rect 3332 2932 3384 2984
rect 3516 2975 3568 2984
rect 3516 2941 3525 2975
rect 3525 2941 3559 2975
rect 3559 2941 3568 2975
rect 3516 2932 3568 2941
rect 4160 3068 4212 3120
rect 4436 3068 4488 3120
rect 6644 3111 6696 3120
rect 6644 3077 6653 3111
rect 6653 3077 6687 3111
rect 6687 3077 6696 3111
rect 6644 3068 6696 3077
rect 9680 3068 9732 3120
rect 4252 3000 4304 3052
rect 4436 2975 4488 2984
rect 4436 2941 4445 2975
rect 4445 2941 4479 2975
rect 4479 2941 4488 2975
rect 4436 2932 4488 2941
rect 4528 2975 4580 2984
rect 4528 2941 4537 2975
rect 4537 2941 4571 2975
rect 4571 2941 4580 2975
rect 4528 2932 4580 2941
rect 5172 2975 5224 2984
rect 5172 2941 5181 2975
rect 5181 2941 5215 2975
rect 5215 2941 5224 2975
rect 5172 2932 5224 2941
rect 5632 2932 5684 2984
rect 6184 3000 6236 3052
rect 6920 3000 6972 3052
rect 7656 3000 7708 3052
rect 11060 3043 11112 3052
rect 11060 3009 11069 3043
rect 11069 3009 11103 3043
rect 11103 3009 11112 3043
rect 11060 3000 11112 3009
rect 12440 3000 12492 3052
rect 15568 3000 15620 3052
rect 6552 2975 6604 2984
rect 6552 2941 6561 2975
rect 6561 2941 6595 2975
rect 6595 2941 6604 2975
rect 6552 2932 6604 2941
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 6828 2932 6880 2941
rect 11888 2932 11940 2984
rect 7656 2907 7708 2916
rect 2412 2839 2464 2848
rect 2412 2805 2421 2839
rect 2421 2805 2455 2839
rect 2455 2805 2464 2839
rect 2412 2796 2464 2805
rect 3516 2796 3568 2848
rect 3976 2796 4028 2848
rect 4896 2796 4948 2848
rect 7656 2873 7665 2907
rect 7665 2873 7699 2907
rect 7699 2873 7708 2907
rect 7656 2864 7708 2873
rect 8668 2864 8720 2916
rect 9772 2864 9824 2916
rect 11704 2864 11756 2916
rect 13820 2864 13872 2916
rect 7380 2796 7432 2848
rect 13728 2796 13780 2848
rect 5980 2694 6032 2746
rect 6044 2694 6096 2746
rect 6108 2694 6160 2746
rect 6172 2694 6224 2746
rect 10979 2694 11031 2746
rect 11043 2694 11095 2746
rect 11107 2694 11159 2746
rect 11171 2694 11223 2746
rect 2964 2592 3016 2644
rect 3976 2592 4028 2644
rect 5632 2635 5684 2644
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 1676 2567 1728 2576
rect 1676 2533 1685 2567
rect 1685 2533 1719 2567
rect 1719 2533 1728 2567
rect 1676 2524 1728 2533
rect 2412 2524 2464 2576
rect 4160 2567 4212 2576
rect 4160 2533 4169 2567
rect 4169 2533 4203 2567
rect 4203 2533 4212 2567
rect 4160 2524 4212 2533
rect 4896 2524 4948 2576
rect 6828 2592 6880 2644
rect 7656 2592 7708 2644
rect 8668 2592 8720 2644
rect 11520 2592 11572 2644
rect 12164 2635 12216 2644
rect 12164 2601 12173 2635
rect 12173 2601 12207 2635
rect 12207 2601 12216 2635
rect 12164 2592 12216 2601
rect 13820 2592 13872 2644
rect 15568 2635 15620 2644
rect 15568 2601 15577 2635
rect 15577 2601 15611 2635
rect 15611 2601 15620 2635
rect 15568 2592 15620 2601
rect 7012 2524 7064 2576
rect 7196 2524 7248 2576
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 6460 2456 6512 2508
rect 10048 2456 10100 2508
rect 11980 2499 12032 2508
rect 11980 2465 11989 2499
rect 11989 2465 12023 2499
rect 12023 2465 12032 2499
rect 11980 2456 12032 2465
rect 12440 2456 12492 2508
rect 13728 2499 13780 2508
rect 13728 2465 13737 2499
rect 13737 2465 13771 2499
rect 13771 2465 13780 2499
rect 13728 2456 13780 2465
rect 15752 2499 15804 2508
rect 15752 2465 15761 2499
rect 15761 2465 15795 2499
rect 15795 2465 15804 2499
rect 15752 2456 15804 2465
rect 6000 2363 6052 2372
rect 6000 2329 6009 2363
rect 6009 2329 6043 2363
rect 6043 2329 6052 2363
rect 6000 2320 6052 2329
rect 3481 2150 3533 2202
rect 3545 2150 3597 2202
rect 3609 2150 3661 2202
rect 3673 2150 3725 2202
rect 8480 2150 8532 2202
rect 8544 2150 8596 2202
rect 8608 2150 8660 2202
rect 8672 2150 8724 2202
rect 13478 2150 13530 2202
rect 13542 2150 13594 2202
rect 13606 2150 13658 2202
rect 13670 2150 13722 2202
<< metal2 >>
rect 5078 18590 5134 19390
rect 11058 18590 11114 19390
rect 16578 18590 16634 19390
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 1412 16658 1440 17711
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1952 14476 2004 14482
rect 1952 14418 2004 14424
rect 1492 13728 1544 13734
rect 1492 13670 1544 13676
rect 1504 13326 1532 13670
rect 1492 13320 1544 13326
rect 1492 13262 1544 13268
rect 1964 12782 1992 14418
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2240 13802 2268 14214
rect 2228 13796 2280 13802
rect 2228 13738 2280 13744
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1688 11150 1716 12174
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1412 8945 1440 9454
rect 1688 8974 1716 11086
rect 1964 10606 1992 12718
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2240 12374 2268 12582
rect 2228 12368 2280 12374
rect 2228 12310 2280 12316
rect 2136 11280 2188 11286
rect 2136 11222 2188 11228
rect 2148 10810 2176 11222
rect 2228 11008 2280 11014
rect 2228 10950 2280 10956
rect 2240 10810 2268 10950
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1964 9994 1992 10542
rect 1952 9988 2004 9994
rect 1952 9930 2004 9936
rect 1964 9518 1992 9930
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1676 8968 1728 8974
rect 1398 8936 1454 8945
rect 1676 8910 1728 8916
rect 1398 8871 1454 8880
rect 1688 5710 1716 8910
rect 1964 6254 1992 9454
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2240 9110 2268 9318
rect 2228 9104 2280 9110
rect 2228 9046 2280 9052
rect 2332 8922 2360 16730
rect 3455 16348 3751 16368
rect 3511 16346 3535 16348
rect 3591 16346 3615 16348
rect 3671 16346 3695 16348
rect 3533 16294 3535 16346
rect 3597 16294 3609 16346
rect 3671 16294 3673 16346
rect 3511 16292 3535 16294
rect 3591 16292 3615 16294
rect 3671 16292 3695 16294
rect 3455 16272 3751 16292
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 3424 16176 3476 16182
rect 3424 16118 3476 16124
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3160 15994 3188 16050
rect 2412 15972 2464 15978
rect 3160 15966 3280 15994
rect 2412 15914 2464 15920
rect 2424 15706 2452 15914
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2884 13734 2912 15438
rect 3252 15366 3280 15966
rect 3436 15570 3464 16118
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 3528 15706 3556 15982
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 3804 15570 3832 16186
rect 4436 16176 4488 16182
rect 4436 16118 4488 16124
rect 4252 15972 4304 15978
rect 4252 15914 4304 15920
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 3792 15564 3844 15570
rect 3792 15506 3844 15512
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3252 13870 3280 15302
rect 3455 15260 3751 15280
rect 3511 15258 3535 15260
rect 3591 15258 3615 15260
rect 3671 15258 3695 15260
rect 3533 15206 3535 15258
rect 3597 15206 3609 15258
rect 3671 15206 3673 15258
rect 3511 15204 3535 15206
rect 3591 15204 3615 15206
rect 3671 15204 3695 15206
rect 3455 15184 3751 15204
rect 3804 14550 3832 15506
rect 4172 14890 4200 15642
rect 4264 15570 4292 15914
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4344 15564 4396 15570
rect 4344 15506 4396 15512
rect 4252 15428 4304 15434
rect 4252 15370 4304 15376
rect 4160 14884 4212 14890
rect 4160 14826 4212 14832
rect 3792 14544 3844 14550
rect 3792 14486 3844 14492
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3344 13938 3372 14214
rect 3455 14172 3751 14192
rect 3511 14170 3535 14172
rect 3591 14170 3615 14172
rect 3671 14170 3695 14172
rect 3533 14118 3535 14170
rect 3597 14118 3609 14170
rect 3671 14118 3673 14170
rect 3511 14116 3535 14118
rect 3591 14116 3615 14118
rect 3671 14116 3695 14118
rect 3455 14096 3751 14116
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3804 13870 3832 14214
rect 3896 14006 3924 14214
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 2872 13728 2924 13734
rect 2872 13670 2924 13676
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 2884 12238 2912 12310
rect 3252 12306 3280 13806
rect 3988 13734 4016 14418
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 4080 14006 4108 14282
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 4172 13938 4200 14826
rect 4264 14346 4292 15370
rect 4356 15162 4384 15506
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4448 14634 4476 16118
rect 4356 14606 4476 14634
rect 4356 14414 4384 14606
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4252 14340 4304 14346
rect 4252 14282 4304 14288
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4068 13864 4120 13870
rect 4264 13818 4292 14282
rect 4120 13812 4292 13818
rect 4068 13806 4292 13812
rect 4080 13790 4292 13806
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3455 13084 3751 13104
rect 3511 13082 3535 13084
rect 3591 13082 3615 13084
rect 3671 13082 3695 13084
rect 3533 13030 3535 13082
rect 3597 13030 3609 13082
rect 3671 13030 3673 13082
rect 3511 13028 3535 13030
rect 3591 13028 3615 13030
rect 3671 13028 3695 13030
rect 3455 13008 3751 13028
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3528 12306 3556 12718
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3896 12442 3924 12650
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3896 12306 3924 12378
rect 3240 12300 3292 12306
rect 3240 12242 3292 12248
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 3455 11996 3751 12016
rect 3511 11994 3535 11996
rect 3591 11994 3615 11996
rect 3671 11994 3695 11996
rect 3533 11942 3535 11994
rect 3597 11942 3609 11994
rect 3671 11942 3673 11994
rect 3511 11940 3535 11942
rect 3591 11940 3615 11942
rect 3671 11940 3695 11942
rect 3455 11920 3751 11940
rect 4080 11830 4108 13790
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4172 12374 4200 12582
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 4252 12368 4304 12374
rect 4356 12356 4384 14350
rect 4448 13326 4476 14486
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4304 12328 4384 12356
rect 4252 12310 4304 12316
rect 2780 11824 2832 11830
rect 2780 11766 2832 11772
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 2792 10538 2820 11766
rect 4264 11200 4292 12310
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4356 11694 4384 12038
rect 4448 11830 4476 12038
rect 4436 11824 4488 11830
rect 4436 11766 4488 11772
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4172 11172 4292 11200
rect 4436 11212 4488 11218
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 3455 10908 3751 10928
rect 3511 10906 3535 10908
rect 3591 10906 3615 10908
rect 3671 10906 3695 10908
rect 3533 10854 3535 10906
rect 3597 10854 3609 10906
rect 3671 10854 3673 10906
rect 3511 10852 3535 10854
rect 3591 10852 3615 10854
rect 3671 10852 3695 10854
rect 3455 10832 3751 10852
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2780 10532 2832 10538
rect 2780 10474 2832 10480
rect 2792 9518 2820 10474
rect 2976 9722 3004 10746
rect 3804 10742 3832 11018
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 3804 10606 3832 10678
rect 3896 10606 3924 11086
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4080 10606 4108 10950
rect 4172 10810 4200 11172
rect 4436 11154 4488 11160
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3240 10600 3292 10606
rect 3424 10600 3476 10606
rect 3292 10560 3424 10588
rect 3240 10542 3292 10548
rect 3424 10542 3476 10548
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 3068 10266 3096 10542
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 3252 9654 3280 10542
rect 3896 10062 3924 10542
rect 4080 10130 4108 10542
rect 4172 10198 4200 10746
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 4356 10130 4384 11018
rect 4448 10606 4476 11154
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4448 10266 4476 10542
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3455 9820 3751 9840
rect 3511 9818 3535 9820
rect 3591 9818 3615 9820
rect 3671 9818 3695 9820
rect 3533 9766 3535 9818
rect 3597 9766 3609 9818
rect 3671 9766 3673 9818
rect 3511 9764 3535 9766
rect 3591 9764 3615 9766
rect 3671 9764 3695 9766
rect 3455 9744 3751 9764
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2516 9178 2544 9318
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2240 8894 2360 8922
rect 2240 8430 2268 8894
rect 3344 8838 3372 9454
rect 4080 9042 4108 10066
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 3455 8732 3751 8752
rect 3511 8730 3535 8732
rect 3591 8730 3615 8732
rect 3671 8730 3695 8732
rect 3533 8678 3535 8730
rect 3597 8678 3609 8730
rect 3671 8678 3673 8730
rect 3511 8676 3535 8678
rect 3591 8676 3615 8678
rect 3671 8676 3695 8678
rect 3455 8656 3751 8676
rect 4172 8498 4200 8774
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 2044 8016 2096 8022
rect 2044 7958 2096 7964
rect 2056 7410 2084 7958
rect 2240 7886 2268 8366
rect 2332 7954 2360 8366
rect 4264 8022 4292 8366
rect 4356 8294 4384 8502
rect 4448 8430 4476 8978
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 4356 7954 4384 8230
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2332 7546 2360 7890
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2608 7274 2636 7822
rect 2700 7410 2728 7890
rect 3160 7478 3188 7890
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 2596 7268 2648 7274
rect 2596 7210 2648 7216
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 2504 6248 2556 6254
rect 2504 6190 2556 6196
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1872 5846 1900 6054
rect 1860 5840 1912 5846
rect 1860 5782 1912 5788
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1688 4146 1716 5646
rect 1964 4690 1992 6190
rect 2516 4758 2544 6190
rect 2608 4826 2636 7210
rect 3068 6322 3096 7210
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 2780 6180 2832 6186
rect 2780 6122 2832 6128
rect 2792 5914 2820 6122
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2884 5846 2912 6054
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2504 4752 2556 4758
rect 2504 4694 2556 4700
rect 3068 4690 3096 6258
rect 3160 6186 3188 7278
rect 3344 7206 3372 7890
rect 4448 7818 4476 8366
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 3455 7644 3751 7664
rect 3511 7642 3535 7644
rect 3591 7642 3615 7644
rect 3671 7642 3695 7644
rect 3533 7590 3535 7642
rect 3597 7590 3609 7642
rect 3671 7590 3673 7642
rect 3511 7588 3535 7590
rect 3591 7588 3615 7590
rect 3671 7588 3695 7590
rect 3455 7568 3751 7588
rect 4540 7342 4568 16730
rect 5092 16658 5120 18590
rect 11072 17626 11100 18590
rect 11072 17598 11376 17626
rect 5954 16892 6250 16912
rect 6010 16890 6034 16892
rect 6090 16890 6114 16892
rect 6170 16890 6194 16892
rect 6032 16838 6034 16890
rect 6096 16838 6108 16890
rect 6170 16838 6172 16890
rect 6010 16836 6034 16838
rect 6090 16836 6114 16838
rect 6170 16836 6194 16838
rect 5954 16816 6250 16836
rect 10953 16892 11249 16912
rect 11009 16890 11033 16892
rect 11089 16890 11113 16892
rect 11169 16890 11193 16892
rect 11031 16838 11033 16890
rect 11095 16838 11107 16890
rect 11169 16838 11171 16890
rect 11009 16836 11033 16838
rect 11089 16836 11113 16838
rect 11169 16836 11193 16838
rect 10953 16816 11249 16836
rect 11348 16794 11376 17598
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 16592 16726 16620 18590
rect 6736 16720 6788 16726
rect 6736 16662 6788 16668
rect 16580 16720 16632 16726
rect 16580 16662 16632 16668
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4632 14958 4660 15846
rect 4724 15706 4752 16050
rect 5080 16040 5132 16046
rect 5000 15988 5080 15994
rect 5000 15982 5132 15988
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5000 15966 5120 15982
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4724 15366 4752 15506
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 5000 15162 5028 15966
rect 5080 15904 5132 15910
rect 5080 15846 5132 15852
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5092 15638 5120 15846
rect 5184 15706 5212 15846
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5080 15632 5132 15638
rect 5080 15574 5132 15580
rect 5264 15360 5316 15366
rect 5368 15314 5396 15982
rect 6564 15910 6592 16050
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 5828 15638 5856 15846
rect 5954 15804 6250 15824
rect 6010 15802 6034 15804
rect 6090 15802 6114 15804
rect 6170 15802 6194 15804
rect 6032 15750 6034 15802
rect 6096 15750 6108 15802
rect 6170 15750 6172 15802
rect 6010 15748 6034 15750
rect 6090 15748 6114 15750
rect 6170 15748 6194 15750
rect 5954 15728 6250 15748
rect 5816 15632 5868 15638
rect 5816 15574 5868 15580
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 5316 15308 5396 15314
rect 5264 15302 5396 15308
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5276 15286 5396 15302
rect 4988 15156 5040 15162
rect 4988 15098 5040 15104
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4632 13870 4660 14894
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 4908 13870 4936 14350
rect 5000 14006 5028 15098
rect 5368 14618 5396 15286
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 4988 14000 5040 14006
rect 4988 13942 5040 13948
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 4724 13394 4752 13806
rect 4908 13530 4936 13806
rect 5000 13734 5028 13942
rect 5368 13870 5396 14350
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5552 13938 5580 14282
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 5368 13394 5396 13806
rect 5552 13394 5580 13874
rect 5644 13530 5672 14214
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4632 10810 4660 12242
rect 4724 12102 4752 13330
rect 5172 12708 5224 12714
rect 5172 12650 5224 12656
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 5000 12306 5028 12378
rect 5184 12306 5212 12650
rect 5368 12442 5396 13330
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4724 11150 4752 12038
rect 5092 11218 5120 12174
rect 5460 12170 5488 12718
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 5552 11914 5580 13330
rect 5736 13326 5764 14418
rect 5828 13938 5856 15302
rect 6472 14890 6500 15506
rect 6460 14884 6512 14890
rect 6460 14826 6512 14832
rect 5954 14716 6250 14736
rect 6010 14714 6034 14716
rect 6090 14714 6114 14716
rect 6170 14714 6194 14716
rect 6032 14662 6034 14714
rect 6096 14662 6108 14714
rect 6170 14662 6172 14714
rect 6010 14660 6034 14662
rect 6090 14660 6114 14662
rect 6170 14660 6194 14662
rect 5954 14640 6250 14660
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 5828 13530 5856 13874
rect 6564 13870 6592 15846
rect 6656 15366 6684 15982
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 5954 13628 6250 13648
rect 6010 13626 6034 13628
rect 6090 13626 6114 13628
rect 6170 13626 6194 13628
rect 6032 13574 6034 13626
rect 6096 13574 6108 13626
rect 6170 13574 6172 13626
rect 6010 13572 6034 13574
rect 6090 13572 6114 13574
rect 6170 13572 6194 13574
rect 5954 13552 6250 13572
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 6288 13258 6316 13330
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6276 13252 6328 13258
rect 6276 13194 6328 13200
rect 6564 12782 6592 13262
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6276 12708 6328 12714
rect 6276 12650 6328 12656
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5736 12306 5764 12582
rect 5954 12540 6250 12560
rect 6010 12538 6034 12540
rect 6090 12538 6114 12540
rect 6170 12538 6194 12540
rect 6032 12486 6034 12538
rect 6096 12486 6108 12538
rect 6170 12486 6172 12538
rect 6010 12484 6034 12486
rect 6090 12484 6114 12486
rect 6170 12484 6194 12486
rect 5954 12464 6250 12484
rect 6092 12368 6144 12374
rect 6144 12328 6224 12356
rect 6092 12310 6144 12316
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5828 11914 5856 12174
rect 5552 11886 5856 11914
rect 6012 11694 6040 12242
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 5368 11354 5396 11630
rect 5448 11552 5500 11558
rect 6196 11540 6224 12328
rect 6288 12170 6316 12650
rect 6564 12306 6592 12718
rect 6748 12434 6776 16662
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 8454 16348 8750 16368
rect 8510 16346 8534 16348
rect 8590 16346 8614 16348
rect 8670 16346 8694 16348
rect 8532 16294 8534 16346
rect 8596 16294 8608 16346
rect 8670 16294 8672 16346
rect 8510 16292 8534 16294
rect 8590 16292 8614 16294
rect 8670 16292 8694 16294
rect 8454 16272 8750 16292
rect 11256 16250 11284 16594
rect 13452 16348 13748 16368
rect 13508 16346 13532 16348
rect 13588 16346 13612 16348
rect 13668 16346 13692 16348
rect 13530 16294 13532 16346
rect 13594 16294 13606 16346
rect 13668 16294 13670 16346
rect 13508 16292 13532 16294
rect 13588 16292 13612 16294
rect 13668 16292 13692 16294
rect 13452 16272 13748 16292
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 9864 16040 9916 16046
rect 9864 15982 9916 15988
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 7024 15706 7052 15982
rect 9220 15972 9272 15978
rect 9220 15914 9272 15920
rect 9232 15706 9260 15914
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 7024 14074 7052 15506
rect 8454 15260 8750 15280
rect 8510 15258 8534 15260
rect 8590 15258 8614 15260
rect 8670 15258 8694 15260
rect 8532 15206 8534 15258
rect 8596 15206 8608 15258
rect 8670 15206 8672 15258
rect 8510 15204 8534 15206
rect 8590 15204 8614 15206
rect 8670 15204 8694 15206
rect 8454 15184 8750 15204
rect 9600 15162 9628 15506
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 6656 12406 6776 12434
rect 6920 12436 6972 12442
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6276 12164 6328 12170
rect 6276 12106 6328 12112
rect 6472 11898 6500 12242
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6276 11552 6328 11558
rect 6196 11512 6276 11540
rect 5448 11494 5500 11500
rect 6276 11494 6328 11500
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5080 11212 5132 11218
rect 5000 11172 5080 11200
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4632 10674 4660 10746
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4632 8838 4660 10610
rect 4724 10130 4752 10950
rect 5000 10810 5028 11172
rect 5080 11154 5132 11160
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 5092 10606 5120 10950
rect 5460 10606 5488 11494
rect 5954 11452 6250 11472
rect 6010 11450 6034 11452
rect 6090 11450 6114 11452
rect 6170 11450 6194 11452
rect 6032 11398 6034 11450
rect 6096 11398 6108 11450
rect 6170 11398 6172 11450
rect 6010 11396 6034 11398
rect 6090 11396 6114 11398
rect 6170 11396 6194 11398
rect 5954 11376 6250 11396
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5276 10198 5304 10542
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5828 10266 5856 10406
rect 5954 10364 6250 10384
rect 6010 10362 6034 10364
rect 6090 10362 6114 10364
rect 6170 10362 6194 10364
rect 6032 10310 6034 10362
rect 6096 10310 6108 10362
rect 6170 10310 6172 10362
rect 6010 10308 6034 10310
rect 6090 10308 6114 10310
rect 6170 10308 6194 10310
rect 5954 10288 6250 10308
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 5828 10130 5856 10202
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4632 8362 4660 8774
rect 4724 8634 4752 8978
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4816 8566 4844 10066
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6380 9586 6408 9862
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 4804 8560 4856 8566
rect 4804 8502 4856 8508
rect 5276 8430 5304 8774
rect 5368 8566 5396 8978
rect 5736 8974 5764 9454
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 5828 9110 5856 9386
rect 5954 9276 6250 9296
rect 6010 9274 6034 9276
rect 6090 9274 6114 9276
rect 6170 9274 6194 9276
rect 6032 9222 6034 9274
rect 6096 9222 6108 9274
rect 6170 9222 6172 9274
rect 6010 9220 6034 9222
rect 6090 9220 6114 9222
rect 6170 9220 6194 9222
rect 5954 9200 6250 9220
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3344 7002 3372 7142
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3884 6724 3936 6730
rect 3884 6666 3936 6672
rect 3455 6556 3751 6576
rect 3511 6554 3535 6556
rect 3591 6554 3615 6556
rect 3671 6554 3695 6556
rect 3533 6502 3535 6554
rect 3597 6502 3609 6554
rect 3671 6502 3673 6554
rect 3511 6500 3535 6502
rect 3591 6500 3615 6502
rect 3671 6500 3695 6502
rect 3455 6480 3751 6500
rect 3896 6254 3924 6666
rect 3988 6254 4016 6938
rect 5092 6934 5120 7890
rect 5080 6928 5132 6934
rect 5080 6870 5132 6876
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 4528 6792 4580 6798
rect 4816 6746 4844 6802
rect 4580 6740 4844 6746
rect 4528 6734 4844 6740
rect 4540 6718 4844 6734
rect 4540 6458 4568 6718
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 5000 6338 5028 6802
rect 5092 6458 5120 6870
rect 5184 6730 5212 8366
rect 5368 8022 5396 8502
rect 5828 8498 5856 8774
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 6104 8430 6132 8774
rect 6656 8566 6684 12406
rect 6920 12378 6972 12384
rect 6932 12238 6960 12378
rect 7024 12306 7052 13806
rect 7208 13190 7236 13806
rect 7196 13184 7248 13190
rect 7248 13144 7328 13172
rect 7196 13126 7248 13132
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6748 11218 6776 11562
rect 6932 11286 6960 12174
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 7024 11014 7052 12242
rect 7116 11801 7144 12718
rect 7300 12714 7328 13144
rect 7196 12708 7248 12714
rect 7196 12650 7248 12656
rect 7288 12708 7340 12714
rect 7288 12650 7340 12656
rect 7102 11792 7158 11801
rect 7102 11727 7158 11736
rect 7116 11218 7144 11727
rect 7208 11354 7236 12650
rect 7576 11354 7604 14350
rect 7668 13326 7696 14894
rect 8220 14482 8248 14894
rect 8852 14884 8904 14890
rect 8852 14826 8904 14832
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8454 14172 8750 14192
rect 8510 14170 8534 14172
rect 8590 14170 8614 14172
rect 8670 14170 8694 14172
rect 8532 14118 8534 14170
rect 8596 14118 8608 14170
rect 8670 14118 8672 14170
rect 8510 14116 8534 14118
rect 8590 14116 8614 14118
rect 8670 14116 8694 14118
rect 8454 14096 8750 14116
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7668 12986 7696 13262
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7668 12374 7696 12786
rect 7760 12646 7788 13466
rect 8864 13394 8892 14826
rect 9048 14074 9076 14894
rect 9140 14618 9168 14894
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9232 13841 9260 13874
rect 9218 13832 9274 13841
rect 9218 13767 9274 13776
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7944 12918 7972 13262
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 7932 12912 7984 12918
rect 7932 12854 7984 12860
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 7116 10742 7144 11154
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 7760 10198 7788 12582
rect 7852 11218 7880 12718
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 7944 12170 7972 12650
rect 8036 12306 8064 12922
rect 8312 12866 8340 13330
rect 8454 13084 8750 13104
rect 8510 13082 8534 13084
rect 8590 13082 8614 13084
rect 8670 13082 8694 13084
rect 8532 13030 8534 13082
rect 8596 13030 8608 13082
rect 8670 13030 8672 13082
rect 8510 13028 8534 13030
rect 8590 13028 8614 13030
rect 8670 13028 8694 13030
rect 8454 13008 8750 13028
rect 8484 12912 8536 12918
rect 8312 12838 8432 12866
rect 8484 12854 8536 12860
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8312 12374 8340 12650
rect 8404 12442 8432 12838
rect 8496 12782 8524 12854
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8116 12368 8168 12374
rect 8116 12310 8168 12316
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8128 12209 8156 12310
rect 8496 12306 8524 12718
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8114 12200 8170 12209
rect 7932 12164 7984 12170
rect 8114 12135 8170 12144
rect 7932 12106 7984 12112
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8312 11898 8340 12038
rect 8454 11996 8750 12016
rect 8510 11994 8534 11996
rect 8590 11994 8614 11996
rect 8670 11994 8694 11996
rect 8532 11942 8534 11994
rect 8596 11942 8608 11994
rect 8670 11942 8672 11994
rect 8510 11940 8534 11942
rect 8590 11940 8614 11942
rect 8670 11940 8694 11942
rect 8454 11920 8750 11940
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8760 11688 8812 11694
rect 8864 11676 8892 13330
rect 9048 12306 9076 13330
rect 9324 13326 9352 13874
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9324 12986 9352 13262
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9324 12306 9352 12922
rect 9416 12850 9444 14010
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9496 13864 9548 13870
rect 9548 13824 9720 13852
rect 9496 13806 9548 13812
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 9312 12300 9364 12306
rect 9416 12288 9444 12786
rect 9588 12300 9640 12306
rect 9416 12260 9588 12288
rect 9312 12242 9364 12248
rect 9588 12242 9640 12248
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8956 11830 8984 12038
rect 8944 11824 8996 11830
rect 8944 11766 8996 11772
rect 8812 11648 8892 11676
rect 8760 11630 8812 11636
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8128 11354 8156 11494
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7852 10606 7880 11154
rect 8128 10810 8156 11290
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 7840 10600 7892 10606
rect 8312 10588 8340 11494
rect 8864 11218 8892 11648
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 8864 11082 8892 11154
rect 8956 11150 8984 11630
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 8454 10908 8750 10928
rect 8510 10906 8534 10908
rect 8590 10906 8614 10908
rect 8670 10906 8694 10908
rect 8532 10854 8534 10906
rect 8596 10854 8608 10906
rect 8670 10854 8672 10906
rect 8510 10852 8534 10854
rect 8590 10852 8614 10854
rect 8670 10852 8694 10854
rect 8454 10832 8750 10852
rect 8392 10600 8444 10606
rect 8312 10560 8392 10588
rect 7840 10542 7892 10548
rect 8392 10542 8444 10548
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7852 9994 7880 10542
rect 8864 10538 8892 11018
rect 8852 10532 8904 10538
rect 8852 10474 8904 10480
rect 7840 9988 7892 9994
rect 7840 9930 7892 9936
rect 8852 9988 8904 9994
rect 8852 9930 8904 9936
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7024 9450 7052 9862
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 6656 8430 6684 8502
rect 6840 8498 6868 8978
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 5460 8294 5488 8366
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5954 8188 6250 8208
rect 6010 8186 6034 8188
rect 6090 8186 6114 8188
rect 6170 8186 6194 8188
rect 6032 8134 6034 8186
rect 6096 8134 6108 8186
rect 6170 8134 6172 8186
rect 6010 8132 6034 8134
rect 6090 8132 6114 8134
rect 6170 8132 6194 8134
rect 5954 8112 6250 8132
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5000 6310 5120 6338
rect 5092 6254 5120 6310
rect 5460 6254 5488 7278
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 3252 5370 3280 5782
rect 3792 5772 3844 5778
rect 3792 5714 3844 5720
rect 3455 5468 3751 5488
rect 3511 5466 3535 5468
rect 3591 5466 3615 5468
rect 3671 5466 3695 5468
rect 3533 5414 3535 5466
rect 3597 5414 3609 5466
rect 3671 5414 3673 5466
rect 3511 5412 3535 5414
rect 3591 5412 3615 5414
rect 3671 5412 3695 5414
rect 3455 5392 3751 5412
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3804 4758 3832 5714
rect 3896 5658 3924 6190
rect 3988 5846 4016 6190
rect 4252 6180 4304 6186
rect 4252 6122 4304 6128
rect 3976 5840 4028 5846
rect 3976 5782 4028 5788
rect 4264 5778 4292 6122
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 3976 5704 4028 5710
rect 3896 5652 3976 5658
rect 3896 5646 4028 5652
rect 3896 5630 4016 5646
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 480 2984 532 2990
rect 480 2926 532 2932
rect 492 800 520 2926
rect 1412 2514 1440 4082
rect 1964 2990 1992 4626
rect 2228 4480 2280 4486
rect 2228 4422 2280 4428
rect 2412 4480 2464 4486
rect 2412 4422 2464 4428
rect 2240 4010 2268 4422
rect 2424 4282 2452 4422
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2228 4004 2280 4010
rect 2228 3946 2280 3952
rect 2792 3058 2820 4626
rect 3068 4282 3096 4626
rect 3455 4380 3751 4400
rect 3511 4378 3535 4380
rect 3591 4378 3615 4380
rect 3671 4378 3695 4380
rect 3533 4326 3535 4378
rect 3597 4326 3609 4378
rect 3671 4326 3673 4378
rect 3511 4324 3535 4326
rect 3591 4324 3615 4326
rect 3671 4324 3695 4326
rect 3455 4304 3751 4324
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3252 3738 3280 4218
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3252 3126 3280 3674
rect 3988 3670 4016 5630
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4172 4826 4200 5034
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 3252 2990 3280 3062
rect 3344 2990 3372 3538
rect 3455 3292 3751 3312
rect 3511 3290 3535 3292
rect 3591 3290 3615 3292
rect 3671 3290 3695 3292
rect 3533 3238 3535 3290
rect 3597 3238 3609 3290
rect 3671 3238 3673 3290
rect 3511 3236 3535 3238
rect 3591 3236 3615 3238
rect 3671 3236 3695 3238
rect 3455 3216 3751 3236
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 1676 2916 1728 2922
rect 1676 2858 1728 2864
rect 1688 2582 1716 2858
rect 2412 2848 2464 2854
rect 2412 2790 2464 2796
rect 2424 2582 2452 2790
rect 2976 2650 3004 2926
rect 3528 2854 3556 2926
rect 3988 2854 4016 3606
rect 4264 3602 4292 5714
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4724 5234 4752 5510
rect 5000 5234 5028 5578
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 5000 4758 5028 5170
rect 4528 4752 4580 4758
rect 4528 4694 4580 4700
rect 4988 4752 5040 4758
rect 4988 4694 5040 4700
rect 4540 4486 4568 4694
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 3988 2650 4016 2790
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 4172 2582 4200 3062
rect 4264 3058 4292 3402
rect 4436 3120 4488 3126
rect 4436 3062 4488 3068
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4448 2990 4476 3062
rect 4540 2990 4568 4422
rect 5092 3194 5120 6190
rect 5552 6186 5580 6802
rect 5644 6390 5672 7890
rect 5828 7546 5856 7890
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5954 7100 6250 7120
rect 6010 7098 6034 7100
rect 6090 7098 6114 7100
rect 6170 7098 6194 7100
rect 6032 7046 6034 7098
rect 6096 7046 6108 7098
rect 6170 7046 6172 7098
rect 6010 7044 6034 7046
rect 6090 7044 6114 7046
rect 6170 7044 6194 7046
rect 5954 7024 6250 7044
rect 6564 7002 6592 8366
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6196 6458 6224 6802
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 5632 6384 5684 6390
rect 5632 6326 5684 6332
rect 5736 6254 5764 6394
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 5184 4622 5212 5238
rect 5552 5030 5580 6122
rect 5632 5840 5684 5846
rect 5632 5782 5684 5788
rect 5644 5098 5672 5782
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5644 4690 5672 5034
rect 5828 4826 5856 6326
rect 5954 6012 6250 6032
rect 6010 6010 6034 6012
rect 6090 6010 6114 6012
rect 6170 6010 6194 6012
rect 6032 5958 6034 6010
rect 6096 5958 6108 6010
rect 6170 5958 6172 6010
rect 6010 5956 6034 5958
rect 6090 5956 6114 5958
rect 6170 5956 6194 5958
rect 5954 5936 6250 5956
rect 6748 5914 6776 6734
rect 6840 6730 6868 8434
rect 6932 8430 6960 9046
rect 7300 8498 7328 9862
rect 7852 9722 7880 9930
rect 8454 9820 8750 9840
rect 8510 9818 8534 9820
rect 8590 9818 8614 9820
rect 8670 9818 8694 9820
rect 8532 9766 8534 9818
rect 8596 9766 8608 9818
rect 8670 9766 8672 9818
rect 8510 9764 8534 9766
rect 8590 9764 8614 9766
rect 8670 9764 8694 9766
rect 8454 9744 8750 9764
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 8864 9450 8892 9930
rect 9048 9518 9076 12242
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9232 11778 9260 12174
rect 9312 12164 9364 12170
rect 9496 12164 9548 12170
rect 9312 12106 9364 12112
rect 9416 12124 9496 12152
rect 9140 11750 9260 11778
rect 9140 11694 9168 11750
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9324 11558 9352 12106
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8128 9178 8156 9386
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 7300 7954 7328 8434
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 8022 7788 8230
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 8128 7886 8156 9114
rect 9140 9042 9168 11018
rect 9324 11014 9352 11494
rect 9416 11354 9444 12124
rect 9496 12106 9548 12112
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9600 11801 9628 11834
rect 9586 11792 9642 11801
rect 9586 11727 9642 11736
rect 9692 11694 9720 13824
rect 9784 13530 9812 13942
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9784 12986 9812 13466
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9784 12442 9812 12718
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9784 12238 9812 12378
rect 9876 12374 9904 15982
rect 10953 15804 11249 15824
rect 11009 15802 11033 15804
rect 11089 15802 11113 15804
rect 11169 15802 11193 15804
rect 11031 15750 11033 15802
rect 11095 15750 11107 15802
rect 11169 15750 11171 15802
rect 11009 15748 11033 15750
rect 11089 15748 11113 15750
rect 11169 15748 11193 15750
rect 10953 15728 11249 15748
rect 13280 15638 13308 15982
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 13556 15570 13584 15846
rect 13740 15706 13768 15846
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13832 15570 13860 15846
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 11612 14884 11664 14890
rect 11612 14826 11664 14832
rect 10953 14716 11249 14736
rect 11009 14714 11033 14716
rect 11089 14714 11113 14716
rect 11169 14714 11193 14716
rect 11031 14662 11033 14714
rect 11095 14662 11107 14714
rect 11169 14662 11171 14714
rect 11009 14660 11033 14662
rect 11089 14660 11113 14662
rect 11169 14660 11193 14662
rect 10953 14640 11249 14660
rect 11624 14618 11652 14826
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 9956 13864 10008 13870
rect 9954 13832 9956 13841
rect 10008 13832 10010 13841
rect 9954 13767 10010 13776
rect 10140 13796 10192 13802
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9876 11898 9904 12106
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9600 11558 9628 11630
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9232 10674 9260 10950
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9324 10606 9352 10950
rect 9600 10810 9628 11154
rect 9784 10810 9812 11154
rect 9876 11082 9904 11834
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9876 10742 9904 11018
rect 9864 10736 9916 10742
rect 9864 10678 9916 10684
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9416 10266 9444 10610
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9416 10062 9444 10202
rect 9968 10169 9996 13767
rect 10140 13738 10192 13744
rect 10048 13388 10100 13394
rect 10152 13376 10180 13738
rect 10953 13628 11249 13648
rect 11009 13626 11033 13628
rect 11089 13626 11113 13628
rect 11169 13626 11193 13628
rect 11031 13574 11033 13626
rect 11095 13574 11107 13626
rect 11169 13574 11171 13626
rect 11009 13572 11033 13574
rect 11089 13572 11113 13574
rect 11169 13572 11193 13574
rect 10953 13552 11249 13572
rect 11348 13394 11376 14418
rect 11796 14340 11848 14346
rect 11796 14282 11848 14288
rect 11808 14074 11836 14282
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11716 13530 11744 13670
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 10100 13348 10180 13376
rect 11336 13388 11388 13394
rect 10048 13330 10100 13336
rect 11336 13330 11388 13336
rect 10953 12540 11249 12560
rect 11009 12538 11033 12540
rect 11089 12538 11113 12540
rect 11169 12538 11193 12540
rect 11031 12486 11033 12538
rect 11095 12486 11107 12538
rect 11169 12486 11171 12538
rect 11009 12484 11033 12486
rect 11089 12484 11113 12486
rect 11169 12484 11193 12486
rect 10953 12464 11249 12484
rect 11348 12442 11376 13330
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10230 12200 10286 12209
rect 10230 12135 10232 12144
rect 10284 12135 10286 12144
rect 10232 12106 10284 12112
rect 10244 10266 10272 12106
rect 11072 11898 11100 12242
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 10416 11824 10468 11830
rect 10416 11766 10468 11772
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 9954 10160 10010 10169
rect 9954 10095 9956 10104
rect 10008 10095 10010 10104
rect 9956 10066 10008 10072
rect 9404 10056 9456 10062
rect 9968 10035 9996 10066
rect 9404 9998 9456 10004
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9692 9178 9720 9454
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 8454 8732 8750 8752
rect 8510 8730 8534 8732
rect 8590 8730 8614 8732
rect 8670 8730 8694 8732
rect 8532 8678 8534 8730
rect 8596 8678 8608 8730
rect 8670 8678 8672 8730
rect 8510 8676 8534 8678
rect 8590 8676 8614 8678
rect 8670 8676 8694 8678
rect 8454 8656 8750 8676
rect 9692 8498 9720 9114
rect 9784 8906 9812 9318
rect 10060 9042 10088 9862
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8404 7954 8432 8298
rect 8680 8090 8708 8366
rect 9692 8090 9720 8434
rect 10060 8430 10088 8978
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 8944 8016 8996 8022
rect 8944 7958 8996 7964
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 7342 8156 7822
rect 8454 7644 8750 7664
rect 8510 7642 8534 7644
rect 8590 7642 8614 7644
rect 8670 7642 8694 7644
rect 8532 7590 8534 7642
rect 8596 7590 8608 7642
rect 8670 7590 8672 7642
rect 8510 7588 8534 7590
rect 8590 7588 8614 7590
rect 8670 7588 8694 7590
rect 8454 7568 8750 7588
rect 8864 7342 8892 7890
rect 8956 7546 8984 7958
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9600 6934 9628 7278
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7576 6458 7604 6598
rect 7760 6458 7788 6666
rect 8454 6556 8750 6576
rect 8510 6554 8534 6556
rect 8590 6554 8614 6556
rect 8670 6554 8694 6556
rect 8532 6502 8534 6554
rect 8596 6502 8608 6554
rect 8670 6502 8672 6554
rect 8510 6500 8534 6502
rect 8590 6500 8614 6502
rect 8670 6500 8694 6502
rect 8454 6480 8750 6500
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 7944 6118 7972 6326
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6288 5370 6316 5714
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6288 5030 6316 5306
rect 6472 5166 6500 5646
rect 6748 5234 6776 5714
rect 7944 5710 7972 6054
rect 8128 5846 8156 6190
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 5954 4924 6250 4944
rect 6010 4922 6034 4924
rect 6090 4922 6114 4924
rect 6170 4922 6194 4924
rect 6032 4870 6034 4922
rect 6096 4870 6108 4922
rect 6170 4870 6172 4922
rect 6010 4868 6034 4870
rect 6090 4868 6114 4870
rect 6170 4868 6194 4870
rect 5954 4848 6250 4868
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5184 2990 5212 4558
rect 5368 4078 5396 4558
rect 5460 4214 5488 4626
rect 5448 4208 5500 4214
rect 5448 4150 5500 4156
rect 5644 4146 5672 4626
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 6368 4004 6420 4010
rect 6368 3946 6420 3952
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 5954 3836 6250 3856
rect 6010 3834 6034 3836
rect 6090 3834 6114 3836
rect 6170 3834 6194 3836
rect 6032 3782 6034 3834
rect 6096 3782 6108 3834
rect 6170 3782 6172 3834
rect 6010 3780 6034 3782
rect 6090 3780 6114 3782
rect 6170 3780 6194 3782
rect 5954 3760 6250 3780
rect 6288 3482 6316 3878
rect 6380 3670 6408 3946
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 6472 3602 6500 5102
rect 6748 5030 6776 5170
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6368 3528 6420 3534
rect 6196 3476 6368 3482
rect 6196 3470 6420 3476
rect 6196 3454 6408 3470
rect 6196 3058 6224 3454
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 4436 2984 4488 2990
rect 4436 2926 4488 2932
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 4908 2582 4936 2790
rect 5644 2650 5672 2926
rect 5954 2748 6250 2768
rect 6010 2746 6034 2748
rect 6090 2746 6114 2748
rect 6170 2746 6194 2748
rect 6032 2694 6034 2746
rect 6096 2694 6108 2746
rect 6170 2694 6172 2746
rect 6010 2692 6034 2694
rect 6090 2692 6114 2694
rect 6170 2692 6194 2694
rect 5954 2672 6250 2692
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 1676 2576 1728 2582
rect 1676 2518 1728 2524
rect 2412 2576 2464 2582
rect 2412 2518 2464 2524
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 6472 2514 6500 3538
rect 6564 2990 6592 3878
rect 6656 3534 6684 4014
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6656 3126 6684 3470
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 6840 2990 6868 3538
rect 6932 3058 6960 4626
rect 7024 3738 7052 5578
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7944 4758 7972 4966
rect 7932 4752 7984 4758
rect 7932 4694 7984 4700
rect 8220 4622 8248 5646
rect 8312 5166 8340 5714
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 8454 5468 8750 5488
rect 8510 5466 8534 5468
rect 8590 5466 8614 5468
rect 8670 5466 8694 5468
rect 8532 5414 8534 5466
rect 8596 5414 8608 5466
rect 8670 5414 8672 5466
rect 8510 5412 8534 5414
rect 8590 5412 8614 5414
rect 8670 5412 8694 5414
rect 8454 5392 8750 5412
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 8760 5296 8812 5302
rect 8760 5238 8812 5244
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7024 3602 7052 3674
rect 7208 3618 7236 4558
rect 7300 4078 7328 4558
rect 8312 4486 8340 5102
rect 8772 4554 8800 5238
rect 9048 5166 9076 5306
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 8760 4548 8812 4554
rect 8760 4490 8812 4496
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8454 4380 8750 4400
rect 8510 4378 8534 4380
rect 8590 4378 8614 4380
rect 8670 4378 8694 4380
rect 8532 4326 8534 4378
rect 8596 4326 8608 4378
rect 8670 4326 8672 4378
rect 8510 4324 8534 4326
rect 8590 4324 8614 4326
rect 8670 4324 8694 4326
rect 8454 4304 8750 4324
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7012 3596 7064 3602
rect 7208 3590 7328 3618
rect 9048 3602 9076 5102
rect 9324 5098 9352 5170
rect 9416 5166 9444 5510
rect 9600 5166 9628 6190
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9876 5846 9904 6054
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 10336 5302 10364 8570
rect 10428 7410 10456 11766
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10520 10606 10548 11630
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10520 9722 10548 10542
rect 10612 10130 10640 11698
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10888 11354 10916 11630
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 10953 11452 11249 11472
rect 11009 11450 11033 11452
rect 11089 11450 11113 11452
rect 11169 11450 11193 11452
rect 11031 11398 11033 11450
rect 11095 11398 11107 11450
rect 11169 11398 11171 11450
rect 11009 11396 11033 11398
rect 11089 11396 11113 11398
rect 11169 11396 11193 11398
rect 10953 11376 11249 11396
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10888 10470 10916 11154
rect 11900 10606 11928 11562
rect 12084 10742 12112 13942
rect 12176 13190 12204 14418
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 12176 12306 12204 13126
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12176 11744 12204 12242
rect 12268 12102 12296 13398
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12360 12170 12388 13330
rect 12452 13326 12480 15506
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 13452 15260 13748 15280
rect 13508 15258 13532 15260
rect 13588 15258 13612 15260
rect 13668 15258 13692 15260
rect 13530 15206 13532 15258
rect 13594 15206 13606 15258
rect 13668 15206 13670 15258
rect 13508 15204 13532 15206
rect 13588 15204 13612 15206
rect 13668 15204 13692 15206
rect 13452 15184 13748 15204
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 13004 14006 13032 14418
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 12992 14000 13044 14006
rect 12992 13942 13044 13948
rect 13004 13394 13032 13942
rect 13372 13870 13400 14350
rect 13452 14172 13748 14192
rect 13508 14170 13532 14172
rect 13588 14170 13612 14172
rect 13668 14170 13692 14172
rect 13530 14118 13532 14170
rect 13594 14118 13606 14170
rect 13668 14118 13670 14170
rect 13508 14116 13532 14118
rect 13588 14116 13612 14118
rect 13668 14116 13692 14118
rect 13452 14096 13748 14116
rect 13832 14006 13860 14554
rect 14200 14550 14228 15438
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 14188 14544 14240 14550
rect 14188 14486 14240 14492
rect 13912 14340 13964 14346
rect 13912 14282 13964 14288
rect 13924 14074 13952 14282
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 14844 14006 14872 14214
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 14832 14000 14884 14006
rect 14832 13942 14884 13948
rect 15028 13870 15056 15370
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 13096 13394 13124 13806
rect 13372 13530 13400 13806
rect 14660 13734 14688 13806
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 14660 13462 14688 13670
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12440 12368 12492 12374
rect 12440 12310 12492 12316
rect 12452 12170 12480 12310
rect 12348 12164 12400 12170
rect 12348 12106 12400 12112
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12256 11756 12308 11762
rect 12176 11716 12256 11744
rect 12256 11698 12308 11704
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 12268 10606 12296 11698
rect 12360 11626 12388 12106
rect 12452 11694 12480 12106
rect 12728 12102 12756 13330
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 12820 12986 12848 13194
rect 13452 13084 13748 13104
rect 13508 13082 13532 13084
rect 13588 13082 13612 13084
rect 13668 13082 13692 13084
rect 13530 13030 13532 13082
rect 13594 13030 13606 13082
rect 13668 13030 13670 13082
rect 13508 13028 13532 13030
rect 13588 13028 13612 13030
rect 13668 13028 13692 13030
rect 13452 13008 13748 13028
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12348 11620 12400 11626
rect 12348 11562 12400 11568
rect 12452 10674 12480 11630
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 10953 10364 11249 10384
rect 11009 10362 11033 10364
rect 11089 10362 11113 10364
rect 11169 10362 11193 10364
rect 11031 10310 11033 10362
rect 11095 10310 11107 10362
rect 11169 10310 11171 10362
rect 11009 10308 11033 10310
rect 11089 10308 11113 10310
rect 11169 10308 11193 10310
rect 10953 10288 11249 10308
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10612 9178 10640 9386
rect 10953 9276 11249 9296
rect 11009 9274 11033 9276
rect 11089 9274 11113 9276
rect 11169 9274 11193 9276
rect 11031 9222 11033 9274
rect 11095 9222 11107 9274
rect 11169 9222 11171 9274
rect 11009 9220 11033 9222
rect 11089 9220 11113 9222
rect 11169 9220 11193 9222
rect 10953 9200 11249 9220
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10612 8634 10640 9114
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10953 8188 11249 8208
rect 11009 8186 11033 8188
rect 11089 8186 11113 8188
rect 11169 8186 11193 8188
rect 11031 8134 11033 8186
rect 11095 8134 11107 8186
rect 11169 8134 11171 8186
rect 11009 8132 11033 8134
rect 11089 8132 11113 8134
rect 11169 8132 11193 8134
rect 10953 8112 11249 8132
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10428 6866 10456 7346
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10704 6934 10732 7142
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10888 6866 10916 7278
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 10953 7100 11249 7120
rect 11009 7098 11033 7100
rect 11089 7098 11113 7100
rect 11169 7098 11193 7100
rect 11031 7046 11033 7098
rect 11095 7046 11107 7098
rect 11169 7046 11171 7098
rect 11009 7044 11033 7046
rect 11089 7044 11113 7046
rect 11169 7044 11193 7046
rect 10953 7024 11249 7044
rect 11440 6866 11468 7142
rect 11716 6866 11744 10406
rect 11900 9994 11928 10542
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12176 10062 12204 10202
rect 12268 10198 12296 10542
rect 12256 10192 12308 10198
rect 12256 10134 12308 10140
rect 12530 10160 12586 10169
rect 12530 10095 12532 10104
rect 12584 10095 12586 10104
rect 12532 10066 12584 10072
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11992 9926 12020 9998
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11808 8430 11836 9862
rect 12728 9674 12756 12038
rect 12820 10130 12848 12922
rect 14936 12782 14964 13194
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 14924 12776 14976 12782
rect 14924 12718 14976 12724
rect 13176 12368 13228 12374
rect 13176 12310 13228 12316
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13004 11014 13032 12174
rect 13188 11694 13216 12310
rect 13372 12306 13400 12718
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13740 12374 13768 12582
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 14936 12306 14964 12718
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 15028 12306 15056 12650
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 13452 11996 13748 12016
rect 13508 11994 13532 11996
rect 13588 11994 13612 11996
rect 13668 11994 13692 11996
rect 13530 11942 13532 11994
rect 13594 11942 13606 11994
rect 13668 11942 13670 11994
rect 13508 11940 13532 11942
rect 13588 11940 13612 11942
rect 13668 11940 13692 11942
rect 13452 11920 13748 11940
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 15028 11286 15056 12038
rect 15016 11280 15068 11286
rect 15016 11222 15068 11228
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 13004 10130 13032 10950
rect 13452 10908 13748 10928
rect 13508 10906 13532 10908
rect 13588 10906 13612 10908
rect 13668 10906 13692 10908
rect 13530 10854 13532 10906
rect 13594 10854 13606 10906
rect 13668 10854 13670 10906
rect 13508 10852 13532 10854
rect 13588 10852 13612 10854
rect 13668 10852 13692 10854
rect 13452 10832 13748 10852
rect 15120 10606 15148 11018
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 15028 10130 15056 10406
rect 15120 10198 15148 10542
rect 15750 10296 15806 10305
rect 15750 10231 15806 10240
rect 15108 10192 15160 10198
rect 15108 10134 15160 10140
rect 15764 10130 15792 10231
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 12820 9926 12848 10066
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 12544 9646 12756 9674
rect 12544 9042 12572 9646
rect 12912 9110 12940 9862
rect 13452 9820 13748 9840
rect 13508 9818 13532 9820
rect 13588 9818 13612 9820
rect 13668 9818 13692 9820
rect 13530 9766 13532 9818
rect 13594 9766 13606 9818
rect 13668 9766 13670 9818
rect 13508 9764 13532 9766
rect 13588 9764 13612 9766
rect 13668 9764 13692 9766
rect 13452 9744 13748 9764
rect 12900 9104 12952 9110
rect 12900 9046 12952 9052
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 12544 8498 12572 8978
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11808 7954 11836 8366
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 13096 7886 13124 8502
rect 13188 8430 13216 8978
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 13280 7954 13308 8774
rect 13372 8566 13400 8910
rect 13452 8732 13748 8752
rect 13508 8730 13532 8732
rect 13588 8730 13612 8732
rect 13668 8730 13692 8732
rect 13530 8678 13532 8730
rect 13594 8678 13606 8730
rect 13668 8678 13670 8730
rect 13508 8676 13532 8678
rect 13588 8676 13612 8678
rect 13668 8676 13692 8678
rect 13452 8656 13748 8676
rect 13360 8560 13412 8566
rect 13360 8502 13412 8508
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13464 8090 13492 8298
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13648 7954 13676 8366
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 13096 7342 13124 7822
rect 13452 7644 13748 7664
rect 13508 7642 13532 7644
rect 13588 7642 13612 7644
rect 13668 7642 13692 7644
rect 13530 7590 13532 7642
rect 13594 7590 13606 7642
rect 13668 7590 13670 7642
rect 13508 7588 13532 7590
rect 13588 7588 13612 7590
rect 13668 7588 13692 7590
rect 13452 7568 13748 7588
rect 13832 7342 13860 9862
rect 15304 9518 15332 9862
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14200 8430 14228 8774
rect 15120 8430 15148 9386
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 14568 7342 14596 8366
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14752 8090 14780 8230
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11716 6254 11744 6802
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 12360 6186 12388 6734
rect 12912 6254 12940 6734
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 13096 6186 13124 7278
rect 14752 7274 14780 7890
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 15028 7478 15056 7686
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 14740 7268 14792 7274
rect 14740 7210 14792 7216
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 13188 6322 13216 6802
rect 13452 6556 13748 6576
rect 13508 6554 13532 6556
rect 13588 6554 13612 6556
rect 13668 6554 13692 6556
rect 13530 6502 13532 6554
rect 13594 6502 13606 6554
rect 13668 6502 13670 6554
rect 13508 6500 13532 6502
rect 13588 6500 13612 6502
rect 13668 6500 13692 6502
rect 13452 6480 13748 6500
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 10953 6012 11249 6032
rect 11009 6010 11033 6012
rect 11089 6010 11113 6012
rect 11169 6010 11193 6012
rect 11031 5958 11033 6010
rect 11095 5958 11107 6010
rect 11169 5958 11171 6010
rect 11009 5956 11033 5958
rect 11089 5956 11113 5958
rect 11169 5956 11193 5958
rect 10953 5936 11249 5956
rect 12360 5778 12388 6122
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5778 13860 6054
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10324 5296 10376 5302
rect 10324 5238 10376 5244
rect 10796 5166 10824 5510
rect 11072 5250 11100 5714
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11256 5370 11284 5510
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 10888 5234 11100 5250
rect 10876 5228 11100 5234
rect 10928 5222 11100 5228
rect 10876 5170 10928 5176
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 7012 3538 7064 3544
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6840 2650 6868 2926
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 7024 2582 7052 3334
rect 7116 3194 7144 3470
rect 7196 3460 7248 3466
rect 7196 3402 7248 3408
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7208 2582 7236 3402
rect 7300 3398 7328 3590
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7392 2854 7420 3470
rect 7668 3058 7696 3470
rect 8454 3292 8750 3312
rect 8510 3290 8534 3292
rect 8590 3290 8614 3292
rect 8670 3290 8694 3292
rect 8532 3238 8534 3290
rect 8596 3238 8608 3290
rect 8670 3238 8672 3290
rect 8510 3236 8534 3238
rect 8590 3236 8614 3238
rect 8670 3236 8694 3238
rect 8454 3216 8750 3236
rect 9140 3194 9168 5034
rect 9324 4826 9352 5034
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 9232 3194 9260 3606
rect 9324 3602 9352 3946
rect 9312 3596 9364 3602
rect 9416 3584 9444 5102
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9600 4826 9628 4966
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9876 4554 9904 5102
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10336 4758 10364 4966
rect 10324 4752 10376 4758
rect 10888 4740 10916 5170
rect 10953 4924 11249 4944
rect 11009 4922 11033 4924
rect 11089 4922 11113 4924
rect 11169 4922 11193 4924
rect 11031 4870 11033 4922
rect 11095 4870 11107 4922
rect 11169 4870 11171 4922
rect 11009 4868 11033 4870
rect 11089 4868 11113 4870
rect 11169 4868 11193 4870
rect 10953 4848 11249 4868
rect 11348 4808 11376 5646
rect 12360 5234 12388 5714
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12544 5166 12572 5578
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 13452 5468 13748 5488
rect 13508 5466 13532 5468
rect 13588 5466 13612 5468
rect 13668 5466 13692 5468
rect 13530 5414 13532 5466
rect 13594 5414 13606 5466
rect 13668 5414 13670 5466
rect 13508 5412 13532 5414
rect 13588 5412 13612 5414
rect 13668 5412 13692 5414
rect 13452 5392 13748 5412
rect 14476 5234 14504 5510
rect 15580 5370 15608 9862
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 11428 5092 11480 5098
rect 11428 5034 11480 5040
rect 11612 5092 11664 5098
rect 11612 5034 11664 5040
rect 11164 4780 11376 4808
rect 10968 4752 11020 4758
rect 10888 4712 10968 4740
rect 10324 4694 10376 4700
rect 10968 4694 11020 4700
rect 11164 4622 11192 4780
rect 11440 4758 11468 5034
rect 11428 4752 11480 4758
rect 11428 4694 11480 4700
rect 11624 4690 11652 5034
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11716 4690 11744 4966
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 9876 3602 9904 4490
rect 11164 4282 11192 4558
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11624 4146 11652 4626
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 11716 4078 11744 4626
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 10953 3836 11249 3856
rect 11009 3834 11033 3836
rect 11089 3834 11113 3836
rect 11169 3834 11193 3836
rect 11031 3782 11033 3834
rect 11095 3782 11107 3834
rect 11169 3782 11171 3834
rect 11009 3780 11033 3782
rect 11089 3780 11113 3782
rect 11169 3780 11193 3782
rect 10953 3760 11249 3780
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 9496 3596 9548 3602
rect 9416 3556 9496 3584
rect 9312 3538 9364 3544
rect 9496 3538 9548 3544
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9692 3126 9720 3334
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 9784 2922 9812 3334
rect 7656 2916 7708 2922
rect 7656 2858 7708 2864
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 7668 2650 7696 2858
rect 8680 2650 8708 2858
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 10060 2514 10088 3538
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 11072 3058 11100 3334
rect 11164 3194 11192 3470
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10953 2748 11249 2768
rect 11009 2746 11033 2748
rect 11089 2746 11113 2748
rect 11169 2746 11193 2748
rect 11031 2694 11033 2746
rect 11095 2694 11107 2746
rect 11169 2694 11171 2746
rect 11009 2692 11033 2694
rect 11089 2692 11113 2694
rect 11169 2692 11193 2694
rect 10953 2672 11249 2692
rect 11532 2650 11560 3606
rect 11716 2922 11744 4014
rect 11900 4010 11928 5102
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12084 4486 12112 4558
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 12084 4078 12112 4422
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11900 3534 11928 3946
rect 11992 3738 12020 4014
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11900 2990 11928 3470
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 11704 2916 11756 2922
rect 11704 2858 11756 2864
rect 12176 2650 12204 5102
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 12452 3058 12480 4218
rect 12544 3670 12572 5102
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13004 4758 13032 4966
rect 13188 4758 13216 5102
rect 12992 4752 13044 4758
rect 12992 4694 13044 4700
rect 13176 4752 13228 4758
rect 13176 4694 13228 4700
rect 13740 4690 13768 5170
rect 14096 5092 14148 5098
rect 14096 5034 14148 5040
rect 14188 5092 14240 5098
rect 14188 5034 14240 5040
rect 14108 4690 14136 5034
rect 14200 4826 14228 5034
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 15580 4690 15608 4966
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 13740 4468 13768 4626
rect 15752 4548 15804 4554
rect 15752 4490 15804 4496
rect 13740 4440 13860 4468
rect 13452 4380 13748 4400
rect 13508 4378 13532 4380
rect 13588 4378 13612 4380
rect 13668 4378 13692 4380
rect 13530 4326 13532 4378
rect 13594 4326 13606 4378
rect 13668 4326 13670 4378
rect 13508 4324 13532 4326
rect 13588 4324 13612 4326
rect 13668 4324 13692 4326
rect 13452 4304 13748 4324
rect 13832 4282 13860 4440
rect 15764 4282 15792 4490
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 13832 4146 13860 4218
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13556 3670 13584 3878
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12544 2774 12572 3606
rect 13832 3602 13860 4082
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13452 3292 13748 3312
rect 13508 3290 13532 3292
rect 13588 3290 13612 3292
rect 13668 3290 13692 3292
rect 13530 3238 13532 3290
rect 13594 3238 13606 3290
rect 13668 3238 13670 3290
rect 13508 3236 13532 3238
rect 13588 3236 13612 3238
rect 13668 3236 13692 3238
rect 13452 3216 13748 3236
rect 14292 3194 14320 3946
rect 14936 3194 14964 3946
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 13820 2916 13872 2922
rect 13820 2858 13872 2864
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 12452 2746 12572 2774
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 12452 2514 12480 2746
rect 13740 2514 13768 2790
rect 13832 2650 13860 2858
rect 15580 2650 15608 2994
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 15568 2644 15620 2650
rect 15568 2586 15620 2592
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 15752 2508 15804 2514
rect 15752 2450 15804 2456
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 3455 2204 3751 2224
rect 3511 2202 3535 2204
rect 3591 2202 3615 2204
rect 3671 2202 3695 2204
rect 3533 2150 3535 2202
rect 3597 2150 3609 2202
rect 3671 2150 3673 2202
rect 3511 2148 3535 2150
rect 3591 2148 3615 2150
rect 3671 2148 3695 2150
rect 3455 2128 3751 2148
rect 6012 800 6040 2314
rect 8454 2204 8750 2224
rect 8510 2202 8534 2204
rect 8590 2202 8614 2204
rect 8670 2202 8694 2204
rect 8532 2150 8534 2202
rect 8596 2150 8608 2202
rect 8670 2150 8672 2202
rect 8510 2148 8534 2150
rect 8590 2148 8614 2150
rect 8670 2148 8694 2150
rect 8454 2128 8750 2148
rect 11992 800 12020 2450
rect 13452 2204 13748 2224
rect 13508 2202 13532 2204
rect 13588 2202 13612 2204
rect 13668 2202 13692 2204
rect 13530 2150 13532 2202
rect 13594 2150 13606 2202
rect 13668 2150 13670 2202
rect 13508 2148 13532 2150
rect 13588 2148 13612 2150
rect 13668 2148 13692 2150
rect 13452 2128 13748 2148
rect 15764 1465 15792 2450
rect 15750 1456 15806 1465
rect 15750 1391 15806 1400
rect 478 0 534 800
rect 5998 0 6054 800
rect 11978 0 12034 800
<< via2 >>
rect 1398 17720 1454 17776
rect 1398 8880 1454 8936
rect 3455 16346 3511 16348
rect 3535 16346 3591 16348
rect 3615 16346 3671 16348
rect 3695 16346 3751 16348
rect 3455 16294 3481 16346
rect 3481 16294 3511 16346
rect 3535 16294 3545 16346
rect 3545 16294 3591 16346
rect 3615 16294 3661 16346
rect 3661 16294 3671 16346
rect 3695 16294 3725 16346
rect 3725 16294 3751 16346
rect 3455 16292 3511 16294
rect 3535 16292 3591 16294
rect 3615 16292 3671 16294
rect 3695 16292 3751 16294
rect 3455 15258 3511 15260
rect 3535 15258 3591 15260
rect 3615 15258 3671 15260
rect 3695 15258 3751 15260
rect 3455 15206 3481 15258
rect 3481 15206 3511 15258
rect 3535 15206 3545 15258
rect 3545 15206 3591 15258
rect 3615 15206 3661 15258
rect 3661 15206 3671 15258
rect 3695 15206 3725 15258
rect 3725 15206 3751 15258
rect 3455 15204 3511 15206
rect 3535 15204 3591 15206
rect 3615 15204 3671 15206
rect 3695 15204 3751 15206
rect 3455 14170 3511 14172
rect 3535 14170 3591 14172
rect 3615 14170 3671 14172
rect 3695 14170 3751 14172
rect 3455 14118 3481 14170
rect 3481 14118 3511 14170
rect 3535 14118 3545 14170
rect 3545 14118 3591 14170
rect 3615 14118 3661 14170
rect 3661 14118 3671 14170
rect 3695 14118 3725 14170
rect 3725 14118 3751 14170
rect 3455 14116 3511 14118
rect 3535 14116 3591 14118
rect 3615 14116 3671 14118
rect 3695 14116 3751 14118
rect 3455 13082 3511 13084
rect 3535 13082 3591 13084
rect 3615 13082 3671 13084
rect 3695 13082 3751 13084
rect 3455 13030 3481 13082
rect 3481 13030 3511 13082
rect 3535 13030 3545 13082
rect 3545 13030 3591 13082
rect 3615 13030 3661 13082
rect 3661 13030 3671 13082
rect 3695 13030 3725 13082
rect 3725 13030 3751 13082
rect 3455 13028 3511 13030
rect 3535 13028 3591 13030
rect 3615 13028 3671 13030
rect 3695 13028 3751 13030
rect 3455 11994 3511 11996
rect 3535 11994 3591 11996
rect 3615 11994 3671 11996
rect 3695 11994 3751 11996
rect 3455 11942 3481 11994
rect 3481 11942 3511 11994
rect 3535 11942 3545 11994
rect 3545 11942 3591 11994
rect 3615 11942 3661 11994
rect 3661 11942 3671 11994
rect 3695 11942 3725 11994
rect 3725 11942 3751 11994
rect 3455 11940 3511 11942
rect 3535 11940 3591 11942
rect 3615 11940 3671 11942
rect 3695 11940 3751 11942
rect 3455 10906 3511 10908
rect 3535 10906 3591 10908
rect 3615 10906 3671 10908
rect 3695 10906 3751 10908
rect 3455 10854 3481 10906
rect 3481 10854 3511 10906
rect 3535 10854 3545 10906
rect 3545 10854 3591 10906
rect 3615 10854 3661 10906
rect 3661 10854 3671 10906
rect 3695 10854 3725 10906
rect 3725 10854 3751 10906
rect 3455 10852 3511 10854
rect 3535 10852 3591 10854
rect 3615 10852 3671 10854
rect 3695 10852 3751 10854
rect 3455 9818 3511 9820
rect 3535 9818 3591 9820
rect 3615 9818 3671 9820
rect 3695 9818 3751 9820
rect 3455 9766 3481 9818
rect 3481 9766 3511 9818
rect 3535 9766 3545 9818
rect 3545 9766 3591 9818
rect 3615 9766 3661 9818
rect 3661 9766 3671 9818
rect 3695 9766 3725 9818
rect 3725 9766 3751 9818
rect 3455 9764 3511 9766
rect 3535 9764 3591 9766
rect 3615 9764 3671 9766
rect 3695 9764 3751 9766
rect 3455 8730 3511 8732
rect 3535 8730 3591 8732
rect 3615 8730 3671 8732
rect 3695 8730 3751 8732
rect 3455 8678 3481 8730
rect 3481 8678 3511 8730
rect 3535 8678 3545 8730
rect 3545 8678 3591 8730
rect 3615 8678 3661 8730
rect 3661 8678 3671 8730
rect 3695 8678 3725 8730
rect 3725 8678 3751 8730
rect 3455 8676 3511 8678
rect 3535 8676 3591 8678
rect 3615 8676 3671 8678
rect 3695 8676 3751 8678
rect 3455 7642 3511 7644
rect 3535 7642 3591 7644
rect 3615 7642 3671 7644
rect 3695 7642 3751 7644
rect 3455 7590 3481 7642
rect 3481 7590 3511 7642
rect 3535 7590 3545 7642
rect 3545 7590 3591 7642
rect 3615 7590 3661 7642
rect 3661 7590 3671 7642
rect 3695 7590 3725 7642
rect 3725 7590 3751 7642
rect 3455 7588 3511 7590
rect 3535 7588 3591 7590
rect 3615 7588 3671 7590
rect 3695 7588 3751 7590
rect 5954 16890 6010 16892
rect 6034 16890 6090 16892
rect 6114 16890 6170 16892
rect 6194 16890 6250 16892
rect 5954 16838 5980 16890
rect 5980 16838 6010 16890
rect 6034 16838 6044 16890
rect 6044 16838 6090 16890
rect 6114 16838 6160 16890
rect 6160 16838 6170 16890
rect 6194 16838 6224 16890
rect 6224 16838 6250 16890
rect 5954 16836 6010 16838
rect 6034 16836 6090 16838
rect 6114 16836 6170 16838
rect 6194 16836 6250 16838
rect 10953 16890 11009 16892
rect 11033 16890 11089 16892
rect 11113 16890 11169 16892
rect 11193 16890 11249 16892
rect 10953 16838 10979 16890
rect 10979 16838 11009 16890
rect 11033 16838 11043 16890
rect 11043 16838 11089 16890
rect 11113 16838 11159 16890
rect 11159 16838 11169 16890
rect 11193 16838 11223 16890
rect 11223 16838 11249 16890
rect 10953 16836 11009 16838
rect 11033 16836 11089 16838
rect 11113 16836 11169 16838
rect 11193 16836 11249 16838
rect 5954 15802 6010 15804
rect 6034 15802 6090 15804
rect 6114 15802 6170 15804
rect 6194 15802 6250 15804
rect 5954 15750 5980 15802
rect 5980 15750 6010 15802
rect 6034 15750 6044 15802
rect 6044 15750 6090 15802
rect 6114 15750 6160 15802
rect 6160 15750 6170 15802
rect 6194 15750 6224 15802
rect 6224 15750 6250 15802
rect 5954 15748 6010 15750
rect 6034 15748 6090 15750
rect 6114 15748 6170 15750
rect 6194 15748 6250 15750
rect 5954 14714 6010 14716
rect 6034 14714 6090 14716
rect 6114 14714 6170 14716
rect 6194 14714 6250 14716
rect 5954 14662 5980 14714
rect 5980 14662 6010 14714
rect 6034 14662 6044 14714
rect 6044 14662 6090 14714
rect 6114 14662 6160 14714
rect 6160 14662 6170 14714
rect 6194 14662 6224 14714
rect 6224 14662 6250 14714
rect 5954 14660 6010 14662
rect 6034 14660 6090 14662
rect 6114 14660 6170 14662
rect 6194 14660 6250 14662
rect 5954 13626 6010 13628
rect 6034 13626 6090 13628
rect 6114 13626 6170 13628
rect 6194 13626 6250 13628
rect 5954 13574 5980 13626
rect 5980 13574 6010 13626
rect 6034 13574 6044 13626
rect 6044 13574 6090 13626
rect 6114 13574 6160 13626
rect 6160 13574 6170 13626
rect 6194 13574 6224 13626
rect 6224 13574 6250 13626
rect 5954 13572 6010 13574
rect 6034 13572 6090 13574
rect 6114 13572 6170 13574
rect 6194 13572 6250 13574
rect 5954 12538 6010 12540
rect 6034 12538 6090 12540
rect 6114 12538 6170 12540
rect 6194 12538 6250 12540
rect 5954 12486 5980 12538
rect 5980 12486 6010 12538
rect 6034 12486 6044 12538
rect 6044 12486 6090 12538
rect 6114 12486 6160 12538
rect 6160 12486 6170 12538
rect 6194 12486 6224 12538
rect 6224 12486 6250 12538
rect 5954 12484 6010 12486
rect 6034 12484 6090 12486
rect 6114 12484 6170 12486
rect 6194 12484 6250 12486
rect 8454 16346 8510 16348
rect 8534 16346 8590 16348
rect 8614 16346 8670 16348
rect 8694 16346 8750 16348
rect 8454 16294 8480 16346
rect 8480 16294 8510 16346
rect 8534 16294 8544 16346
rect 8544 16294 8590 16346
rect 8614 16294 8660 16346
rect 8660 16294 8670 16346
rect 8694 16294 8724 16346
rect 8724 16294 8750 16346
rect 8454 16292 8510 16294
rect 8534 16292 8590 16294
rect 8614 16292 8670 16294
rect 8694 16292 8750 16294
rect 13452 16346 13508 16348
rect 13532 16346 13588 16348
rect 13612 16346 13668 16348
rect 13692 16346 13748 16348
rect 13452 16294 13478 16346
rect 13478 16294 13508 16346
rect 13532 16294 13542 16346
rect 13542 16294 13588 16346
rect 13612 16294 13658 16346
rect 13658 16294 13668 16346
rect 13692 16294 13722 16346
rect 13722 16294 13748 16346
rect 13452 16292 13508 16294
rect 13532 16292 13588 16294
rect 13612 16292 13668 16294
rect 13692 16292 13748 16294
rect 8454 15258 8510 15260
rect 8534 15258 8590 15260
rect 8614 15258 8670 15260
rect 8694 15258 8750 15260
rect 8454 15206 8480 15258
rect 8480 15206 8510 15258
rect 8534 15206 8544 15258
rect 8544 15206 8590 15258
rect 8614 15206 8660 15258
rect 8660 15206 8670 15258
rect 8694 15206 8724 15258
rect 8724 15206 8750 15258
rect 8454 15204 8510 15206
rect 8534 15204 8590 15206
rect 8614 15204 8670 15206
rect 8694 15204 8750 15206
rect 5954 11450 6010 11452
rect 6034 11450 6090 11452
rect 6114 11450 6170 11452
rect 6194 11450 6250 11452
rect 5954 11398 5980 11450
rect 5980 11398 6010 11450
rect 6034 11398 6044 11450
rect 6044 11398 6090 11450
rect 6114 11398 6160 11450
rect 6160 11398 6170 11450
rect 6194 11398 6224 11450
rect 6224 11398 6250 11450
rect 5954 11396 6010 11398
rect 6034 11396 6090 11398
rect 6114 11396 6170 11398
rect 6194 11396 6250 11398
rect 5954 10362 6010 10364
rect 6034 10362 6090 10364
rect 6114 10362 6170 10364
rect 6194 10362 6250 10364
rect 5954 10310 5980 10362
rect 5980 10310 6010 10362
rect 6034 10310 6044 10362
rect 6044 10310 6090 10362
rect 6114 10310 6160 10362
rect 6160 10310 6170 10362
rect 6194 10310 6224 10362
rect 6224 10310 6250 10362
rect 5954 10308 6010 10310
rect 6034 10308 6090 10310
rect 6114 10308 6170 10310
rect 6194 10308 6250 10310
rect 5954 9274 6010 9276
rect 6034 9274 6090 9276
rect 6114 9274 6170 9276
rect 6194 9274 6250 9276
rect 5954 9222 5980 9274
rect 5980 9222 6010 9274
rect 6034 9222 6044 9274
rect 6044 9222 6090 9274
rect 6114 9222 6160 9274
rect 6160 9222 6170 9274
rect 6194 9222 6224 9274
rect 6224 9222 6250 9274
rect 5954 9220 6010 9222
rect 6034 9220 6090 9222
rect 6114 9220 6170 9222
rect 6194 9220 6250 9222
rect 3455 6554 3511 6556
rect 3535 6554 3591 6556
rect 3615 6554 3671 6556
rect 3695 6554 3751 6556
rect 3455 6502 3481 6554
rect 3481 6502 3511 6554
rect 3535 6502 3545 6554
rect 3545 6502 3591 6554
rect 3615 6502 3661 6554
rect 3661 6502 3671 6554
rect 3695 6502 3725 6554
rect 3725 6502 3751 6554
rect 3455 6500 3511 6502
rect 3535 6500 3591 6502
rect 3615 6500 3671 6502
rect 3695 6500 3751 6502
rect 7102 11736 7158 11792
rect 8454 14170 8510 14172
rect 8534 14170 8590 14172
rect 8614 14170 8670 14172
rect 8694 14170 8750 14172
rect 8454 14118 8480 14170
rect 8480 14118 8510 14170
rect 8534 14118 8544 14170
rect 8544 14118 8590 14170
rect 8614 14118 8660 14170
rect 8660 14118 8670 14170
rect 8694 14118 8724 14170
rect 8724 14118 8750 14170
rect 8454 14116 8510 14118
rect 8534 14116 8590 14118
rect 8614 14116 8670 14118
rect 8694 14116 8750 14118
rect 9218 13776 9274 13832
rect 8454 13082 8510 13084
rect 8534 13082 8590 13084
rect 8614 13082 8670 13084
rect 8694 13082 8750 13084
rect 8454 13030 8480 13082
rect 8480 13030 8510 13082
rect 8534 13030 8544 13082
rect 8544 13030 8590 13082
rect 8614 13030 8660 13082
rect 8660 13030 8670 13082
rect 8694 13030 8724 13082
rect 8724 13030 8750 13082
rect 8454 13028 8510 13030
rect 8534 13028 8590 13030
rect 8614 13028 8670 13030
rect 8694 13028 8750 13030
rect 8114 12144 8170 12200
rect 8454 11994 8510 11996
rect 8534 11994 8590 11996
rect 8614 11994 8670 11996
rect 8694 11994 8750 11996
rect 8454 11942 8480 11994
rect 8480 11942 8510 11994
rect 8534 11942 8544 11994
rect 8544 11942 8590 11994
rect 8614 11942 8660 11994
rect 8660 11942 8670 11994
rect 8694 11942 8724 11994
rect 8724 11942 8750 11994
rect 8454 11940 8510 11942
rect 8534 11940 8590 11942
rect 8614 11940 8670 11942
rect 8694 11940 8750 11942
rect 8454 10906 8510 10908
rect 8534 10906 8590 10908
rect 8614 10906 8670 10908
rect 8694 10906 8750 10908
rect 8454 10854 8480 10906
rect 8480 10854 8510 10906
rect 8534 10854 8544 10906
rect 8544 10854 8590 10906
rect 8614 10854 8660 10906
rect 8660 10854 8670 10906
rect 8694 10854 8724 10906
rect 8724 10854 8750 10906
rect 8454 10852 8510 10854
rect 8534 10852 8590 10854
rect 8614 10852 8670 10854
rect 8694 10852 8750 10854
rect 5954 8186 6010 8188
rect 6034 8186 6090 8188
rect 6114 8186 6170 8188
rect 6194 8186 6250 8188
rect 5954 8134 5980 8186
rect 5980 8134 6010 8186
rect 6034 8134 6044 8186
rect 6044 8134 6090 8186
rect 6114 8134 6160 8186
rect 6160 8134 6170 8186
rect 6194 8134 6224 8186
rect 6224 8134 6250 8186
rect 5954 8132 6010 8134
rect 6034 8132 6090 8134
rect 6114 8132 6170 8134
rect 6194 8132 6250 8134
rect 3455 5466 3511 5468
rect 3535 5466 3591 5468
rect 3615 5466 3671 5468
rect 3695 5466 3751 5468
rect 3455 5414 3481 5466
rect 3481 5414 3511 5466
rect 3535 5414 3545 5466
rect 3545 5414 3591 5466
rect 3615 5414 3661 5466
rect 3661 5414 3671 5466
rect 3695 5414 3725 5466
rect 3725 5414 3751 5466
rect 3455 5412 3511 5414
rect 3535 5412 3591 5414
rect 3615 5412 3671 5414
rect 3695 5412 3751 5414
rect 3455 4378 3511 4380
rect 3535 4378 3591 4380
rect 3615 4378 3671 4380
rect 3695 4378 3751 4380
rect 3455 4326 3481 4378
rect 3481 4326 3511 4378
rect 3535 4326 3545 4378
rect 3545 4326 3591 4378
rect 3615 4326 3661 4378
rect 3661 4326 3671 4378
rect 3695 4326 3725 4378
rect 3725 4326 3751 4378
rect 3455 4324 3511 4326
rect 3535 4324 3591 4326
rect 3615 4324 3671 4326
rect 3695 4324 3751 4326
rect 3455 3290 3511 3292
rect 3535 3290 3591 3292
rect 3615 3290 3671 3292
rect 3695 3290 3751 3292
rect 3455 3238 3481 3290
rect 3481 3238 3511 3290
rect 3535 3238 3545 3290
rect 3545 3238 3591 3290
rect 3615 3238 3661 3290
rect 3661 3238 3671 3290
rect 3695 3238 3725 3290
rect 3725 3238 3751 3290
rect 3455 3236 3511 3238
rect 3535 3236 3591 3238
rect 3615 3236 3671 3238
rect 3695 3236 3751 3238
rect 5954 7098 6010 7100
rect 6034 7098 6090 7100
rect 6114 7098 6170 7100
rect 6194 7098 6250 7100
rect 5954 7046 5980 7098
rect 5980 7046 6010 7098
rect 6034 7046 6044 7098
rect 6044 7046 6090 7098
rect 6114 7046 6160 7098
rect 6160 7046 6170 7098
rect 6194 7046 6224 7098
rect 6224 7046 6250 7098
rect 5954 7044 6010 7046
rect 6034 7044 6090 7046
rect 6114 7044 6170 7046
rect 6194 7044 6250 7046
rect 5954 6010 6010 6012
rect 6034 6010 6090 6012
rect 6114 6010 6170 6012
rect 6194 6010 6250 6012
rect 5954 5958 5980 6010
rect 5980 5958 6010 6010
rect 6034 5958 6044 6010
rect 6044 5958 6090 6010
rect 6114 5958 6160 6010
rect 6160 5958 6170 6010
rect 6194 5958 6224 6010
rect 6224 5958 6250 6010
rect 5954 5956 6010 5958
rect 6034 5956 6090 5958
rect 6114 5956 6170 5958
rect 6194 5956 6250 5958
rect 8454 9818 8510 9820
rect 8534 9818 8590 9820
rect 8614 9818 8670 9820
rect 8694 9818 8750 9820
rect 8454 9766 8480 9818
rect 8480 9766 8510 9818
rect 8534 9766 8544 9818
rect 8544 9766 8590 9818
rect 8614 9766 8660 9818
rect 8660 9766 8670 9818
rect 8694 9766 8724 9818
rect 8724 9766 8750 9818
rect 8454 9764 8510 9766
rect 8534 9764 8590 9766
rect 8614 9764 8670 9766
rect 8694 9764 8750 9766
rect 9586 11736 9642 11792
rect 10953 15802 11009 15804
rect 11033 15802 11089 15804
rect 11113 15802 11169 15804
rect 11193 15802 11249 15804
rect 10953 15750 10979 15802
rect 10979 15750 11009 15802
rect 11033 15750 11043 15802
rect 11043 15750 11089 15802
rect 11113 15750 11159 15802
rect 11159 15750 11169 15802
rect 11193 15750 11223 15802
rect 11223 15750 11249 15802
rect 10953 15748 11009 15750
rect 11033 15748 11089 15750
rect 11113 15748 11169 15750
rect 11193 15748 11249 15750
rect 10953 14714 11009 14716
rect 11033 14714 11089 14716
rect 11113 14714 11169 14716
rect 11193 14714 11249 14716
rect 10953 14662 10979 14714
rect 10979 14662 11009 14714
rect 11033 14662 11043 14714
rect 11043 14662 11089 14714
rect 11113 14662 11159 14714
rect 11159 14662 11169 14714
rect 11193 14662 11223 14714
rect 11223 14662 11249 14714
rect 10953 14660 11009 14662
rect 11033 14660 11089 14662
rect 11113 14660 11169 14662
rect 11193 14660 11249 14662
rect 9954 13812 9956 13832
rect 9956 13812 10008 13832
rect 10008 13812 10010 13832
rect 9954 13776 10010 13812
rect 10953 13626 11009 13628
rect 11033 13626 11089 13628
rect 11113 13626 11169 13628
rect 11193 13626 11249 13628
rect 10953 13574 10979 13626
rect 10979 13574 11009 13626
rect 11033 13574 11043 13626
rect 11043 13574 11089 13626
rect 11113 13574 11159 13626
rect 11159 13574 11169 13626
rect 11193 13574 11223 13626
rect 11223 13574 11249 13626
rect 10953 13572 11009 13574
rect 11033 13572 11089 13574
rect 11113 13572 11169 13574
rect 11193 13572 11249 13574
rect 10953 12538 11009 12540
rect 11033 12538 11089 12540
rect 11113 12538 11169 12540
rect 11193 12538 11249 12540
rect 10953 12486 10979 12538
rect 10979 12486 11009 12538
rect 11033 12486 11043 12538
rect 11043 12486 11089 12538
rect 11113 12486 11159 12538
rect 11159 12486 11169 12538
rect 11193 12486 11223 12538
rect 11223 12486 11249 12538
rect 10953 12484 11009 12486
rect 11033 12484 11089 12486
rect 11113 12484 11169 12486
rect 11193 12484 11249 12486
rect 10230 12164 10286 12200
rect 10230 12144 10232 12164
rect 10232 12144 10284 12164
rect 10284 12144 10286 12164
rect 9954 10124 10010 10160
rect 9954 10104 9956 10124
rect 9956 10104 10008 10124
rect 10008 10104 10010 10124
rect 8454 8730 8510 8732
rect 8534 8730 8590 8732
rect 8614 8730 8670 8732
rect 8694 8730 8750 8732
rect 8454 8678 8480 8730
rect 8480 8678 8510 8730
rect 8534 8678 8544 8730
rect 8544 8678 8590 8730
rect 8614 8678 8660 8730
rect 8660 8678 8670 8730
rect 8694 8678 8724 8730
rect 8724 8678 8750 8730
rect 8454 8676 8510 8678
rect 8534 8676 8590 8678
rect 8614 8676 8670 8678
rect 8694 8676 8750 8678
rect 8454 7642 8510 7644
rect 8534 7642 8590 7644
rect 8614 7642 8670 7644
rect 8694 7642 8750 7644
rect 8454 7590 8480 7642
rect 8480 7590 8510 7642
rect 8534 7590 8544 7642
rect 8544 7590 8590 7642
rect 8614 7590 8660 7642
rect 8660 7590 8670 7642
rect 8694 7590 8724 7642
rect 8724 7590 8750 7642
rect 8454 7588 8510 7590
rect 8534 7588 8590 7590
rect 8614 7588 8670 7590
rect 8694 7588 8750 7590
rect 8454 6554 8510 6556
rect 8534 6554 8590 6556
rect 8614 6554 8670 6556
rect 8694 6554 8750 6556
rect 8454 6502 8480 6554
rect 8480 6502 8510 6554
rect 8534 6502 8544 6554
rect 8544 6502 8590 6554
rect 8614 6502 8660 6554
rect 8660 6502 8670 6554
rect 8694 6502 8724 6554
rect 8724 6502 8750 6554
rect 8454 6500 8510 6502
rect 8534 6500 8590 6502
rect 8614 6500 8670 6502
rect 8694 6500 8750 6502
rect 5954 4922 6010 4924
rect 6034 4922 6090 4924
rect 6114 4922 6170 4924
rect 6194 4922 6250 4924
rect 5954 4870 5980 4922
rect 5980 4870 6010 4922
rect 6034 4870 6044 4922
rect 6044 4870 6090 4922
rect 6114 4870 6160 4922
rect 6160 4870 6170 4922
rect 6194 4870 6224 4922
rect 6224 4870 6250 4922
rect 5954 4868 6010 4870
rect 6034 4868 6090 4870
rect 6114 4868 6170 4870
rect 6194 4868 6250 4870
rect 5954 3834 6010 3836
rect 6034 3834 6090 3836
rect 6114 3834 6170 3836
rect 6194 3834 6250 3836
rect 5954 3782 5980 3834
rect 5980 3782 6010 3834
rect 6034 3782 6044 3834
rect 6044 3782 6090 3834
rect 6114 3782 6160 3834
rect 6160 3782 6170 3834
rect 6194 3782 6224 3834
rect 6224 3782 6250 3834
rect 5954 3780 6010 3782
rect 6034 3780 6090 3782
rect 6114 3780 6170 3782
rect 6194 3780 6250 3782
rect 5954 2746 6010 2748
rect 6034 2746 6090 2748
rect 6114 2746 6170 2748
rect 6194 2746 6250 2748
rect 5954 2694 5980 2746
rect 5980 2694 6010 2746
rect 6034 2694 6044 2746
rect 6044 2694 6090 2746
rect 6114 2694 6160 2746
rect 6160 2694 6170 2746
rect 6194 2694 6224 2746
rect 6224 2694 6250 2746
rect 5954 2692 6010 2694
rect 6034 2692 6090 2694
rect 6114 2692 6170 2694
rect 6194 2692 6250 2694
rect 8454 5466 8510 5468
rect 8534 5466 8590 5468
rect 8614 5466 8670 5468
rect 8694 5466 8750 5468
rect 8454 5414 8480 5466
rect 8480 5414 8510 5466
rect 8534 5414 8544 5466
rect 8544 5414 8590 5466
rect 8614 5414 8660 5466
rect 8660 5414 8670 5466
rect 8694 5414 8724 5466
rect 8724 5414 8750 5466
rect 8454 5412 8510 5414
rect 8534 5412 8590 5414
rect 8614 5412 8670 5414
rect 8694 5412 8750 5414
rect 8454 4378 8510 4380
rect 8534 4378 8590 4380
rect 8614 4378 8670 4380
rect 8694 4378 8750 4380
rect 8454 4326 8480 4378
rect 8480 4326 8510 4378
rect 8534 4326 8544 4378
rect 8544 4326 8590 4378
rect 8614 4326 8660 4378
rect 8660 4326 8670 4378
rect 8694 4326 8724 4378
rect 8724 4326 8750 4378
rect 8454 4324 8510 4326
rect 8534 4324 8590 4326
rect 8614 4324 8670 4326
rect 8694 4324 8750 4326
rect 10953 11450 11009 11452
rect 11033 11450 11089 11452
rect 11113 11450 11169 11452
rect 11193 11450 11249 11452
rect 10953 11398 10979 11450
rect 10979 11398 11009 11450
rect 11033 11398 11043 11450
rect 11043 11398 11089 11450
rect 11113 11398 11159 11450
rect 11159 11398 11169 11450
rect 11193 11398 11223 11450
rect 11223 11398 11249 11450
rect 10953 11396 11009 11398
rect 11033 11396 11089 11398
rect 11113 11396 11169 11398
rect 11193 11396 11249 11398
rect 13452 15258 13508 15260
rect 13532 15258 13588 15260
rect 13612 15258 13668 15260
rect 13692 15258 13748 15260
rect 13452 15206 13478 15258
rect 13478 15206 13508 15258
rect 13532 15206 13542 15258
rect 13542 15206 13588 15258
rect 13612 15206 13658 15258
rect 13658 15206 13668 15258
rect 13692 15206 13722 15258
rect 13722 15206 13748 15258
rect 13452 15204 13508 15206
rect 13532 15204 13588 15206
rect 13612 15204 13668 15206
rect 13692 15204 13748 15206
rect 13452 14170 13508 14172
rect 13532 14170 13588 14172
rect 13612 14170 13668 14172
rect 13692 14170 13748 14172
rect 13452 14118 13478 14170
rect 13478 14118 13508 14170
rect 13532 14118 13542 14170
rect 13542 14118 13588 14170
rect 13612 14118 13658 14170
rect 13658 14118 13668 14170
rect 13692 14118 13722 14170
rect 13722 14118 13748 14170
rect 13452 14116 13508 14118
rect 13532 14116 13588 14118
rect 13612 14116 13668 14118
rect 13692 14116 13748 14118
rect 13452 13082 13508 13084
rect 13532 13082 13588 13084
rect 13612 13082 13668 13084
rect 13692 13082 13748 13084
rect 13452 13030 13478 13082
rect 13478 13030 13508 13082
rect 13532 13030 13542 13082
rect 13542 13030 13588 13082
rect 13612 13030 13658 13082
rect 13658 13030 13668 13082
rect 13692 13030 13722 13082
rect 13722 13030 13748 13082
rect 13452 13028 13508 13030
rect 13532 13028 13588 13030
rect 13612 13028 13668 13030
rect 13692 13028 13748 13030
rect 10953 10362 11009 10364
rect 11033 10362 11089 10364
rect 11113 10362 11169 10364
rect 11193 10362 11249 10364
rect 10953 10310 10979 10362
rect 10979 10310 11009 10362
rect 11033 10310 11043 10362
rect 11043 10310 11089 10362
rect 11113 10310 11159 10362
rect 11159 10310 11169 10362
rect 11193 10310 11223 10362
rect 11223 10310 11249 10362
rect 10953 10308 11009 10310
rect 11033 10308 11089 10310
rect 11113 10308 11169 10310
rect 11193 10308 11249 10310
rect 10953 9274 11009 9276
rect 11033 9274 11089 9276
rect 11113 9274 11169 9276
rect 11193 9274 11249 9276
rect 10953 9222 10979 9274
rect 10979 9222 11009 9274
rect 11033 9222 11043 9274
rect 11043 9222 11089 9274
rect 11113 9222 11159 9274
rect 11159 9222 11169 9274
rect 11193 9222 11223 9274
rect 11223 9222 11249 9274
rect 10953 9220 11009 9222
rect 11033 9220 11089 9222
rect 11113 9220 11169 9222
rect 11193 9220 11249 9222
rect 10953 8186 11009 8188
rect 11033 8186 11089 8188
rect 11113 8186 11169 8188
rect 11193 8186 11249 8188
rect 10953 8134 10979 8186
rect 10979 8134 11009 8186
rect 11033 8134 11043 8186
rect 11043 8134 11089 8186
rect 11113 8134 11159 8186
rect 11159 8134 11169 8186
rect 11193 8134 11223 8186
rect 11223 8134 11249 8186
rect 10953 8132 11009 8134
rect 11033 8132 11089 8134
rect 11113 8132 11169 8134
rect 11193 8132 11249 8134
rect 10953 7098 11009 7100
rect 11033 7098 11089 7100
rect 11113 7098 11169 7100
rect 11193 7098 11249 7100
rect 10953 7046 10979 7098
rect 10979 7046 11009 7098
rect 11033 7046 11043 7098
rect 11043 7046 11089 7098
rect 11113 7046 11159 7098
rect 11159 7046 11169 7098
rect 11193 7046 11223 7098
rect 11223 7046 11249 7098
rect 10953 7044 11009 7046
rect 11033 7044 11089 7046
rect 11113 7044 11169 7046
rect 11193 7044 11249 7046
rect 12530 10124 12586 10160
rect 12530 10104 12532 10124
rect 12532 10104 12584 10124
rect 12584 10104 12586 10124
rect 13452 11994 13508 11996
rect 13532 11994 13588 11996
rect 13612 11994 13668 11996
rect 13692 11994 13748 11996
rect 13452 11942 13478 11994
rect 13478 11942 13508 11994
rect 13532 11942 13542 11994
rect 13542 11942 13588 11994
rect 13612 11942 13658 11994
rect 13658 11942 13668 11994
rect 13692 11942 13722 11994
rect 13722 11942 13748 11994
rect 13452 11940 13508 11942
rect 13532 11940 13588 11942
rect 13612 11940 13668 11942
rect 13692 11940 13748 11942
rect 13452 10906 13508 10908
rect 13532 10906 13588 10908
rect 13612 10906 13668 10908
rect 13692 10906 13748 10908
rect 13452 10854 13478 10906
rect 13478 10854 13508 10906
rect 13532 10854 13542 10906
rect 13542 10854 13588 10906
rect 13612 10854 13658 10906
rect 13658 10854 13668 10906
rect 13692 10854 13722 10906
rect 13722 10854 13748 10906
rect 13452 10852 13508 10854
rect 13532 10852 13588 10854
rect 13612 10852 13668 10854
rect 13692 10852 13748 10854
rect 15750 10240 15806 10296
rect 13452 9818 13508 9820
rect 13532 9818 13588 9820
rect 13612 9818 13668 9820
rect 13692 9818 13748 9820
rect 13452 9766 13478 9818
rect 13478 9766 13508 9818
rect 13532 9766 13542 9818
rect 13542 9766 13588 9818
rect 13612 9766 13658 9818
rect 13658 9766 13668 9818
rect 13692 9766 13722 9818
rect 13722 9766 13748 9818
rect 13452 9764 13508 9766
rect 13532 9764 13588 9766
rect 13612 9764 13668 9766
rect 13692 9764 13748 9766
rect 13452 8730 13508 8732
rect 13532 8730 13588 8732
rect 13612 8730 13668 8732
rect 13692 8730 13748 8732
rect 13452 8678 13478 8730
rect 13478 8678 13508 8730
rect 13532 8678 13542 8730
rect 13542 8678 13588 8730
rect 13612 8678 13658 8730
rect 13658 8678 13668 8730
rect 13692 8678 13722 8730
rect 13722 8678 13748 8730
rect 13452 8676 13508 8678
rect 13532 8676 13588 8678
rect 13612 8676 13668 8678
rect 13692 8676 13748 8678
rect 13452 7642 13508 7644
rect 13532 7642 13588 7644
rect 13612 7642 13668 7644
rect 13692 7642 13748 7644
rect 13452 7590 13478 7642
rect 13478 7590 13508 7642
rect 13532 7590 13542 7642
rect 13542 7590 13588 7642
rect 13612 7590 13658 7642
rect 13658 7590 13668 7642
rect 13692 7590 13722 7642
rect 13722 7590 13748 7642
rect 13452 7588 13508 7590
rect 13532 7588 13588 7590
rect 13612 7588 13668 7590
rect 13692 7588 13748 7590
rect 13452 6554 13508 6556
rect 13532 6554 13588 6556
rect 13612 6554 13668 6556
rect 13692 6554 13748 6556
rect 13452 6502 13478 6554
rect 13478 6502 13508 6554
rect 13532 6502 13542 6554
rect 13542 6502 13588 6554
rect 13612 6502 13658 6554
rect 13658 6502 13668 6554
rect 13692 6502 13722 6554
rect 13722 6502 13748 6554
rect 13452 6500 13508 6502
rect 13532 6500 13588 6502
rect 13612 6500 13668 6502
rect 13692 6500 13748 6502
rect 10953 6010 11009 6012
rect 11033 6010 11089 6012
rect 11113 6010 11169 6012
rect 11193 6010 11249 6012
rect 10953 5958 10979 6010
rect 10979 5958 11009 6010
rect 11033 5958 11043 6010
rect 11043 5958 11089 6010
rect 11113 5958 11159 6010
rect 11159 5958 11169 6010
rect 11193 5958 11223 6010
rect 11223 5958 11249 6010
rect 10953 5956 11009 5958
rect 11033 5956 11089 5958
rect 11113 5956 11169 5958
rect 11193 5956 11249 5958
rect 8454 3290 8510 3292
rect 8534 3290 8590 3292
rect 8614 3290 8670 3292
rect 8694 3290 8750 3292
rect 8454 3238 8480 3290
rect 8480 3238 8510 3290
rect 8534 3238 8544 3290
rect 8544 3238 8590 3290
rect 8614 3238 8660 3290
rect 8660 3238 8670 3290
rect 8694 3238 8724 3290
rect 8724 3238 8750 3290
rect 8454 3236 8510 3238
rect 8534 3236 8590 3238
rect 8614 3236 8670 3238
rect 8694 3236 8750 3238
rect 10953 4922 11009 4924
rect 11033 4922 11089 4924
rect 11113 4922 11169 4924
rect 11193 4922 11249 4924
rect 10953 4870 10979 4922
rect 10979 4870 11009 4922
rect 11033 4870 11043 4922
rect 11043 4870 11089 4922
rect 11113 4870 11159 4922
rect 11159 4870 11169 4922
rect 11193 4870 11223 4922
rect 11223 4870 11249 4922
rect 10953 4868 11009 4870
rect 11033 4868 11089 4870
rect 11113 4868 11169 4870
rect 11193 4868 11249 4870
rect 13452 5466 13508 5468
rect 13532 5466 13588 5468
rect 13612 5466 13668 5468
rect 13692 5466 13748 5468
rect 13452 5414 13478 5466
rect 13478 5414 13508 5466
rect 13532 5414 13542 5466
rect 13542 5414 13588 5466
rect 13612 5414 13658 5466
rect 13658 5414 13668 5466
rect 13692 5414 13722 5466
rect 13722 5414 13748 5466
rect 13452 5412 13508 5414
rect 13532 5412 13588 5414
rect 13612 5412 13668 5414
rect 13692 5412 13748 5414
rect 10953 3834 11009 3836
rect 11033 3834 11089 3836
rect 11113 3834 11169 3836
rect 11193 3834 11249 3836
rect 10953 3782 10979 3834
rect 10979 3782 11009 3834
rect 11033 3782 11043 3834
rect 11043 3782 11089 3834
rect 11113 3782 11159 3834
rect 11159 3782 11169 3834
rect 11193 3782 11223 3834
rect 11223 3782 11249 3834
rect 10953 3780 11009 3782
rect 11033 3780 11089 3782
rect 11113 3780 11169 3782
rect 11193 3780 11249 3782
rect 10953 2746 11009 2748
rect 11033 2746 11089 2748
rect 11113 2746 11169 2748
rect 11193 2746 11249 2748
rect 10953 2694 10979 2746
rect 10979 2694 11009 2746
rect 11033 2694 11043 2746
rect 11043 2694 11089 2746
rect 11113 2694 11159 2746
rect 11159 2694 11169 2746
rect 11193 2694 11223 2746
rect 11223 2694 11249 2746
rect 10953 2692 11009 2694
rect 11033 2692 11089 2694
rect 11113 2692 11169 2694
rect 11193 2692 11249 2694
rect 13452 4378 13508 4380
rect 13532 4378 13588 4380
rect 13612 4378 13668 4380
rect 13692 4378 13748 4380
rect 13452 4326 13478 4378
rect 13478 4326 13508 4378
rect 13532 4326 13542 4378
rect 13542 4326 13588 4378
rect 13612 4326 13658 4378
rect 13658 4326 13668 4378
rect 13692 4326 13722 4378
rect 13722 4326 13748 4378
rect 13452 4324 13508 4326
rect 13532 4324 13588 4326
rect 13612 4324 13668 4326
rect 13692 4324 13748 4326
rect 13452 3290 13508 3292
rect 13532 3290 13588 3292
rect 13612 3290 13668 3292
rect 13692 3290 13748 3292
rect 13452 3238 13478 3290
rect 13478 3238 13508 3290
rect 13532 3238 13542 3290
rect 13542 3238 13588 3290
rect 13612 3238 13658 3290
rect 13658 3238 13668 3290
rect 13692 3238 13722 3290
rect 13722 3238 13748 3290
rect 13452 3236 13508 3238
rect 13532 3236 13588 3238
rect 13612 3236 13668 3238
rect 13692 3236 13748 3238
rect 3455 2202 3511 2204
rect 3535 2202 3591 2204
rect 3615 2202 3671 2204
rect 3695 2202 3751 2204
rect 3455 2150 3481 2202
rect 3481 2150 3511 2202
rect 3535 2150 3545 2202
rect 3545 2150 3591 2202
rect 3615 2150 3661 2202
rect 3661 2150 3671 2202
rect 3695 2150 3725 2202
rect 3725 2150 3751 2202
rect 3455 2148 3511 2150
rect 3535 2148 3591 2150
rect 3615 2148 3671 2150
rect 3695 2148 3751 2150
rect 8454 2202 8510 2204
rect 8534 2202 8590 2204
rect 8614 2202 8670 2204
rect 8694 2202 8750 2204
rect 8454 2150 8480 2202
rect 8480 2150 8510 2202
rect 8534 2150 8544 2202
rect 8544 2150 8590 2202
rect 8614 2150 8660 2202
rect 8660 2150 8670 2202
rect 8694 2150 8724 2202
rect 8724 2150 8750 2202
rect 8454 2148 8510 2150
rect 8534 2148 8590 2150
rect 8614 2148 8670 2150
rect 8694 2148 8750 2150
rect 13452 2202 13508 2204
rect 13532 2202 13588 2204
rect 13612 2202 13668 2204
rect 13692 2202 13748 2204
rect 13452 2150 13478 2202
rect 13478 2150 13508 2202
rect 13532 2150 13542 2202
rect 13542 2150 13588 2202
rect 13612 2150 13658 2202
rect 13658 2150 13668 2202
rect 13692 2150 13722 2202
rect 13722 2150 13748 2202
rect 13452 2148 13508 2150
rect 13532 2148 13588 2150
rect 13612 2148 13668 2150
rect 13692 2148 13748 2150
rect 15750 1400 15806 1456
<< metal3 >>
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 5942 16896 6262 16897
rect 5942 16832 5950 16896
rect 6014 16832 6030 16896
rect 6094 16832 6110 16896
rect 6174 16832 6190 16896
rect 6254 16832 6262 16896
rect 5942 16831 6262 16832
rect 10941 16896 11261 16897
rect 10941 16832 10949 16896
rect 11013 16832 11029 16896
rect 11093 16832 11109 16896
rect 11173 16832 11189 16896
rect 11253 16832 11261 16896
rect 10941 16831 11261 16832
rect 3443 16352 3763 16353
rect 3443 16288 3451 16352
rect 3515 16288 3531 16352
rect 3595 16288 3611 16352
rect 3675 16288 3691 16352
rect 3755 16288 3763 16352
rect 3443 16287 3763 16288
rect 8442 16352 8762 16353
rect 8442 16288 8450 16352
rect 8514 16288 8530 16352
rect 8594 16288 8610 16352
rect 8674 16288 8690 16352
rect 8754 16288 8762 16352
rect 8442 16287 8762 16288
rect 13440 16352 13760 16353
rect 13440 16288 13448 16352
rect 13512 16288 13528 16352
rect 13592 16288 13608 16352
rect 13672 16288 13688 16352
rect 13752 16288 13760 16352
rect 13440 16287 13760 16288
rect 5942 15808 6262 15809
rect 5942 15744 5950 15808
rect 6014 15744 6030 15808
rect 6094 15744 6110 15808
rect 6174 15744 6190 15808
rect 6254 15744 6262 15808
rect 5942 15743 6262 15744
rect 10941 15808 11261 15809
rect 10941 15744 10949 15808
rect 11013 15744 11029 15808
rect 11093 15744 11109 15808
rect 11173 15744 11189 15808
rect 11253 15744 11261 15808
rect 10941 15743 11261 15744
rect 3443 15264 3763 15265
rect 3443 15200 3451 15264
rect 3515 15200 3531 15264
rect 3595 15200 3611 15264
rect 3675 15200 3691 15264
rect 3755 15200 3763 15264
rect 3443 15199 3763 15200
rect 8442 15264 8762 15265
rect 8442 15200 8450 15264
rect 8514 15200 8530 15264
rect 8594 15200 8610 15264
rect 8674 15200 8690 15264
rect 8754 15200 8762 15264
rect 8442 15199 8762 15200
rect 13440 15264 13760 15265
rect 13440 15200 13448 15264
rect 13512 15200 13528 15264
rect 13592 15200 13608 15264
rect 13672 15200 13688 15264
rect 13752 15200 13760 15264
rect 13440 15199 13760 15200
rect 5942 14720 6262 14721
rect 5942 14656 5950 14720
rect 6014 14656 6030 14720
rect 6094 14656 6110 14720
rect 6174 14656 6190 14720
rect 6254 14656 6262 14720
rect 5942 14655 6262 14656
rect 10941 14720 11261 14721
rect 10941 14656 10949 14720
rect 11013 14656 11029 14720
rect 11093 14656 11109 14720
rect 11173 14656 11189 14720
rect 11253 14656 11261 14720
rect 10941 14655 11261 14656
rect 3443 14176 3763 14177
rect 3443 14112 3451 14176
rect 3515 14112 3531 14176
rect 3595 14112 3611 14176
rect 3675 14112 3691 14176
rect 3755 14112 3763 14176
rect 3443 14111 3763 14112
rect 8442 14176 8762 14177
rect 8442 14112 8450 14176
rect 8514 14112 8530 14176
rect 8594 14112 8610 14176
rect 8674 14112 8690 14176
rect 8754 14112 8762 14176
rect 8442 14111 8762 14112
rect 13440 14176 13760 14177
rect 13440 14112 13448 14176
rect 13512 14112 13528 14176
rect 13592 14112 13608 14176
rect 13672 14112 13688 14176
rect 13752 14112 13760 14176
rect 13440 14111 13760 14112
rect 9213 13834 9279 13837
rect 9949 13834 10015 13837
rect 9213 13832 10015 13834
rect 9213 13776 9218 13832
rect 9274 13776 9954 13832
rect 10010 13776 10015 13832
rect 9213 13774 10015 13776
rect 9213 13771 9279 13774
rect 9949 13771 10015 13774
rect 5942 13632 6262 13633
rect 5942 13568 5950 13632
rect 6014 13568 6030 13632
rect 6094 13568 6110 13632
rect 6174 13568 6190 13632
rect 6254 13568 6262 13632
rect 5942 13567 6262 13568
rect 10941 13632 11261 13633
rect 10941 13568 10949 13632
rect 11013 13568 11029 13632
rect 11093 13568 11109 13632
rect 11173 13568 11189 13632
rect 11253 13568 11261 13632
rect 10941 13567 11261 13568
rect 3443 13088 3763 13089
rect 3443 13024 3451 13088
rect 3515 13024 3531 13088
rect 3595 13024 3611 13088
rect 3675 13024 3691 13088
rect 3755 13024 3763 13088
rect 3443 13023 3763 13024
rect 8442 13088 8762 13089
rect 8442 13024 8450 13088
rect 8514 13024 8530 13088
rect 8594 13024 8610 13088
rect 8674 13024 8690 13088
rect 8754 13024 8762 13088
rect 8442 13023 8762 13024
rect 13440 13088 13760 13089
rect 13440 13024 13448 13088
rect 13512 13024 13528 13088
rect 13592 13024 13608 13088
rect 13672 13024 13688 13088
rect 13752 13024 13760 13088
rect 13440 13023 13760 13024
rect 5942 12544 6262 12545
rect 5942 12480 5950 12544
rect 6014 12480 6030 12544
rect 6094 12480 6110 12544
rect 6174 12480 6190 12544
rect 6254 12480 6262 12544
rect 5942 12479 6262 12480
rect 10941 12544 11261 12545
rect 10941 12480 10949 12544
rect 11013 12480 11029 12544
rect 11093 12480 11109 12544
rect 11173 12480 11189 12544
rect 11253 12480 11261 12544
rect 10941 12479 11261 12480
rect 8109 12202 8175 12205
rect 10225 12202 10291 12205
rect 8109 12200 10291 12202
rect 8109 12144 8114 12200
rect 8170 12144 10230 12200
rect 10286 12144 10291 12200
rect 8109 12142 10291 12144
rect 8109 12139 8175 12142
rect 10225 12139 10291 12142
rect 3443 12000 3763 12001
rect 3443 11936 3451 12000
rect 3515 11936 3531 12000
rect 3595 11936 3611 12000
rect 3675 11936 3691 12000
rect 3755 11936 3763 12000
rect 3443 11935 3763 11936
rect 8442 12000 8762 12001
rect 8442 11936 8450 12000
rect 8514 11936 8530 12000
rect 8594 11936 8610 12000
rect 8674 11936 8690 12000
rect 8754 11936 8762 12000
rect 8442 11935 8762 11936
rect 13440 12000 13760 12001
rect 13440 11936 13448 12000
rect 13512 11936 13528 12000
rect 13592 11936 13608 12000
rect 13672 11936 13688 12000
rect 13752 11936 13760 12000
rect 13440 11935 13760 11936
rect 7097 11794 7163 11797
rect 9581 11794 9647 11797
rect 7097 11792 9647 11794
rect 7097 11736 7102 11792
rect 7158 11736 9586 11792
rect 9642 11736 9647 11792
rect 7097 11734 9647 11736
rect 7097 11731 7163 11734
rect 9581 11731 9647 11734
rect 5942 11456 6262 11457
rect 5942 11392 5950 11456
rect 6014 11392 6030 11456
rect 6094 11392 6110 11456
rect 6174 11392 6190 11456
rect 6254 11392 6262 11456
rect 5942 11391 6262 11392
rect 10941 11456 11261 11457
rect 10941 11392 10949 11456
rect 11013 11392 11029 11456
rect 11093 11392 11109 11456
rect 11173 11392 11189 11456
rect 11253 11392 11261 11456
rect 10941 11391 11261 11392
rect 3443 10912 3763 10913
rect 3443 10848 3451 10912
rect 3515 10848 3531 10912
rect 3595 10848 3611 10912
rect 3675 10848 3691 10912
rect 3755 10848 3763 10912
rect 3443 10847 3763 10848
rect 8442 10912 8762 10913
rect 8442 10848 8450 10912
rect 8514 10848 8530 10912
rect 8594 10848 8610 10912
rect 8674 10848 8690 10912
rect 8754 10848 8762 10912
rect 8442 10847 8762 10848
rect 13440 10912 13760 10913
rect 13440 10848 13448 10912
rect 13512 10848 13528 10912
rect 13592 10848 13608 10912
rect 13672 10848 13688 10912
rect 13752 10848 13760 10912
rect 13440 10847 13760 10848
rect 5942 10368 6262 10369
rect 5942 10304 5950 10368
rect 6014 10304 6030 10368
rect 6094 10304 6110 10368
rect 6174 10304 6190 10368
rect 6254 10304 6262 10368
rect 5942 10303 6262 10304
rect 10941 10368 11261 10369
rect 10941 10304 10949 10368
rect 11013 10304 11029 10368
rect 11093 10304 11109 10368
rect 11173 10304 11189 10368
rect 11253 10304 11261 10368
rect 10941 10303 11261 10304
rect 15745 10298 15811 10301
rect 16446 10298 17246 10328
rect 15745 10296 17246 10298
rect 15745 10240 15750 10296
rect 15806 10240 17246 10296
rect 15745 10238 17246 10240
rect 15745 10235 15811 10238
rect 16446 10208 17246 10238
rect 9949 10162 10015 10165
rect 12525 10162 12591 10165
rect 9949 10160 12591 10162
rect 9949 10104 9954 10160
rect 10010 10104 12530 10160
rect 12586 10104 12591 10160
rect 9949 10102 12591 10104
rect 9949 10099 10015 10102
rect 12525 10099 12591 10102
rect 3443 9824 3763 9825
rect 3443 9760 3451 9824
rect 3515 9760 3531 9824
rect 3595 9760 3611 9824
rect 3675 9760 3691 9824
rect 3755 9760 3763 9824
rect 3443 9759 3763 9760
rect 8442 9824 8762 9825
rect 8442 9760 8450 9824
rect 8514 9760 8530 9824
rect 8594 9760 8610 9824
rect 8674 9760 8690 9824
rect 8754 9760 8762 9824
rect 8442 9759 8762 9760
rect 13440 9824 13760 9825
rect 13440 9760 13448 9824
rect 13512 9760 13528 9824
rect 13592 9760 13608 9824
rect 13672 9760 13688 9824
rect 13752 9760 13760 9824
rect 13440 9759 13760 9760
rect 5942 9280 6262 9281
rect 5942 9216 5950 9280
rect 6014 9216 6030 9280
rect 6094 9216 6110 9280
rect 6174 9216 6190 9280
rect 6254 9216 6262 9280
rect 5942 9215 6262 9216
rect 10941 9280 11261 9281
rect 10941 9216 10949 9280
rect 11013 9216 11029 9280
rect 11093 9216 11109 9280
rect 11173 9216 11189 9280
rect 11253 9216 11261 9280
rect 10941 9215 11261 9216
rect 0 8938 800 8968
rect 1393 8938 1459 8941
rect 0 8936 1459 8938
rect 0 8880 1398 8936
rect 1454 8880 1459 8936
rect 0 8878 1459 8880
rect 0 8848 800 8878
rect 1393 8875 1459 8878
rect 3443 8736 3763 8737
rect 3443 8672 3451 8736
rect 3515 8672 3531 8736
rect 3595 8672 3611 8736
rect 3675 8672 3691 8736
rect 3755 8672 3763 8736
rect 3443 8671 3763 8672
rect 8442 8736 8762 8737
rect 8442 8672 8450 8736
rect 8514 8672 8530 8736
rect 8594 8672 8610 8736
rect 8674 8672 8690 8736
rect 8754 8672 8762 8736
rect 8442 8671 8762 8672
rect 13440 8736 13760 8737
rect 13440 8672 13448 8736
rect 13512 8672 13528 8736
rect 13592 8672 13608 8736
rect 13672 8672 13688 8736
rect 13752 8672 13760 8736
rect 13440 8671 13760 8672
rect 5942 8192 6262 8193
rect 5942 8128 5950 8192
rect 6014 8128 6030 8192
rect 6094 8128 6110 8192
rect 6174 8128 6190 8192
rect 6254 8128 6262 8192
rect 5942 8127 6262 8128
rect 10941 8192 11261 8193
rect 10941 8128 10949 8192
rect 11013 8128 11029 8192
rect 11093 8128 11109 8192
rect 11173 8128 11189 8192
rect 11253 8128 11261 8192
rect 10941 8127 11261 8128
rect 3443 7648 3763 7649
rect 3443 7584 3451 7648
rect 3515 7584 3531 7648
rect 3595 7584 3611 7648
rect 3675 7584 3691 7648
rect 3755 7584 3763 7648
rect 3443 7583 3763 7584
rect 8442 7648 8762 7649
rect 8442 7584 8450 7648
rect 8514 7584 8530 7648
rect 8594 7584 8610 7648
rect 8674 7584 8690 7648
rect 8754 7584 8762 7648
rect 8442 7583 8762 7584
rect 13440 7648 13760 7649
rect 13440 7584 13448 7648
rect 13512 7584 13528 7648
rect 13592 7584 13608 7648
rect 13672 7584 13688 7648
rect 13752 7584 13760 7648
rect 13440 7583 13760 7584
rect 5942 7104 6262 7105
rect 5942 7040 5950 7104
rect 6014 7040 6030 7104
rect 6094 7040 6110 7104
rect 6174 7040 6190 7104
rect 6254 7040 6262 7104
rect 5942 7039 6262 7040
rect 10941 7104 11261 7105
rect 10941 7040 10949 7104
rect 11013 7040 11029 7104
rect 11093 7040 11109 7104
rect 11173 7040 11189 7104
rect 11253 7040 11261 7104
rect 10941 7039 11261 7040
rect 3443 6560 3763 6561
rect 3443 6496 3451 6560
rect 3515 6496 3531 6560
rect 3595 6496 3611 6560
rect 3675 6496 3691 6560
rect 3755 6496 3763 6560
rect 3443 6495 3763 6496
rect 8442 6560 8762 6561
rect 8442 6496 8450 6560
rect 8514 6496 8530 6560
rect 8594 6496 8610 6560
rect 8674 6496 8690 6560
rect 8754 6496 8762 6560
rect 8442 6495 8762 6496
rect 13440 6560 13760 6561
rect 13440 6496 13448 6560
rect 13512 6496 13528 6560
rect 13592 6496 13608 6560
rect 13672 6496 13688 6560
rect 13752 6496 13760 6560
rect 13440 6495 13760 6496
rect 5942 6016 6262 6017
rect 5942 5952 5950 6016
rect 6014 5952 6030 6016
rect 6094 5952 6110 6016
rect 6174 5952 6190 6016
rect 6254 5952 6262 6016
rect 5942 5951 6262 5952
rect 10941 6016 11261 6017
rect 10941 5952 10949 6016
rect 11013 5952 11029 6016
rect 11093 5952 11109 6016
rect 11173 5952 11189 6016
rect 11253 5952 11261 6016
rect 10941 5951 11261 5952
rect 3443 5472 3763 5473
rect 3443 5408 3451 5472
rect 3515 5408 3531 5472
rect 3595 5408 3611 5472
rect 3675 5408 3691 5472
rect 3755 5408 3763 5472
rect 3443 5407 3763 5408
rect 8442 5472 8762 5473
rect 8442 5408 8450 5472
rect 8514 5408 8530 5472
rect 8594 5408 8610 5472
rect 8674 5408 8690 5472
rect 8754 5408 8762 5472
rect 8442 5407 8762 5408
rect 13440 5472 13760 5473
rect 13440 5408 13448 5472
rect 13512 5408 13528 5472
rect 13592 5408 13608 5472
rect 13672 5408 13688 5472
rect 13752 5408 13760 5472
rect 13440 5407 13760 5408
rect 5942 4928 6262 4929
rect 5942 4864 5950 4928
rect 6014 4864 6030 4928
rect 6094 4864 6110 4928
rect 6174 4864 6190 4928
rect 6254 4864 6262 4928
rect 5942 4863 6262 4864
rect 10941 4928 11261 4929
rect 10941 4864 10949 4928
rect 11013 4864 11029 4928
rect 11093 4864 11109 4928
rect 11173 4864 11189 4928
rect 11253 4864 11261 4928
rect 10941 4863 11261 4864
rect 3443 4384 3763 4385
rect 3443 4320 3451 4384
rect 3515 4320 3531 4384
rect 3595 4320 3611 4384
rect 3675 4320 3691 4384
rect 3755 4320 3763 4384
rect 3443 4319 3763 4320
rect 8442 4384 8762 4385
rect 8442 4320 8450 4384
rect 8514 4320 8530 4384
rect 8594 4320 8610 4384
rect 8674 4320 8690 4384
rect 8754 4320 8762 4384
rect 8442 4319 8762 4320
rect 13440 4384 13760 4385
rect 13440 4320 13448 4384
rect 13512 4320 13528 4384
rect 13592 4320 13608 4384
rect 13672 4320 13688 4384
rect 13752 4320 13760 4384
rect 13440 4319 13760 4320
rect 5942 3840 6262 3841
rect 5942 3776 5950 3840
rect 6014 3776 6030 3840
rect 6094 3776 6110 3840
rect 6174 3776 6190 3840
rect 6254 3776 6262 3840
rect 5942 3775 6262 3776
rect 10941 3840 11261 3841
rect 10941 3776 10949 3840
rect 11013 3776 11029 3840
rect 11093 3776 11109 3840
rect 11173 3776 11189 3840
rect 11253 3776 11261 3840
rect 10941 3775 11261 3776
rect 3443 3296 3763 3297
rect 3443 3232 3451 3296
rect 3515 3232 3531 3296
rect 3595 3232 3611 3296
rect 3675 3232 3691 3296
rect 3755 3232 3763 3296
rect 3443 3231 3763 3232
rect 8442 3296 8762 3297
rect 8442 3232 8450 3296
rect 8514 3232 8530 3296
rect 8594 3232 8610 3296
rect 8674 3232 8690 3296
rect 8754 3232 8762 3296
rect 8442 3231 8762 3232
rect 13440 3296 13760 3297
rect 13440 3232 13448 3296
rect 13512 3232 13528 3296
rect 13592 3232 13608 3296
rect 13672 3232 13688 3296
rect 13752 3232 13760 3296
rect 13440 3231 13760 3232
rect 5942 2752 6262 2753
rect 5942 2688 5950 2752
rect 6014 2688 6030 2752
rect 6094 2688 6110 2752
rect 6174 2688 6190 2752
rect 6254 2688 6262 2752
rect 5942 2687 6262 2688
rect 10941 2752 11261 2753
rect 10941 2688 10949 2752
rect 11013 2688 11029 2752
rect 11093 2688 11109 2752
rect 11173 2688 11189 2752
rect 11253 2688 11261 2752
rect 10941 2687 11261 2688
rect 3443 2208 3763 2209
rect 3443 2144 3451 2208
rect 3515 2144 3531 2208
rect 3595 2144 3611 2208
rect 3675 2144 3691 2208
rect 3755 2144 3763 2208
rect 3443 2143 3763 2144
rect 8442 2208 8762 2209
rect 8442 2144 8450 2208
rect 8514 2144 8530 2208
rect 8594 2144 8610 2208
rect 8674 2144 8690 2208
rect 8754 2144 8762 2208
rect 8442 2143 8762 2144
rect 13440 2208 13760 2209
rect 13440 2144 13448 2208
rect 13512 2144 13528 2208
rect 13592 2144 13608 2208
rect 13672 2144 13688 2208
rect 13752 2144 13760 2208
rect 13440 2143 13760 2144
rect 15745 1458 15811 1461
rect 16446 1458 17246 1488
rect 15745 1456 17246 1458
rect 15745 1400 15750 1456
rect 15806 1400 17246 1456
rect 15745 1398 17246 1400
rect 15745 1395 15811 1398
rect 16446 1368 17246 1398
<< via3 >>
rect 5950 16892 6014 16896
rect 5950 16836 5954 16892
rect 5954 16836 6010 16892
rect 6010 16836 6014 16892
rect 5950 16832 6014 16836
rect 6030 16892 6094 16896
rect 6030 16836 6034 16892
rect 6034 16836 6090 16892
rect 6090 16836 6094 16892
rect 6030 16832 6094 16836
rect 6110 16892 6174 16896
rect 6110 16836 6114 16892
rect 6114 16836 6170 16892
rect 6170 16836 6174 16892
rect 6110 16832 6174 16836
rect 6190 16892 6254 16896
rect 6190 16836 6194 16892
rect 6194 16836 6250 16892
rect 6250 16836 6254 16892
rect 6190 16832 6254 16836
rect 10949 16892 11013 16896
rect 10949 16836 10953 16892
rect 10953 16836 11009 16892
rect 11009 16836 11013 16892
rect 10949 16832 11013 16836
rect 11029 16892 11093 16896
rect 11029 16836 11033 16892
rect 11033 16836 11089 16892
rect 11089 16836 11093 16892
rect 11029 16832 11093 16836
rect 11109 16892 11173 16896
rect 11109 16836 11113 16892
rect 11113 16836 11169 16892
rect 11169 16836 11173 16892
rect 11109 16832 11173 16836
rect 11189 16892 11253 16896
rect 11189 16836 11193 16892
rect 11193 16836 11249 16892
rect 11249 16836 11253 16892
rect 11189 16832 11253 16836
rect 3451 16348 3515 16352
rect 3451 16292 3455 16348
rect 3455 16292 3511 16348
rect 3511 16292 3515 16348
rect 3451 16288 3515 16292
rect 3531 16348 3595 16352
rect 3531 16292 3535 16348
rect 3535 16292 3591 16348
rect 3591 16292 3595 16348
rect 3531 16288 3595 16292
rect 3611 16348 3675 16352
rect 3611 16292 3615 16348
rect 3615 16292 3671 16348
rect 3671 16292 3675 16348
rect 3611 16288 3675 16292
rect 3691 16348 3755 16352
rect 3691 16292 3695 16348
rect 3695 16292 3751 16348
rect 3751 16292 3755 16348
rect 3691 16288 3755 16292
rect 8450 16348 8514 16352
rect 8450 16292 8454 16348
rect 8454 16292 8510 16348
rect 8510 16292 8514 16348
rect 8450 16288 8514 16292
rect 8530 16348 8594 16352
rect 8530 16292 8534 16348
rect 8534 16292 8590 16348
rect 8590 16292 8594 16348
rect 8530 16288 8594 16292
rect 8610 16348 8674 16352
rect 8610 16292 8614 16348
rect 8614 16292 8670 16348
rect 8670 16292 8674 16348
rect 8610 16288 8674 16292
rect 8690 16348 8754 16352
rect 8690 16292 8694 16348
rect 8694 16292 8750 16348
rect 8750 16292 8754 16348
rect 8690 16288 8754 16292
rect 13448 16348 13512 16352
rect 13448 16292 13452 16348
rect 13452 16292 13508 16348
rect 13508 16292 13512 16348
rect 13448 16288 13512 16292
rect 13528 16348 13592 16352
rect 13528 16292 13532 16348
rect 13532 16292 13588 16348
rect 13588 16292 13592 16348
rect 13528 16288 13592 16292
rect 13608 16348 13672 16352
rect 13608 16292 13612 16348
rect 13612 16292 13668 16348
rect 13668 16292 13672 16348
rect 13608 16288 13672 16292
rect 13688 16348 13752 16352
rect 13688 16292 13692 16348
rect 13692 16292 13748 16348
rect 13748 16292 13752 16348
rect 13688 16288 13752 16292
rect 5950 15804 6014 15808
rect 5950 15748 5954 15804
rect 5954 15748 6010 15804
rect 6010 15748 6014 15804
rect 5950 15744 6014 15748
rect 6030 15804 6094 15808
rect 6030 15748 6034 15804
rect 6034 15748 6090 15804
rect 6090 15748 6094 15804
rect 6030 15744 6094 15748
rect 6110 15804 6174 15808
rect 6110 15748 6114 15804
rect 6114 15748 6170 15804
rect 6170 15748 6174 15804
rect 6110 15744 6174 15748
rect 6190 15804 6254 15808
rect 6190 15748 6194 15804
rect 6194 15748 6250 15804
rect 6250 15748 6254 15804
rect 6190 15744 6254 15748
rect 10949 15804 11013 15808
rect 10949 15748 10953 15804
rect 10953 15748 11009 15804
rect 11009 15748 11013 15804
rect 10949 15744 11013 15748
rect 11029 15804 11093 15808
rect 11029 15748 11033 15804
rect 11033 15748 11089 15804
rect 11089 15748 11093 15804
rect 11029 15744 11093 15748
rect 11109 15804 11173 15808
rect 11109 15748 11113 15804
rect 11113 15748 11169 15804
rect 11169 15748 11173 15804
rect 11109 15744 11173 15748
rect 11189 15804 11253 15808
rect 11189 15748 11193 15804
rect 11193 15748 11249 15804
rect 11249 15748 11253 15804
rect 11189 15744 11253 15748
rect 3451 15260 3515 15264
rect 3451 15204 3455 15260
rect 3455 15204 3511 15260
rect 3511 15204 3515 15260
rect 3451 15200 3515 15204
rect 3531 15260 3595 15264
rect 3531 15204 3535 15260
rect 3535 15204 3591 15260
rect 3591 15204 3595 15260
rect 3531 15200 3595 15204
rect 3611 15260 3675 15264
rect 3611 15204 3615 15260
rect 3615 15204 3671 15260
rect 3671 15204 3675 15260
rect 3611 15200 3675 15204
rect 3691 15260 3755 15264
rect 3691 15204 3695 15260
rect 3695 15204 3751 15260
rect 3751 15204 3755 15260
rect 3691 15200 3755 15204
rect 8450 15260 8514 15264
rect 8450 15204 8454 15260
rect 8454 15204 8510 15260
rect 8510 15204 8514 15260
rect 8450 15200 8514 15204
rect 8530 15260 8594 15264
rect 8530 15204 8534 15260
rect 8534 15204 8590 15260
rect 8590 15204 8594 15260
rect 8530 15200 8594 15204
rect 8610 15260 8674 15264
rect 8610 15204 8614 15260
rect 8614 15204 8670 15260
rect 8670 15204 8674 15260
rect 8610 15200 8674 15204
rect 8690 15260 8754 15264
rect 8690 15204 8694 15260
rect 8694 15204 8750 15260
rect 8750 15204 8754 15260
rect 8690 15200 8754 15204
rect 13448 15260 13512 15264
rect 13448 15204 13452 15260
rect 13452 15204 13508 15260
rect 13508 15204 13512 15260
rect 13448 15200 13512 15204
rect 13528 15260 13592 15264
rect 13528 15204 13532 15260
rect 13532 15204 13588 15260
rect 13588 15204 13592 15260
rect 13528 15200 13592 15204
rect 13608 15260 13672 15264
rect 13608 15204 13612 15260
rect 13612 15204 13668 15260
rect 13668 15204 13672 15260
rect 13608 15200 13672 15204
rect 13688 15260 13752 15264
rect 13688 15204 13692 15260
rect 13692 15204 13748 15260
rect 13748 15204 13752 15260
rect 13688 15200 13752 15204
rect 5950 14716 6014 14720
rect 5950 14660 5954 14716
rect 5954 14660 6010 14716
rect 6010 14660 6014 14716
rect 5950 14656 6014 14660
rect 6030 14716 6094 14720
rect 6030 14660 6034 14716
rect 6034 14660 6090 14716
rect 6090 14660 6094 14716
rect 6030 14656 6094 14660
rect 6110 14716 6174 14720
rect 6110 14660 6114 14716
rect 6114 14660 6170 14716
rect 6170 14660 6174 14716
rect 6110 14656 6174 14660
rect 6190 14716 6254 14720
rect 6190 14660 6194 14716
rect 6194 14660 6250 14716
rect 6250 14660 6254 14716
rect 6190 14656 6254 14660
rect 10949 14716 11013 14720
rect 10949 14660 10953 14716
rect 10953 14660 11009 14716
rect 11009 14660 11013 14716
rect 10949 14656 11013 14660
rect 11029 14716 11093 14720
rect 11029 14660 11033 14716
rect 11033 14660 11089 14716
rect 11089 14660 11093 14716
rect 11029 14656 11093 14660
rect 11109 14716 11173 14720
rect 11109 14660 11113 14716
rect 11113 14660 11169 14716
rect 11169 14660 11173 14716
rect 11109 14656 11173 14660
rect 11189 14716 11253 14720
rect 11189 14660 11193 14716
rect 11193 14660 11249 14716
rect 11249 14660 11253 14716
rect 11189 14656 11253 14660
rect 3451 14172 3515 14176
rect 3451 14116 3455 14172
rect 3455 14116 3511 14172
rect 3511 14116 3515 14172
rect 3451 14112 3515 14116
rect 3531 14172 3595 14176
rect 3531 14116 3535 14172
rect 3535 14116 3591 14172
rect 3591 14116 3595 14172
rect 3531 14112 3595 14116
rect 3611 14172 3675 14176
rect 3611 14116 3615 14172
rect 3615 14116 3671 14172
rect 3671 14116 3675 14172
rect 3611 14112 3675 14116
rect 3691 14172 3755 14176
rect 3691 14116 3695 14172
rect 3695 14116 3751 14172
rect 3751 14116 3755 14172
rect 3691 14112 3755 14116
rect 8450 14172 8514 14176
rect 8450 14116 8454 14172
rect 8454 14116 8510 14172
rect 8510 14116 8514 14172
rect 8450 14112 8514 14116
rect 8530 14172 8594 14176
rect 8530 14116 8534 14172
rect 8534 14116 8590 14172
rect 8590 14116 8594 14172
rect 8530 14112 8594 14116
rect 8610 14172 8674 14176
rect 8610 14116 8614 14172
rect 8614 14116 8670 14172
rect 8670 14116 8674 14172
rect 8610 14112 8674 14116
rect 8690 14172 8754 14176
rect 8690 14116 8694 14172
rect 8694 14116 8750 14172
rect 8750 14116 8754 14172
rect 8690 14112 8754 14116
rect 13448 14172 13512 14176
rect 13448 14116 13452 14172
rect 13452 14116 13508 14172
rect 13508 14116 13512 14172
rect 13448 14112 13512 14116
rect 13528 14172 13592 14176
rect 13528 14116 13532 14172
rect 13532 14116 13588 14172
rect 13588 14116 13592 14172
rect 13528 14112 13592 14116
rect 13608 14172 13672 14176
rect 13608 14116 13612 14172
rect 13612 14116 13668 14172
rect 13668 14116 13672 14172
rect 13608 14112 13672 14116
rect 13688 14172 13752 14176
rect 13688 14116 13692 14172
rect 13692 14116 13748 14172
rect 13748 14116 13752 14172
rect 13688 14112 13752 14116
rect 5950 13628 6014 13632
rect 5950 13572 5954 13628
rect 5954 13572 6010 13628
rect 6010 13572 6014 13628
rect 5950 13568 6014 13572
rect 6030 13628 6094 13632
rect 6030 13572 6034 13628
rect 6034 13572 6090 13628
rect 6090 13572 6094 13628
rect 6030 13568 6094 13572
rect 6110 13628 6174 13632
rect 6110 13572 6114 13628
rect 6114 13572 6170 13628
rect 6170 13572 6174 13628
rect 6110 13568 6174 13572
rect 6190 13628 6254 13632
rect 6190 13572 6194 13628
rect 6194 13572 6250 13628
rect 6250 13572 6254 13628
rect 6190 13568 6254 13572
rect 10949 13628 11013 13632
rect 10949 13572 10953 13628
rect 10953 13572 11009 13628
rect 11009 13572 11013 13628
rect 10949 13568 11013 13572
rect 11029 13628 11093 13632
rect 11029 13572 11033 13628
rect 11033 13572 11089 13628
rect 11089 13572 11093 13628
rect 11029 13568 11093 13572
rect 11109 13628 11173 13632
rect 11109 13572 11113 13628
rect 11113 13572 11169 13628
rect 11169 13572 11173 13628
rect 11109 13568 11173 13572
rect 11189 13628 11253 13632
rect 11189 13572 11193 13628
rect 11193 13572 11249 13628
rect 11249 13572 11253 13628
rect 11189 13568 11253 13572
rect 3451 13084 3515 13088
rect 3451 13028 3455 13084
rect 3455 13028 3511 13084
rect 3511 13028 3515 13084
rect 3451 13024 3515 13028
rect 3531 13084 3595 13088
rect 3531 13028 3535 13084
rect 3535 13028 3591 13084
rect 3591 13028 3595 13084
rect 3531 13024 3595 13028
rect 3611 13084 3675 13088
rect 3611 13028 3615 13084
rect 3615 13028 3671 13084
rect 3671 13028 3675 13084
rect 3611 13024 3675 13028
rect 3691 13084 3755 13088
rect 3691 13028 3695 13084
rect 3695 13028 3751 13084
rect 3751 13028 3755 13084
rect 3691 13024 3755 13028
rect 8450 13084 8514 13088
rect 8450 13028 8454 13084
rect 8454 13028 8510 13084
rect 8510 13028 8514 13084
rect 8450 13024 8514 13028
rect 8530 13084 8594 13088
rect 8530 13028 8534 13084
rect 8534 13028 8590 13084
rect 8590 13028 8594 13084
rect 8530 13024 8594 13028
rect 8610 13084 8674 13088
rect 8610 13028 8614 13084
rect 8614 13028 8670 13084
rect 8670 13028 8674 13084
rect 8610 13024 8674 13028
rect 8690 13084 8754 13088
rect 8690 13028 8694 13084
rect 8694 13028 8750 13084
rect 8750 13028 8754 13084
rect 8690 13024 8754 13028
rect 13448 13084 13512 13088
rect 13448 13028 13452 13084
rect 13452 13028 13508 13084
rect 13508 13028 13512 13084
rect 13448 13024 13512 13028
rect 13528 13084 13592 13088
rect 13528 13028 13532 13084
rect 13532 13028 13588 13084
rect 13588 13028 13592 13084
rect 13528 13024 13592 13028
rect 13608 13084 13672 13088
rect 13608 13028 13612 13084
rect 13612 13028 13668 13084
rect 13668 13028 13672 13084
rect 13608 13024 13672 13028
rect 13688 13084 13752 13088
rect 13688 13028 13692 13084
rect 13692 13028 13748 13084
rect 13748 13028 13752 13084
rect 13688 13024 13752 13028
rect 5950 12540 6014 12544
rect 5950 12484 5954 12540
rect 5954 12484 6010 12540
rect 6010 12484 6014 12540
rect 5950 12480 6014 12484
rect 6030 12540 6094 12544
rect 6030 12484 6034 12540
rect 6034 12484 6090 12540
rect 6090 12484 6094 12540
rect 6030 12480 6094 12484
rect 6110 12540 6174 12544
rect 6110 12484 6114 12540
rect 6114 12484 6170 12540
rect 6170 12484 6174 12540
rect 6110 12480 6174 12484
rect 6190 12540 6254 12544
rect 6190 12484 6194 12540
rect 6194 12484 6250 12540
rect 6250 12484 6254 12540
rect 6190 12480 6254 12484
rect 10949 12540 11013 12544
rect 10949 12484 10953 12540
rect 10953 12484 11009 12540
rect 11009 12484 11013 12540
rect 10949 12480 11013 12484
rect 11029 12540 11093 12544
rect 11029 12484 11033 12540
rect 11033 12484 11089 12540
rect 11089 12484 11093 12540
rect 11029 12480 11093 12484
rect 11109 12540 11173 12544
rect 11109 12484 11113 12540
rect 11113 12484 11169 12540
rect 11169 12484 11173 12540
rect 11109 12480 11173 12484
rect 11189 12540 11253 12544
rect 11189 12484 11193 12540
rect 11193 12484 11249 12540
rect 11249 12484 11253 12540
rect 11189 12480 11253 12484
rect 3451 11996 3515 12000
rect 3451 11940 3455 11996
rect 3455 11940 3511 11996
rect 3511 11940 3515 11996
rect 3451 11936 3515 11940
rect 3531 11996 3595 12000
rect 3531 11940 3535 11996
rect 3535 11940 3591 11996
rect 3591 11940 3595 11996
rect 3531 11936 3595 11940
rect 3611 11996 3675 12000
rect 3611 11940 3615 11996
rect 3615 11940 3671 11996
rect 3671 11940 3675 11996
rect 3611 11936 3675 11940
rect 3691 11996 3755 12000
rect 3691 11940 3695 11996
rect 3695 11940 3751 11996
rect 3751 11940 3755 11996
rect 3691 11936 3755 11940
rect 8450 11996 8514 12000
rect 8450 11940 8454 11996
rect 8454 11940 8510 11996
rect 8510 11940 8514 11996
rect 8450 11936 8514 11940
rect 8530 11996 8594 12000
rect 8530 11940 8534 11996
rect 8534 11940 8590 11996
rect 8590 11940 8594 11996
rect 8530 11936 8594 11940
rect 8610 11996 8674 12000
rect 8610 11940 8614 11996
rect 8614 11940 8670 11996
rect 8670 11940 8674 11996
rect 8610 11936 8674 11940
rect 8690 11996 8754 12000
rect 8690 11940 8694 11996
rect 8694 11940 8750 11996
rect 8750 11940 8754 11996
rect 8690 11936 8754 11940
rect 13448 11996 13512 12000
rect 13448 11940 13452 11996
rect 13452 11940 13508 11996
rect 13508 11940 13512 11996
rect 13448 11936 13512 11940
rect 13528 11996 13592 12000
rect 13528 11940 13532 11996
rect 13532 11940 13588 11996
rect 13588 11940 13592 11996
rect 13528 11936 13592 11940
rect 13608 11996 13672 12000
rect 13608 11940 13612 11996
rect 13612 11940 13668 11996
rect 13668 11940 13672 11996
rect 13608 11936 13672 11940
rect 13688 11996 13752 12000
rect 13688 11940 13692 11996
rect 13692 11940 13748 11996
rect 13748 11940 13752 11996
rect 13688 11936 13752 11940
rect 5950 11452 6014 11456
rect 5950 11396 5954 11452
rect 5954 11396 6010 11452
rect 6010 11396 6014 11452
rect 5950 11392 6014 11396
rect 6030 11452 6094 11456
rect 6030 11396 6034 11452
rect 6034 11396 6090 11452
rect 6090 11396 6094 11452
rect 6030 11392 6094 11396
rect 6110 11452 6174 11456
rect 6110 11396 6114 11452
rect 6114 11396 6170 11452
rect 6170 11396 6174 11452
rect 6110 11392 6174 11396
rect 6190 11452 6254 11456
rect 6190 11396 6194 11452
rect 6194 11396 6250 11452
rect 6250 11396 6254 11452
rect 6190 11392 6254 11396
rect 10949 11452 11013 11456
rect 10949 11396 10953 11452
rect 10953 11396 11009 11452
rect 11009 11396 11013 11452
rect 10949 11392 11013 11396
rect 11029 11452 11093 11456
rect 11029 11396 11033 11452
rect 11033 11396 11089 11452
rect 11089 11396 11093 11452
rect 11029 11392 11093 11396
rect 11109 11452 11173 11456
rect 11109 11396 11113 11452
rect 11113 11396 11169 11452
rect 11169 11396 11173 11452
rect 11109 11392 11173 11396
rect 11189 11452 11253 11456
rect 11189 11396 11193 11452
rect 11193 11396 11249 11452
rect 11249 11396 11253 11452
rect 11189 11392 11253 11396
rect 3451 10908 3515 10912
rect 3451 10852 3455 10908
rect 3455 10852 3511 10908
rect 3511 10852 3515 10908
rect 3451 10848 3515 10852
rect 3531 10908 3595 10912
rect 3531 10852 3535 10908
rect 3535 10852 3591 10908
rect 3591 10852 3595 10908
rect 3531 10848 3595 10852
rect 3611 10908 3675 10912
rect 3611 10852 3615 10908
rect 3615 10852 3671 10908
rect 3671 10852 3675 10908
rect 3611 10848 3675 10852
rect 3691 10908 3755 10912
rect 3691 10852 3695 10908
rect 3695 10852 3751 10908
rect 3751 10852 3755 10908
rect 3691 10848 3755 10852
rect 8450 10908 8514 10912
rect 8450 10852 8454 10908
rect 8454 10852 8510 10908
rect 8510 10852 8514 10908
rect 8450 10848 8514 10852
rect 8530 10908 8594 10912
rect 8530 10852 8534 10908
rect 8534 10852 8590 10908
rect 8590 10852 8594 10908
rect 8530 10848 8594 10852
rect 8610 10908 8674 10912
rect 8610 10852 8614 10908
rect 8614 10852 8670 10908
rect 8670 10852 8674 10908
rect 8610 10848 8674 10852
rect 8690 10908 8754 10912
rect 8690 10852 8694 10908
rect 8694 10852 8750 10908
rect 8750 10852 8754 10908
rect 8690 10848 8754 10852
rect 13448 10908 13512 10912
rect 13448 10852 13452 10908
rect 13452 10852 13508 10908
rect 13508 10852 13512 10908
rect 13448 10848 13512 10852
rect 13528 10908 13592 10912
rect 13528 10852 13532 10908
rect 13532 10852 13588 10908
rect 13588 10852 13592 10908
rect 13528 10848 13592 10852
rect 13608 10908 13672 10912
rect 13608 10852 13612 10908
rect 13612 10852 13668 10908
rect 13668 10852 13672 10908
rect 13608 10848 13672 10852
rect 13688 10908 13752 10912
rect 13688 10852 13692 10908
rect 13692 10852 13748 10908
rect 13748 10852 13752 10908
rect 13688 10848 13752 10852
rect 5950 10364 6014 10368
rect 5950 10308 5954 10364
rect 5954 10308 6010 10364
rect 6010 10308 6014 10364
rect 5950 10304 6014 10308
rect 6030 10364 6094 10368
rect 6030 10308 6034 10364
rect 6034 10308 6090 10364
rect 6090 10308 6094 10364
rect 6030 10304 6094 10308
rect 6110 10364 6174 10368
rect 6110 10308 6114 10364
rect 6114 10308 6170 10364
rect 6170 10308 6174 10364
rect 6110 10304 6174 10308
rect 6190 10364 6254 10368
rect 6190 10308 6194 10364
rect 6194 10308 6250 10364
rect 6250 10308 6254 10364
rect 6190 10304 6254 10308
rect 10949 10364 11013 10368
rect 10949 10308 10953 10364
rect 10953 10308 11009 10364
rect 11009 10308 11013 10364
rect 10949 10304 11013 10308
rect 11029 10364 11093 10368
rect 11029 10308 11033 10364
rect 11033 10308 11089 10364
rect 11089 10308 11093 10364
rect 11029 10304 11093 10308
rect 11109 10364 11173 10368
rect 11109 10308 11113 10364
rect 11113 10308 11169 10364
rect 11169 10308 11173 10364
rect 11109 10304 11173 10308
rect 11189 10364 11253 10368
rect 11189 10308 11193 10364
rect 11193 10308 11249 10364
rect 11249 10308 11253 10364
rect 11189 10304 11253 10308
rect 3451 9820 3515 9824
rect 3451 9764 3455 9820
rect 3455 9764 3511 9820
rect 3511 9764 3515 9820
rect 3451 9760 3515 9764
rect 3531 9820 3595 9824
rect 3531 9764 3535 9820
rect 3535 9764 3591 9820
rect 3591 9764 3595 9820
rect 3531 9760 3595 9764
rect 3611 9820 3675 9824
rect 3611 9764 3615 9820
rect 3615 9764 3671 9820
rect 3671 9764 3675 9820
rect 3611 9760 3675 9764
rect 3691 9820 3755 9824
rect 3691 9764 3695 9820
rect 3695 9764 3751 9820
rect 3751 9764 3755 9820
rect 3691 9760 3755 9764
rect 8450 9820 8514 9824
rect 8450 9764 8454 9820
rect 8454 9764 8510 9820
rect 8510 9764 8514 9820
rect 8450 9760 8514 9764
rect 8530 9820 8594 9824
rect 8530 9764 8534 9820
rect 8534 9764 8590 9820
rect 8590 9764 8594 9820
rect 8530 9760 8594 9764
rect 8610 9820 8674 9824
rect 8610 9764 8614 9820
rect 8614 9764 8670 9820
rect 8670 9764 8674 9820
rect 8610 9760 8674 9764
rect 8690 9820 8754 9824
rect 8690 9764 8694 9820
rect 8694 9764 8750 9820
rect 8750 9764 8754 9820
rect 8690 9760 8754 9764
rect 13448 9820 13512 9824
rect 13448 9764 13452 9820
rect 13452 9764 13508 9820
rect 13508 9764 13512 9820
rect 13448 9760 13512 9764
rect 13528 9820 13592 9824
rect 13528 9764 13532 9820
rect 13532 9764 13588 9820
rect 13588 9764 13592 9820
rect 13528 9760 13592 9764
rect 13608 9820 13672 9824
rect 13608 9764 13612 9820
rect 13612 9764 13668 9820
rect 13668 9764 13672 9820
rect 13608 9760 13672 9764
rect 13688 9820 13752 9824
rect 13688 9764 13692 9820
rect 13692 9764 13748 9820
rect 13748 9764 13752 9820
rect 13688 9760 13752 9764
rect 5950 9276 6014 9280
rect 5950 9220 5954 9276
rect 5954 9220 6010 9276
rect 6010 9220 6014 9276
rect 5950 9216 6014 9220
rect 6030 9276 6094 9280
rect 6030 9220 6034 9276
rect 6034 9220 6090 9276
rect 6090 9220 6094 9276
rect 6030 9216 6094 9220
rect 6110 9276 6174 9280
rect 6110 9220 6114 9276
rect 6114 9220 6170 9276
rect 6170 9220 6174 9276
rect 6110 9216 6174 9220
rect 6190 9276 6254 9280
rect 6190 9220 6194 9276
rect 6194 9220 6250 9276
rect 6250 9220 6254 9276
rect 6190 9216 6254 9220
rect 10949 9276 11013 9280
rect 10949 9220 10953 9276
rect 10953 9220 11009 9276
rect 11009 9220 11013 9276
rect 10949 9216 11013 9220
rect 11029 9276 11093 9280
rect 11029 9220 11033 9276
rect 11033 9220 11089 9276
rect 11089 9220 11093 9276
rect 11029 9216 11093 9220
rect 11109 9276 11173 9280
rect 11109 9220 11113 9276
rect 11113 9220 11169 9276
rect 11169 9220 11173 9276
rect 11109 9216 11173 9220
rect 11189 9276 11253 9280
rect 11189 9220 11193 9276
rect 11193 9220 11249 9276
rect 11249 9220 11253 9276
rect 11189 9216 11253 9220
rect 3451 8732 3515 8736
rect 3451 8676 3455 8732
rect 3455 8676 3511 8732
rect 3511 8676 3515 8732
rect 3451 8672 3515 8676
rect 3531 8732 3595 8736
rect 3531 8676 3535 8732
rect 3535 8676 3591 8732
rect 3591 8676 3595 8732
rect 3531 8672 3595 8676
rect 3611 8732 3675 8736
rect 3611 8676 3615 8732
rect 3615 8676 3671 8732
rect 3671 8676 3675 8732
rect 3611 8672 3675 8676
rect 3691 8732 3755 8736
rect 3691 8676 3695 8732
rect 3695 8676 3751 8732
rect 3751 8676 3755 8732
rect 3691 8672 3755 8676
rect 8450 8732 8514 8736
rect 8450 8676 8454 8732
rect 8454 8676 8510 8732
rect 8510 8676 8514 8732
rect 8450 8672 8514 8676
rect 8530 8732 8594 8736
rect 8530 8676 8534 8732
rect 8534 8676 8590 8732
rect 8590 8676 8594 8732
rect 8530 8672 8594 8676
rect 8610 8732 8674 8736
rect 8610 8676 8614 8732
rect 8614 8676 8670 8732
rect 8670 8676 8674 8732
rect 8610 8672 8674 8676
rect 8690 8732 8754 8736
rect 8690 8676 8694 8732
rect 8694 8676 8750 8732
rect 8750 8676 8754 8732
rect 8690 8672 8754 8676
rect 13448 8732 13512 8736
rect 13448 8676 13452 8732
rect 13452 8676 13508 8732
rect 13508 8676 13512 8732
rect 13448 8672 13512 8676
rect 13528 8732 13592 8736
rect 13528 8676 13532 8732
rect 13532 8676 13588 8732
rect 13588 8676 13592 8732
rect 13528 8672 13592 8676
rect 13608 8732 13672 8736
rect 13608 8676 13612 8732
rect 13612 8676 13668 8732
rect 13668 8676 13672 8732
rect 13608 8672 13672 8676
rect 13688 8732 13752 8736
rect 13688 8676 13692 8732
rect 13692 8676 13748 8732
rect 13748 8676 13752 8732
rect 13688 8672 13752 8676
rect 5950 8188 6014 8192
rect 5950 8132 5954 8188
rect 5954 8132 6010 8188
rect 6010 8132 6014 8188
rect 5950 8128 6014 8132
rect 6030 8188 6094 8192
rect 6030 8132 6034 8188
rect 6034 8132 6090 8188
rect 6090 8132 6094 8188
rect 6030 8128 6094 8132
rect 6110 8188 6174 8192
rect 6110 8132 6114 8188
rect 6114 8132 6170 8188
rect 6170 8132 6174 8188
rect 6110 8128 6174 8132
rect 6190 8188 6254 8192
rect 6190 8132 6194 8188
rect 6194 8132 6250 8188
rect 6250 8132 6254 8188
rect 6190 8128 6254 8132
rect 10949 8188 11013 8192
rect 10949 8132 10953 8188
rect 10953 8132 11009 8188
rect 11009 8132 11013 8188
rect 10949 8128 11013 8132
rect 11029 8188 11093 8192
rect 11029 8132 11033 8188
rect 11033 8132 11089 8188
rect 11089 8132 11093 8188
rect 11029 8128 11093 8132
rect 11109 8188 11173 8192
rect 11109 8132 11113 8188
rect 11113 8132 11169 8188
rect 11169 8132 11173 8188
rect 11109 8128 11173 8132
rect 11189 8188 11253 8192
rect 11189 8132 11193 8188
rect 11193 8132 11249 8188
rect 11249 8132 11253 8188
rect 11189 8128 11253 8132
rect 3451 7644 3515 7648
rect 3451 7588 3455 7644
rect 3455 7588 3511 7644
rect 3511 7588 3515 7644
rect 3451 7584 3515 7588
rect 3531 7644 3595 7648
rect 3531 7588 3535 7644
rect 3535 7588 3591 7644
rect 3591 7588 3595 7644
rect 3531 7584 3595 7588
rect 3611 7644 3675 7648
rect 3611 7588 3615 7644
rect 3615 7588 3671 7644
rect 3671 7588 3675 7644
rect 3611 7584 3675 7588
rect 3691 7644 3755 7648
rect 3691 7588 3695 7644
rect 3695 7588 3751 7644
rect 3751 7588 3755 7644
rect 3691 7584 3755 7588
rect 8450 7644 8514 7648
rect 8450 7588 8454 7644
rect 8454 7588 8510 7644
rect 8510 7588 8514 7644
rect 8450 7584 8514 7588
rect 8530 7644 8594 7648
rect 8530 7588 8534 7644
rect 8534 7588 8590 7644
rect 8590 7588 8594 7644
rect 8530 7584 8594 7588
rect 8610 7644 8674 7648
rect 8610 7588 8614 7644
rect 8614 7588 8670 7644
rect 8670 7588 8674 7644
rect 8610 7584 8674 7588
rect 8690 7644 8754 7648
rect 8690 7588 8694 7644
rect 8694 7588 8750 7644
rect 8750 7588 8754 7644
rect 8690 7584 8754 7588
rect 13448 7644 13512 7648
rect 13448 7588 13452 7644
rect 13452 7588 13508 7644
rect 13508 7588 13512 7644
rect 13448 7584 13512 7588
rect 13528 7644 13592 7648
rect 13528 7588 13532 7644
rect 13532 7588 13588 7644
rect 13588 7588 13592 7644
rect 13528 7584 13592 7588
rect 13608 7644 13672 7648
rect 13608 7588 13612 7644
rect 13612 7588 13668 7644
rect 13668 7588 13672 7644
rect 13608 7584 13672 7588
rect 13688 7644 13752 7648
rect 13688 7588 13692 7644
rect 13692 7588 13748 7644
rect 13748 7588 13752 7644
rect 13688 7584 13752 7588
rect 5950 7100 6014 7104
rect 5950 7044 5954 7100
rect 5954 7044 6010 7100
rect 6010 7044 6014 7100
rect 5950 7040 6014 7044
rect 6030 7100 6094 7104
rect 6030 7044 6034 7100
rect 6034 7044 6090 7100
rect 6090 7044 6094 7100
rect 6030 7040 6094 7044
rect 6110 7100 6174 7104
rect 6110 7044 6114 7100
rect 6114 7044 6170 7100
rect 6170 7044 6174 7100
rect 6110 7040 6174 7044
rect 6190 7100 6254 7104
rect 6190 7044 6194 7100
rect 6194 7044 6250 7100
rect 6250 7044 6254 7100
rect 6190 7040 6254 7044
rect 10949 7100 11013 7104
rect 10949 7044 10953 7100
rect 10953 7044 11009 7100
rect 11009 7044 11013 7100
rect 10949 7040 11013 7044
rect 11029 7100 11093 7104
rect 11029 7044 11033 7100
rect 11033 7044 11089 7100
rect 11089 7044 11093 7100
rect 11029 7040 11093 7044
rect 11109 7100 11173 7104
rect 11109 7044 11113 7100
rect 11113 7044 11169 7100
rect 11169 7044 11173 7100
rect 11109 7040 11173 7044
rect 11189 7100 11253 7104
rect 11189 7044 11193 7100
rect 11193 7044 11249 7100
rect 11249 7044 11253 7100
rect 11189 7040 11253 7044
rect 3451 6556 3515 6560
rect 3451 6500 3455 6556
rect 3455 6500 3511 6556
rect 3511 6500 3515 6556
rect 3451 6496 3515 6500
rect 3531 6556 3595 6560
rect 3531 6500 3535 6556
rect 3535 6500 3591 6556
rect 3591 6500 3595 6556
rect 3531 6496 3595 6500
rect 3611 6556 3675 6560
rect 3611 6500 3615 6556
rect 3615 6500 3671 6556
rect 3671 6500 3675 6556
rect 3611 6496 3675 6500
rect 3691 6556 3755 6560
rect 3691 6500 3695 6556
rect 3695 6500 3751 6556
rect 3751 6500 3755 6556
rect 3691 6496 3755 6500
rect 8450 6556 8514 6560
rect 8450 6500 8454 6556
rect 8454 6500 8510 6556
rect 8510 6500 8514 6556
rect 8450 6496 8514 6500
rect 8530 6556 8594 6560
rect 8530 6500 8534 6556
rect 8534 6500 8590 6556
rect 8590 6500 8594 6556
rect 8530 6496 8594 6500
rect 8610 6556 8674 6560
rect 8610 6500 8614 6556
rect 8614 6500 8670 6556
rect 8670 6500 8674 6556
rect 8610 6496 8674 6500
rect 8690 6556 8754 6560
rect 8690 6500 8694 6556
rect 8694 6500 8750 6556
rect 8750 6500 8754 6556
rect 8690 6496 8754 6500
rect 13448 6556 13512 6560
rect 13448 6500 13452 6556
rect 13452 6500 13508 6556
rect 13508 6500 13512 6556
rect 13448 6496 13512 6500
rect 13528 6556 13592 6560
rect 13528 6500 13532 6556
rect 13532 6500 13588 6556
rect 13588 6500 13592 6556
rect 13528 6496 13592 6500
rect 13608 6556 13672 6560
rect 13608 6500 13612 6556
rect 13612 6500 13668 6556
rect 13668 6500 13672 6556
rect 13608 6496 13672 6500
rect 13688 6556 13752 6560
rect 13688 6500 13692 6556
rect 13692 6500 13748 6556
rect 13748 6500 13752 6556
rect 13688 6496 13752 6500
rect 5950 6012 6014 6016
rect 5950 5956 5954 6012
rect 5954 5956 6010 6012
rect 6010 5956 6014 6012
rect 5950 5952 6014 5956
rect 6030 6012 6094 6016
rect 6030 5956 6034 6012
rect 6034 5956 6090 6012
rect 6090 5956 6094 6012
rect 6030 5952 6094 5956
rect 6110 6012 6174 6016
rect 6110 5956 6114 6012
rect 6114 5956 6170 6012
rect 6170 5956 6174 6012
rect 6110 5952 6174 5956
rect 6190 6012 6254 6016
rect 6190 5956 6194 6012
rect 6194 5956 6250 6012
rect 6250 5956 6254 6012
rect 6190 5952 6254 5956
rect 10949 6012 11013 6016
rect 10949 5956 10953 6012
rect 10953 5956 11009 6012
rect 11009 5956 11013 6012
rect 10949 5952 11013 5956
rect 11029 6012 11093 6016
rect 11029 5956 11033 6012
rect 11033 5956 11089 6012
rect 11089 5956 11093 6012
rect 11029 5952 11093 5956
rect 11109 6012 11173 6016
rect 11109 5956 11113 6012
rect 11113 5956 11169 6012
rect 11169 5956 11173 6012
rect 11109 5952 11173 5956
rect 11189 6012 11253 6016
rect 11189 5956 11193 6012
rect 11193 5956 11249 6012
rect 11249 5956 11253 6012
rect 11189 5952 11253 5956
rect 3451 5468 3515 5472
rect 3451 5412 3455 5468
rect 3455 5412 3511 5468
rect 3511 5412 3515 5468
rect 3451 5408 3515 5412
rect 3531 5468 3595 5472
rect 3531 5412 3535 5468
rect 3535 5412 3591 5468
rect 3591 5412 3595 5468
rect 3531 5408 3595 5412
rect 3611 5468 3675 5472
rect 3611 5412 3615 5468
rect 3615 5412 3671 5468
rect 3671 5412 3675 5468
rect 3611 5408 3675 5412
rect 3691 5468 3755 5472
rect 3691 5412 3695 5468
rect 3695 5412 3751 5468
rect 3751 5412 3755 5468
rect 3691 5408 3755 5412
rect 8450 5468 8514 5472
rect 8450 5412 8454 5468
rect 8454 5412 8510 5468
rect 8510 5412 8514 5468
rect 8450 5408 8514 5412
rect 8530 5468 8594 5472
rect 8530 5412 8534 5468
rect 8534 5412 8590 5468
rect 8590 5412 8594 5468
rect 8530 5408 8594 5412
rect 8610 5468 8674 5472
rect 8610 5412 8614 5468
rect 8614 5412 8670 5468
rect 8670 5412 8674 5468
rect 8610 5408 8674 5412
rect 8690 5468 8754 5472
rect 8690 5412 8694 5468
rect 8694 5412 8750 5468
rect 8750 5412 8754 5468
rect 8690 5408 8754 5412
rect 13448 5468 13512 5472
rect 13448 5412 13452 5468
rect 13452 5412 13508 5468
rect 13508 5412 13512 5468
rect 13448 5408 13512 5412
rect 13528 5468 13592 5472
rect 13528 5412 13532 5468
rect 13532 5412 13588 5468
rect 13588 5412 13592 5468
rect 13528 5408 13592 5412
rect 13608 5468 13672 5472
rect 13608 5412 13612 5468
rect 13612 5412 13668 5468
rect 13668 5412 13672 5468
rect 13608 5408 13672 5412
rect 13688 5468 13752 5472
rect 13688 5412 13692 5468
rect 13692 5412 13748 5468
rect 13748 5412 13752 5468
rect 13688 5408 13752 5412
rect 5950 4924 6014 4928
rect 5950 4868 5954 4924
rect 5954 4868 6010 4924
rect 6010 4868 6014 4924
rect 5950 4864 6014 4868
rect 6030 4924 6094 4928
rect 6030 4868 6034 4924
rect 6034 4868 6090 4924
rect 6090 4868 6094 4924
rect 6030 4864 6094 4868
rect 6110 4924 6174 4928
rect 6110 4868 6114 4924
rect 6114 4868 6170 4924
rect 6170 4868 6174 4924
rect 6110 4864 6174 4868
rect 6190 4924 6254 4928
rect 6190 4868 6194 4924
rect 6194 4868 6250 4924
rect 6250 4868 6254 4924
rect 6190 4864 6254 4868
rect 10949 4924 11013 4928
rect 10949 4868 10953 4924
rect 10953 4868 11009 4924
rect 11009 4868 11013 4924
rect 10949 4864 11013 4868
rect 11029 4924 11093 4928
rect 11029 4868 11033 4924
rect 11033 4868 11089 4924
rect 11089 4868 11093 4924
rect 11029 4864 11093 4868
rect 11109 4924 11173 4928
rect 11109 4868 11113 4924
rect 11113 4868 11169 4924
rect 11169 4868 11173 4924
rect 11109 4864 11173 4868
rect 11189 4924 11253 4928
rect 11189 4868 11193 4924
rect 11193 4868 11249 4924
rect 11249 4868 11253 4924
rect 11189 4864 11253 4868
rect 3451 4380 3515 4384
rect 3451 4324 3455 4380
rect 3455 4324 3511 4380
rect 3511 4324 3515 4380
rect 3451 4320 3515 4324
rect 3531 4380 3595 4384
rect 3531 4324 3535 4380
rect 3535 4324 3591 4380
rect 3591 4324 3595 4380
rect 3531 4320 3595 4324
rect 3611 4380 3675 4384
rect 3611 4324 3615 4380
rect 3615 4324 3671 4380
rect 3671 4324 3675 4380
rect 3611 4320 3675 4324
rect 3691 4380 3755 4384
rect 3691 4324 3695 4380
rect 3695 4324 3751 4380
rect 3751 4324 3755 4380
rect 3691 4320 3755 4324
rect 8450 4380 8514 4384
rect 8450 4324 8454 4380
rect 8454 4324 8510 4380
rect 8510 4324 8514 4380
rect 8450 4320 8514 4324
rect 8530 4380 8594 4384
rect 8530 4324 8534 4380
rect 8534 4324 8590 4380
rect 8590 4324 8594 4380
rect 8530 4320 8594 4324
rect 8610 4380 8674 4384
rect 8610 4324 8614 4380
rect 8614 4324 8670 4380
rect 8670 4324 8674 4380
rect 8610 4320 8674 4324
rect 8690 4380 8754 4384
rect 8690 4324 8694 4380
rect 8694 4324 8750 4380
rect 8750 4324 8754 4380
rect 8690 4320 8754 4324
rect 13448 4380 13512 4384
rect 13448 4324 13452 4380
rect 13452 4324 13508 4380
rect 13508 4324 13512 4380
rect 13448 4320 13512 4324
rect 13528 4380 13592 4384
rect 13528 4324 13532 4380
rect 13532 4324 13588 4380
rect 13588 4324 13592 4380
rect 13528 4320 13592 4324
rect 13608 4380 13672 4384
rect 13608 4324 13612 4380
rect 13612 4324 13668 4380
rect 13668 4324 13672 4380
rect 13608 4320 13672 4324
rect 13688 4380 13752 4384
rect 13688 4324 13692 4380
rect 13692 4324 13748 4380
rect 13748 4324 13752 4380
rect 13688 4320 13752 4324
rect 5950 3836 6014 3840
rect 5950 3780 5954 3836
rect 5954 3780 6010 3836
rect 6010 3780 6014 3836
rect 5950 3776 6014 3780
rect 6030 3836 6094 3840
rect 6030 3780 6034 3836
rect 6034 3780 6090 3836
rect 6090 3780 6094 3836
rect 6030 3776 6094 3780
rect 6110 3836 6174 3840
rect 6110 3780 6114 3836
rect 6114 3780 6170 3836
rect 6170 3780 6174 3836
rect 6110 3776 6174 3780
rect 6190 3836 6254 3840
rect 6190 3780 6194 3836
rect 6194 3780 6250 3836
rect 6250 3780 6254 3836
rect 6190 3776 6254 3780
rect 10949 3836 11013 3840
rect 10949 3780 10953 3836
rect 10953 3780 11009 3836
rect 11009 3780 11013 3836
rect 10949 3776 11013 3780
rect 11029 3836 11093 3840
rect 11029 3780 11033 3836
rect 11033 3780 11089 3836
rect 11089 3780 11093 3836
rect 11029 3776 11093 3780
rect 11109 3836 11173 3840
rect 11109 3780 11113 3836
rect 11113 3780 11169 3836
rect 11169 3780 11173 3836
rect 11109 3776 11173 3780
rect 11189 3836 11253 3840
rect 11189 3780 11193 3836
rect 11193 3780 11249 3836
rect 11249 3780 11253 3836
rect 11189 3776 11253 3780
rect 3451 3292 3515 3296
rect 3451 3236 3455 3292
rect 3455 3236 3511 3292
rect 3511 3236 3515 3292
rect 3451 3232 3515 3236
rect 3531 3292 3595 3296
rect 3531 3236 3535 3292
rect 3535 3236 3591 3292
rect 3591 3236 3595 3292
rect 3531 3232 3595 3236
rect 3611 3292 3675 3296
rect 3611 3236 3615 3292
rect 3615 3236 3671 3292
rect 3671 3236 3675 3292
rect 3611 3232 3675 3236
rect 3691 3292 3755 3296
rect 3691 3236 3695 3292
rect 3695 3236 3751 3292
rect 3751 3236 3755 3292
rect 3691 3232 3755 3236
rect 8450 3292 8514 3296
rect 8450 3236 8454 3292
rect 8454 3236 8510 3292
rect 8510 3236 8514 3292
rect 8450 3232 8514 3236
rect 8530 3292 8594 3296
rect 8530 3236 8534 3292
rect 8534 3236 8590 3292
rect 8590 3236 8594 3292
rect 8530 3232 8594 3236
rect 8610 3292 8674 3296
rect 8610 3236 8614 3292
rect 8614 3236 8670 3292
rect 8670 3236 8674 3292
rect 8610 3232 8674 3236
rect 8690 3292 8754 3296
rect 8690 3236 8694 3292
rect 8694 3236 8750 3292
rect 8750 3236 8754 3292
rect 8690 3232 8754 3236
rect 13448 3292 13512 3296
rect 13448 3236 13452 3292
rect 13452 3236 13508 3292
rect 13508 3236 13512 3292
rect 13448 3232 13512 3236
rect 13528 3292 13592 3296
rect 13528 3236 13532 3292
rect 13532 3236 13588 3292
rect 13588 3236 13592 3292
rect 13528 3232 13592 3236
rect 13608 3292 13672 3296
rect 13608 3236 13612 3292
rect 13612 3236 13668 3292
rect 13668 3236 13672 3292
rect 13608 3232 13672 3236
rect 13688 3292 13752 3296
rect 13688 3236 13692 3292
rect 13692 3236 13748 3292
rect 13748 3236 13752 3292
rect 13688 3232 13752 3236
rect 5950 2748 6014 2752
rect 5950 2692 5954 2748
rect 5954 2692 6010 2748
rect 6010 2692 6014 2748
rect 5950 2688 6014 2692
rect 6030 2748 6094 2752
rect 6030 2692 6034 2748
rect 6034 2692 6090 2748
rect 6090 2692 6094 2748
rect 6030 2688 6094 2692
rect 6110 2748 6174 2752
rect 6110 2692 6114 2748
rect 6114 2692 6170 2748
rect 6170 2692 6174 2748
rect 6110 2688 6174 2692
rect 6190 2748 6254 2752
rect 6190 2692 6194 2748
rect 6194 2692 6250 2748
rect 6250 2692 6254 2748
rect 6190 2688 6254 2692
rect 10949 2748 11013 2752
rect 10949 2692 10953 2748
rect 10953 2692 11009 2748
rect 11009 2692 11013 2748
rect 10949 2688 11013 2692
rect 11029 2748 11093 2752
rect 11029 2692 11033 2748
rect 11033 2692 11089 2748
rect 11089 2692 11093 2748
rect 11029 2688 11093 2692
rect 11109 2748 11173 2752
rect 11109 2692 11113 2748
rect 11113 2692 11169 2748
rect 11169 2692 11173 2748
rect 11109 2688 11173 2692
rect 11189 2748 11253 2752
rect 11189 2692 11193 2748
rect 11193 2692 11249 2748
rect 11249 2692 11253 2748
rect 11189 2688 11253 2692
rect 3451 2204 3515 2208
rect 3451 2148 3455 2204
rect 3455 2148 3511 2204
rect 3511 2148 3515 2204
rect 3451 2144 3515 2148
rect 3531 2204 3595 2208
rect 3531 2148 3535 2204
rect 3535 2148 3591 2204
rect 3591 2148 3595 2204
rect 3531 2144 3595 2148
rect 3611 2204 3675 2208
rect 3611 2148 3615 2204
rect 3615 2148 3671 2204
rect 3671 2148 3675 2204
rect 3611 2144 3675 2148
rect 3691 2204 3755 2208
rect 3691 2148 3695 2204
rect 3695 2148 3751 2204
rect 3751 2148 3755 2204
rect 3691 2144 3755 2148
rect 8450 2204 8514 2208
rect 8450 2148 8454 2204
rect 8454 2148 8510 2204
rect 8510 2148 8514 2204
rect 8450 2144 8514 2148
rect 8530 2204 8594 2208
rect 8530 2148 8534 2204
rect 8534 2148 8590 2204
rect 8590 2148 8594 2204
rect 8530 2144 8594 2148
rect 8610 2204 8674 2208
rect 8610 2148 8614 2204
rect 8614 2148 8670 2204
rect 8670 2148 8674 2204
rect 8610 2144 8674 2148
rect 8690 2204 8754 2208
rect 8690 2148 8694 2204
rect 8694 2148 8750 2204
rect 8750 2148 8754 2204
rect 8690 2144 8754 2148
rect 13448 2204 13512 2208
rect 13448 2148 13452 2204
rect 13452 2148 13508 2204
rect 13508 2148 13512 2204
rect 13448 2144 13512 2148
rect 13528 2204 13592 2208
rect 13528 2148 13532 2204
rect 13532 2148 13588 2204
rect 13588 2148 13592 2204
rect 13528 2144 13592 2148
rect 13608 2204 13672 2208
rect 13608 2148 13612 2204
rect 13612 2148 13668 2204
rect 13668 2148 13672 2204
rect 13608 2144 13672 2148
rect 13688 2204 13752 2208
rect 13688 2148 13692 2204
rect 13692 2148 13748 2204
rect 13748 2148 13752 2204
rect 13688 2144 13752 2148
<< metal4 >>
rect 3443 16352 3763 16912
rect 3443 16288 3451 16352
rect 3515 16288 3531 16352
rect 3595 16288 3611 16352
rect 3675 16288 3691 16352
rect 3755 16288 3763 16352
rect 3443 15264 3763 16288
rect 3443 15200 3451 15264
rect 3515 15200 3531 15264
rect 3595 15200 3611 15264
rect 3675 15200 3691 15264
rect 3755 15200 3763 15264
rect 3443 14486 3763 15200
rect 3443 14250 3485 14486
rect 3721 14250 3763 14486
rect 3443 14176 3763 14250
rect 3443 14112 3451 14176
rect 3515 14112 3531 14176
rect 3595 14112 3611 14176
rect 3675 14112 3691 14176
rect 3755 14112 3763 14176
rect 3443 13088 3763 14112
rect 3443 13024 3451 13088
rect 3515 13024 3531 13088
rect 3595 13024 3611 13088
rect 3675 13024 3691 13088
rect 3755 13024 3763 13088
rect 3443 12000 3763 13024
rect 3443 11936 3451 12000
rect 3515 11936 3531 12000
rect 3595 11936 3611 12000
rect 3675 11936 3691 12000
rect 3755 11936 3763 12000
rect 3443 10912 3763 11936
rect 3443 10848 3451 10912
rect 3515 10848 3531 10912
rect 3595 10848 3611 10912
rect 3675 10848 3691 10912
rect 3755 10848 3763 10912
rect 3443 9824 3763 10848
rect 3443 9760 3451 9824
rect 3515 9760 3531 9824
rect 3595 9760 3611 9824
rect 3675 9760 3691 9824
rect 3755 9760 3763 9824
rect 3443 9590 3763 9760
rect 3443 9354 3485 9590
rect 3721 9354 3763 9590
rect 3443 8736 3763 9354
rect 3443 8672 3451 8736
rect 3515 8672 3531 8736
rect 3595 8672 3611 8736
rect 3675 8672 3691 8736
rect 3755 8672 3763 8736
rect 3443 7648 3763 8672
rect 3443 7584 3451 7648
rect 3515 7584 3531 7648
rect 3595 7584 3611 7648
rect 3675 7584 3691 7648
rect 3755 7584 3763 7648
rect 3443 6560 3763 7584
rect 3443 6496 3451 6560
rect 3515 6496 3531 6560
rect 3595 6496 3611 6560
rect 3675 6496 3691 6560
rect 3755 6496 3763 6560
rect 3443 5472 3763 6496
rect 3443 5408 3451 5472
rect 3515 5408 3531 5472
rect 3595 5408 3611 5472
rect 3675 5408 3691 5472
rect 3755 5408 3763 5472
rect 3443 4694 3763 5408
rect 3443 4458 3485 4694
rect 3721 4458 3763 4694
rect 3443 4384 3763 4458
rect 3443 4320 3451 4384
rect 3515 4320 3531 4384
rect 3595 4320 3611 4384
rect 3675 4320 3691 4384
rect 3755 4320 3763 4384
rect 3443 3296 3763 4320
rect 3443 3232 3451 3296
rect 3515 3232 3531 3296
rect 3595 3232 3611 3296
rect 3675 3232 3691 3296
rect 3755 3232 3763 3296
rect 3443 2208 3763 3232
rect 3443 2144 3451 2208
rect 3515 2144 3531 2208
rect 3595 2144 3611 2208
rect 3675 2144 3691 2208
rect 3755 2144 3763 2208
rect 3443 2128 3763 2144
rect 5942 16896 6263 16912
rect 5942 16832 5950 16896
rect 6014 16832 6030 16896
rect 6094 16832 6110 16896
rect 6174 16832 6190 16896
rect 6254 16832 6263 16896
rect 5942 15808 6263 16832
rect 5942 15744 5950 15808
rect 6014 15744 6030 15808
rect 6094 15744 6110 15808
rect 6174 15744 6190 15808
rect 6254 15744 6263 15808
rect 5942 14720 6263 15744
rect 5942 14656 5950 14720
rect 6014 14656 6030 14720
rect 6094 14656 6110 14720
rect 6174 14656 6190 14720
rect 6254 14656 6263 14720
rect 5942 13632 6263 14656
rect 5942 13568 5950 13632
rect 6014 13568 6030 13632
rect 6094 13568 6110 13632
rect 6174 13568 6190 13632
rect 6254 13568 6263 13632
rect 5942 12544 6263 13568
rect 5942 12480 5950 12544
rect 6014 12480 6030 12544
rect 6094 12480 6110 12544
rect 6174 12480 6190 12544
rect 6254 12480 6263 12544
rect 5942 12038 6263 12480
rect 5942 11802 5984 12038
rect 6220 11802 6263 12038
rect 5942 11456 6263 11802
rect 5942 11392 5950 11456
rect 6014 11392 6030 11456
rect 6094 11392 6110 11456
rect 6174 11392 6190 11456
rect 6254 11392 6263 11456
rect 5942 10368 6263 11392
rect 5942 10304 5950 10368
rect 6014 10304 6030 10368
rect 6094 10304 6110 10368
rect 6174 10304 6190 10368
rect 6254 10304 6263 10368
rect 5942 9280 6263 10304
rect 5942 9216 5950 9280
rect 6014 9216 6030 9280
rect 6094 9216 6110 9280
rect 6174 9216 6190 9280
rect 6254 9216 6263 9280
rect 5942 8192 6263 9216
rect 5942 8128 5950 8192
rect 6014 8128 6030 8192
rect 6094 8128 6110 8192
rect 6174 8128 6190 8192
rect 6254 8128 6263 8192
rect 5942 7142 6263 8128
rect 5942 7104 5984 7142
rect 6220 7104 6263 7142
rect 5942 7040 5950 7104
rect 6254 7040 6263 7104
rect 5942 6906 5984 7040
rect 6220 6906 6263 7040
rect 5942 6016 6263 6906
rect 5942 5952 5950 6016
rect 6014 5952 6030 6016
rect 6094 5952 6110 6016
rect 6174 5952 6190 6016
rect 6254 5952 6263 6016
rect 5942 4928 6263 5952
rect 5942 4864 5950 4928
rect 6014 4864 6030 4928
rect 6094 4864 6110 4928
rect 6174 4864 6190 4928
rect 6254 4864 6263 4928
rect 5942 3840 6263 4864
rect 5942 3776 5950 3840
rect 6014 3776 6030 3840
rect 6094 3776 6110 3840
rect 6174 3776 6190 3840
rect 6254 3776 6263 3840
rect 5942 2752 6263 3776
rect 5942 2688 5950 2752
rect 6014 2688 6030 2752
rect 6094 2688 6110 2752
rect 6174 2688 6190 2752
rect 6254 2688 6263 2752
rect 5942 2128 6263 2688
rect 8442 16352 8762 16912
rect 8442 16288 8450 16352
rect 8514 16288 8530 16352
rect 8594 16288 8610 16352
rect 8674 16288 8690 16352
rect 8754 16288 8762 16352
rect 8442 15264 8762 16288
rect 8442 15200 8450 15264
rect 8514 15200 8530 15264
rect 8594 15200 8610 15264
rect 8674 15200 8690 15264
rect 8754 15200 8762 15264
rect 8442 14486 8762 15200
rect 8442 14250 8484 14486
rect 8720 14250 8762 14486
rect 8442 14176 8762 14250
rect 8442 14112 8450 14176
rect 8514 14112 8530 14176
rect 8594 14112 8610 14176
rect 8674 14112 8690 14176
rect 8754 14112 8762 14176
rect 8442 13088 8762 14112
rect 8442 13024 8450 13088
rect 8514 13024 8530 13088
rect 8594 13024 8610 13088
rect 8674 13024 8690 13088
rect 8754 13024 8762 13088
rect 8442 12000 8762 13024
rect 8442 11936 8450 12000
rect 8514 11936 8530 12000
rect 8594 11936 8610 12000
rect 8674 11936 8690 12000
rect 8754 11936 8762 12000
rect 8442 10912 8762 11936
rect 8442 10848 8450 10912
rect 8514 10848 8530 10912
rect 8594 10848 8610 10912
rect 8674 10848 8690 10912
rect 8754 10848 8762 10912
rect 8442 9824 8762 10848
rect 8442 9760 8450 9824
rect 8514 9760 8530 9824
rect 8594 9760 8610 9824
rect 8674 9760 8690 9824
rect 8754 9760 8762 9824
rect 8442 9590 8762 9760
rect 8442 9354 8484 9590
rect 8720 9354 8762 9590
rect 8442 8736 8762 9354
rect 8442 8672 8450 8736
rect 8514 8672 8530 8736
rect 8594 8672 8610 8736
rect 8674 8672 8690 8736
rect 8754 8672 8762 8736
rect 8442 7648 8762 8672
rect 8442 7584 8450 7648
rect 8514 7584 8530 7648
rect 8594 7584 8610 7648
rect 8674 7584 8690 7648
rect 8754 7584 8762 7648
rect 8442 6560 8762 7584
rect 8442 6496 8450 6560
rect 8514 6496 8530 6560
rect 8594 6496 8610 6560
rect 8674 6496 8690 6560
rect 8754 6496 8762 6560
rect 8442 5472 8762 6496
rect 8442 5408 8450 5472
rect 8514 5408 8530 5472
rect 8594 5408 8610 5472
rect 8674 5408 8690 5472
rect 8754 5408 8762 5472
rect 8442 4694 8762 5408
rect 8442 4458 8484 4694
rect 8720 4458 8762 4694
rect 8442 4384 8762 4458
rect 8442 4320 8450 4384
rect 8514 4320 8530 4384
rect 8594 4320 8610 4384
rect 8674 4320 8690 4384
rect 8754 4320 8762 4384
rect 8442 3296 8762 4320
rect 8442 3232 8450 3296
rect 8514 3232 8530 3296
rect 8594 3232 8610 3296
rect 8674 3232 8690 3296
rect 8754 3232 8762 3296
rect 8442 2208 8762 3232
rect 8442 2144 8450 2208
rect 8514 2144 8530 2208
rect 8594 2144 8610 2208
rect 8674 2144 8690 2208
rect 8754 2144 8762 2208
rect 8442 2128 8762 2144
rect 10941 16896 11261 16912
rect 10941 16832 10949 16896
rect 11013 16832 11029 16896
rect 11093 16832 11109 16896
rect 11173 16832 11189 16896
rect 11253 16832 11261 16896
rect 10941 15808 11261 16832
rect 10941 15744 10949 15808
rect 11013 15744 11029 15808
rect 11093 15744 11109 15808
rect 11173 15744 11189 15808
rect 11253 15744 11261 15808
rect 10941 14720 11261 15744
rect 10941 14656 10949 14720
rect 11013 14656 11029 14720
rect 11093 14656 11109 14720
rect 11173 14656 11189 14720
rect 11253 14656 11261 14720
rect 10941 13632 11261 14656
rect 10941 13568 10949 13632
rect 11013 13568 11029 13632
rect 11093 13568 11109 13632
rect 11173 13568 11189 13632
rect 11253 13568 11261 13632
rect 10941 12544 11261 13568
rect 10941 12480 10949 12544
rect 11013 12480 11029 12544
rect 11093 12480 11109 12544
rect 11173 12480 11189 12544
rect 11253 12480 11261 12544
rect 10941 12038 11261 12480
rect 10941 11802 10983 12038
rect 11219 11802 11261 12038
rect 10941 11456 11261 11802
rect 10941 11392 10949 11456
rect 11013 11392 11029 11456
rect 11093 11392 11109 11456
rect 11173 11392 11189 11456
rect 11253 11392 11261 11456
rect 10941 10368 11261 11392
rect 10941 10304 10949 10368
rect 11013 10304 11029 10368
rect 11093 10304 11109 10368
rect 11173 10304 11189 10368
rect 11253 10304 11261 10368
rect 10941 9280 11261 10304
rect 10941 9216 10949 9280
rect 11013 9216 11029 9280
rect 11093 9216 11109 9280
rect 11173 9216 11189 9280
rect 11253 9216 11261 9280
rect 10941 8192 11261 9216
rect 10941 8128 10949 8192
rect 11013 8128 11029 8192
rect 11093 8128 11109 8192
rect 11173 8128 11189 8192
rect 11253 8128 11261 8192
rect 10941 7142 11261 8128
rect 10941 7104 10983 7142
rect 11219 7104 11261 7142
rect 10941 7040 10949 7104
rect 11253 7040 11261 7104
rect 10941 6906 10983 7040
rect 11219 6906 11261 7040
rect 10941 6016 11261 6906
rect 10941 5952 10949 6016
rect 11013 5952 11029 6016
rect 11093 5952 11109 6016
rect 11173 5952 11189 6016
rect 11253 5952 11261 6016
rect 10941 4928 11261 5952
rect 10941 4864 10949 4928
rect 11013 4864 11029 4928
rect 11093 4864 11109 4928
rect 11173 4864 11189 4928
rect 11253 4864 11261 4928
rect 10941 3840 11261 4864
rect 10941 3776 10949 3840
rect 11013 3776 11029 3840
rect 11093 3776 11109 3840
rect 11173 3776 11189 3840
rect 11253 3776 11261 3840
rect 10941 2752 11261 3776
rect 10941 2688 10949 2752
rect 11013 2688 11029 2752
rect 11093 2688 11109 2752
rect 11173 2688 11189 2752
rect 11253 2688 11261 2752
rect 10941 2128 11261 2688
rect 13440 16352 13761 16912
rect 13440 16288 13448 16352
rect 13512 16288 13528 16352
rect 13592 16288 13608 16352
rect 13672 16288 13688 16352
rect 13752 16288 13761 16352
rect 13440 15264 13761 16288
rect 13440 15200 13448 15264
rect 13512 15200 13528 15264
rect 13592 15200 13608 15264
rect 13672 15200 13688 15264
rect 13752 15200 13761 15264
rect 13440 14486 13761 15200
rect 13440 14250 13482 14486
rect 13718 14250 13761 14486
rect 13440 14176 13761 14250
rect 13440 14112 13448 14176
rect 13512 14112 13528 14176
rect 13592 14112 13608 14176
rect 13672 14112 13688 14176
rect 13752 14112 13761 14176
rect 13440 13088 13761 14112
rect 13440 13024 13448 13088
rect 13512 13024 13528 13088
rect 13592 13024 13608 13088
rect 13672 13024 13688 13088
rect 13752 13024 13761 13088
rect 13440 12000 13761 13024
rect 13440 11936 13448 12000
rect 13512 11936 13528 12000
rect 13592 11936 13608 12000
rect 13672 11936 13688 12000
rect 13752 11936 13761 12000
rect 13440 10912 13761 11936
rect 13440 10848 13448 10912
rect 13512 10848 13528 10912
rect 13592 10848 13608 10912
rect 13672 10848 13688 10912
rect 13752 10848 13761 10912
rect 13440 9824 13761 10848
rect 13440 9760 13448 9824
rect 13512 9760 13528 9824
rect 13592 9760 13608 9824
rect 13672 9760 13688 9824
rect 13752 9760 13761 9824
rect 13440 9590 13761 9760
rect 13440 9354 13482 9590
rect 13718 9354 13761 9590
rect 13440 8736 13761 9354
rect 13440 8672 13448 8736
rect 13512 8672 13528 8736
rect 13592 8672 13608 8736
rect 13672 8672 13688 8736
rect 13752 8672 13761 8736
rect 13440 7648 13761 8672
rect 13440 7584 13448 7648
rect 13512 7584 13528 7648
rect 13592 7584 13608 7648
rect 13672 7584 13688 7648
rect 13752 7584 13761 7648
rect 13440 6560 13761 7584
rect 13440 6496 13448 6560
rect 13512 6496 13528 6560
rect 13592 6496 13608 6560
rect 13672 6496 13688 6560
rect 13752 6496 13761 6560
rect 13440 5472 13761 6496
rect 13440 5408 13448 5472
rect 13512 5408 13528 5472
rect 13592 5408 13608 5472
rect 13672 5408 13688 5472
rect 13752 5408 13761 5472
rect 13440 4694 13761 5408
rect 13440 4458 13482 4694
rect 13718 4458 13761 4694
rect 13440 4384 13761 4458
rect 13440 4320 13448 4384
rect 13512 4320 13528 4384
rect 13592 4320 13608 4384
rect 13672 4320 13688 4384
rect 13752 4320 13761 4384
rect 13440 3296 13761 4320
rect 13440 3232 13448 3296
rect 13512 3232 13528 3296
rect 13592 3232 13608 3296
rect 13672 3232 13688 3296
rect 13752 3232 13761 3296
rect 13440 2208 13761 3232
rect 13440 2144 13448 2208
rect 13512 2144 13528 2208
rect 13592 2144 13608 2208
rect 13672 2144 13688 2208
rect 13752 2144 13761 2208
rect 13440 2128 13761 2144
<< via4 >>
rect 3485 14250 3721 14486
rect 3485 9354 3721 9590
rect 3485 4458 3721 4694
rect 5984 11802 6220 12038
rect 5984 7104 6220 7142
rect 5984 7040 6014 7104
rect 6014 7040 6030 7104
rect 6030 7040 6094 7104
rect 6094 7040 6110 7104
rect 6110 7040 6174 7104
rect 6174 7040 6190 7104
rect 6190 7040 6220 7104
rect 5984 6906 6220 7040
rect 8484 14250 8720 14486
rect 8484 9354 8720 9590
rect 8484 4458 8720 4694
rect 10983 11802 11219 12038
rect 10983 7104 11219 7142
rect 10983 7040 11013 7104
rect 11013 7040 11029 7104
rect 11029 7040 11093 7104
rect 11093 7040 11109 7104
rect 11109 7040 11173 7104
rect 11173 7040 11189 7104
rect 11189 7040 11219 7104
rect 10983 6906 11219 7040
rect 13482 14250 13718 14486
rect 13482 9354 13718 9590
rect 13482 4458 13718 4694
<< metal5 >>
rect 1104 14486 16100 14528
rect 1104 14250 3485 14486
rect 3721 14250 8484 14486
rect 8720 14250 13482 14486
rect 13718 14250 16100 14486
rect 1104 14208 16100 14250
rect 1104 12038 16100 12080
rect 1104 11802 5984 12038
rect 6220 11802 10983 12038
rect 11219 11802 16100 12038
rect 1104 11760 16100 11802
rect 1104 9590 16100 9632
rect 1104 9354 3485 9590
rect 3721 9354 8484 9590
rect 8720 9354 13482 9590
rect 13718 9354 16100 9590
rect 1104 9312 16100 9354
rect 1104 7142 16100 7184
rect 1104 6906 5984 7142
rect 6220 6906 10983 7142
rect 11219 6906 16100 7142
rect 1104 6864 16100 6906
rect 1104 4694 16100 4736
rect 1104 4458 3485 4694
rect 3721 4458 8484 4694
rect 8720 4458 13482 4694
rect 13718 4458 16100 4694
rect 1104 4416 16100 4458
use sky130_fd_sc_hd__o221a_1  _245_
timestamp 1623890261
transform -1 0 3496 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _293_
timestamp 1623890261
transform -1 0 2484 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _310_
timestamp 1623890261
transform 1 0 1380 0 -1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1623890261
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1623890261
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1623890261
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_6
timestamp 1623890261
transform 1 0 1656 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15
timestamp 1623890261
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _243_
timestamp 1623890261
transform -1 0 3772 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _251_
timestamp 1623890261
transform 1 0 3864 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1623890261
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1623890261
transform 1 0 3312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28
timestamp 1623890261
transform 1 0 3680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_29
timestamp 1623890261
transform 1 0 3772 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1623890261
transform -1 0 4968 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _296_
timestamp 1623890261
transform 1 0 4968 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_38
timestamp 1623890261
transform 1 0 4600 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1623890261
transform 1 0 5244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _307_
timestamp 1623890261
transform 1 0 3864 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _142_
timestamp 1623890261
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _247_
timestamp 1623890261
transform 1 0 5980 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp 1623890261
transform -1 0 5980 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output9
timestamp 1623890261
transform -1 0 6348 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_49
timestamp 1623890261
transform 1 0 5612 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1623890261
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1623890261
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1623890261
transform 1 0 6348 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59
timestamp 1623890261
transform 1 0 6532 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_58
timestamp 1623890261
transform 1 0 6440 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _241_
timestamp 1623890261
transform 1 0 6532 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _141_
timestamp 1623890261
transform -1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _250_
timestamp 1623890261
transform 1 0 7084 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1623890261
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70
timestamp 1623890261
transform 1 0 7544 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  _308_
timestamp 1623890261
transform 1 0 7360 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _295_
timestamp 1623890261
transform -1 0 8648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _319_
timestamp 1623890261
transform -1 0 11132 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1623890261
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78
timestamp 1623890261
transform 1 0 8280 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_82
timestamp 1623890261
transform 1 0 8648 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86
timestamp 1623890261
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_88
timestamp 1623890261
transform 1 0 9200 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100
timestamp 1623890261
transform 1 0 10304 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _158_
timestamp 1623890261
transform -1 0 11592 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _279_
timestamp 1623890261
transform -1 0 11316 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1623890261
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1623890261
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1623890261
transform 1 0 11960 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111
timestamp 1623890261
transform 1 0 11316 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115
timestamp 1623890261
transform 1 0 11684 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1623890261
transform 1 0 11868 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_115
timestamp 1623890261
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _299_
timestamp 1623890261
transform -1 0 13984 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _304_
timestamp 1623890261
transform 1 0 12788 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_0_121
timestamp 1623890261
transform 1 0 12236 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_133
timestamp 1623890261
transform 1 0 13340 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_140
timestamp 1623890261
transform 1 0 13984 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1623890261
transform -1 0 14996 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1623890261
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144
timestamp 1623890261
transform 1 0 14352 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_146
timestamp 1623890261
transform 1 0 14536 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_147
timestamp 1623890261
transform 1 0 14628 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_151
timestamp 1623890261
transform 1 0 14996 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1623890261
transform -1 0 16100 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1623890261
transform -1 0 16100 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1623890261
transform 1 0 15548 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_154
timestamp 1623890261
transform 1 0 15272 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_159
timestamp 1623890261
transform 1 0 15732 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1623890261
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1623890261
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1623890261
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _246_
timestamp 1623890261
transform 1 0 3956 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1623890261
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1623890261
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_30
timestamp 1623890261
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_38
timestamp 1623890261
transform 1 0 4600 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _248_
timestamp 1623890261
transform 1 0 7084 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _249_
timestamp 1623890261
transform 1 0 6256 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_2_50
timestamp 1623890261
transform 1 0 5704 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp 1623890261
transform -1 0 8740 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _163_
timestamp 1623890261
transform 1 0 9108 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _284_
timestamp 1623890261
transform 1 0 9844 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1623890261
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_72
timestamp 1623890261
transform 1 0 7728 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_83
timestamp 1623890261
transform 1 0 8740 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_94
timestamp 1623890261
transform 1 0 9752 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _324_
timestamp 1623890261
transform 1 0 10212 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _325_
timestamp 1623890261
transform -1 0 13892 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_2_98
timestamp 1623890261
transform 1 0 10120 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1623890261
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_139
timestamp 1623890261
transform 1 0 13892 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1623890261
transform -1 0 16100 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_144
timestamp 1623890261
transform 1 0 14352 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_156
timestamp 1623890261
transform 1 0 15456 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _311_
timestamp 1623890261
transform 1 0 1380 0 1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1623890261
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _167_
timestamp 1623890261
transform -1 0 6164 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_24
timestamp 1623890261
transform 1 0 3312 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_36
timestamp 1623890261
transform 1 0 4416 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_44
timestamp 1623890261
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _140_
timestamp 1623890261
transform -1 0 7360 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1623890261
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_55
timestamp 1623890261
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_58
timestamp 1623890261
transform 1 0 6440 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_64
timestamp 1623890261
transform 1 0 6992 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_68
timestamp 1623890261
transform 1 0 7360 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_80
timestamp 1623890261
transform 1 0 8464 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_92
timestamp 1623890261
transform 1 0 9568 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _157_
timestamp 1623890261
transform 1 0 11684 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1623890261
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1623890261
transform 1 0 10672 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_112
timestamp 1623890261
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _305_
timestamp 1623890261
transform 1 0 13984 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_3_122
timestamp 1623890261
transform 1 0 12328 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_134
timestamp 1623890261
transform 1 0 13432 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1623890261
transform -1 0 16100 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp 1623890261
transform -1 0 3036 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _244_
timestamp 1623890261
transform 1 0 2392 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp 1623890261
transform -1 0 2300 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1623890261
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1623890261
transform 1 0 1380 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_9
timestamp 1623890261
transform 1 0 1932 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_13
timestamp 1623890261
transform 1 0 2300 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_21
timestamp 1623890261
transform 1 0 3036 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _182_
timestamp 1623890261
transform -1 0 6256 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  _281_
timestamp 1623890261
transform 1 0 4140 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1623890261
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_30
timestamp 1623890261
transform 1 0 3864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_36
timestamp 1623890261
transform 1 0 4416 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_42
timestamp 1623890261
transform 1 0 4968 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _309_
timestamp 1623890261
transform 1 0 6900 0 -1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_6  FILLER_4_56
timestamp 1623890261
transform 1 0 6256 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_62
timestamp 1623890261
transform 1 0 6808 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _320_
timestamp 1623890261
transform -1 0 11224 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1623890261
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_87
timestamp 1623890261
transform 1 0 9108 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _154_
timestamp 1623890261
transform 1 0 11316 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _326_
timestamp 1623890261
transform -1 0 13800 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_4_110
timestamp 1623890261
transform 1 0 11224 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _297_
timestamp 1623890261
transform -1 0 14260 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1623890261
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1623890261
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _152_
timestamp 1623890261
transform -1 0 15824 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1623890261
transform -1 0 16100 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _322_
timestamp 1623890261
transform -1 0 5060 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1623890261
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1623890261
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 1623890261
transform 1 0 2484 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2ai_1  _180_
timestamp 1623890261
transform -1 0 5888 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_5_43
timestamp 1623890261
transform 1 0 5060 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__o2bb2a_1  _168_
timestamp 1623890261
transform 1 0 6440 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1623890261
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1623890261
transform 1 0 5888 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_56
timestamp 1623890261
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_66
timestamp 1623890261
transform 1 0 7176 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _162_
timestamp 1623890261
transform 1 0 9016 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp 1623890261
transform 1 0 8004 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_74
timestamp 1623890261
transform 1 0 7912 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_78
timestamp 1623890261
transform 1 0 8280 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_93
timestamp 1623890261
transform 1 0 9660 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _155_
timestamp 1623890261
transform -1 0 12788 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _200_
timestamp 1623890261
transform -1 0 11592 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _283_
timestamp 1623890261
transform 1 0 10304 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1623890261
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_99
timestamp 1623890261
transform 1 0 10212 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_103
timestamp 1623890261
transform 1 0 10580 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_115
timestamp 1623890261
transform 1 0 11684 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _301_
timestamp 1623890261
transform 1 0 12972 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _306_
timestamp 1623890261
transform 1 0 13800 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 1623890261
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_132
timestamp 1623890261
transform 1 0 13248 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1623890261
transform -1 0 16100 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_158
timestamp 1623890261
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _159_
timestamp 1623890261
transform 1 0 2484 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _280_
timestamp 1623890261
transform 1 0 1932 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _323_
timestamp 1623890261
transform -1 0 3220 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1623890261
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1623890261
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_23
timestamp 1623890261
transform 1 0 3220 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1623890261
transform 1 0 1380 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_12
timestamp 1623890261
transform 1 0 2208 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_22
timestamp 1623890261
transform 1 0 3128 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _160_
timestamp 1623890261
transform 1 0 3864 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _164_
timestamp 1623890261
transform -1 0 4140 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _184_
timestamp 1623890261
transform -1 0 5704 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1623890261
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_37
timestamp 1623890261
transform 1 0 4508 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_33
timestamp 1623890261
transform 1 0 4140 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _169_
timestamp 1623890261
transform 1 0 6256 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _181_
timestamp 1623890261
transform -1 0 5980 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1623890261
transform 1 0 5980 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1623890261
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_49
timestamp 1623890261
transform 1 0 5612 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_55
timestamp 1623890261
transform 1 0 6164 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_56
timestamp 1623890261
transform 1 0 6256 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_58
timestamp 1623890261
transform 1 0 6440 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _171_
timestamp 1623890261
transform 1 0 6992 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_63
timestamp 1623890261
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _161_
timestamp 1623890261
transform 1 0 8280 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _166_
timestamp 1623890261
transform 1 0 8096 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _173_
timestamp 1623890261
transform 1 0 7728 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_75
timestamp 1623890261
transform 1 0 8004 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 1623890261
transform -1 0 9844 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1623890261
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1623890261
transform 1 0 8924 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_91
timestamp 1623890261
transform 1 0 9476 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _321_
timestamp 1623890261
transform -1 0 10948 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_7_79
timestamp 1623890261
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_95
timestamp 1623890261
transform 1 0 9844 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_4  _153_
timestamp 1623890261
transform 1 0 11132 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_8  _156_
timestamp 1623890261
transform 1 0 12052 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  ringosc.iss.ctrlen0
timestamp 1623890261
transform 1 0 11684 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1623890261
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_107
timestamp 1623890261
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_116
timestamp 1623890261
transform 1 0 11776 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_107
timestamp 1623890261
transform 1 0 10948 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 1623890261
transform 1 0 11500 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00
timestamp 1623890261
transform 1 0 13616 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1
timestamp 1623890261
transform 1 0 13156 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb0
timestamp 1623890261
transform 1 0 12144 0 1 5984
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1623890261
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_132
timestamp 1623890261
transform 1 0 13248 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_140
timestamp 1623890261
transform 1 0 13984 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_134
timestamp 1623890261
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_140
timestamp 1623890261
transform 1 0 13984 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01
timestamp 1623890261
transform 1 0 14352 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1623890261
transform -1 0 16100 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1623890261
transform -1 0 16100 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_157
timestamp 1623890261
transform 1 0 15548 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_152
timestamp 1623890261
transform 1 0 15088 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1623890261
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1623890261
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1623890261
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _165_
timestamp 1623890261
transform -1 0 5152 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _185_
timestamp 1623890261
transform 1 0 5152 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _187_
timestamp 1623890261
transform 1 0 3864 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1623890261
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1623890261
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _170_
timestamp 1623890261
transform 1 0 7268 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _172_
timestamp 1623890261
transform -1 0 6532 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _174_
timestamp 1623890261
transform 1 0 6532 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_48
timestamp 1623890261
transform 1 0 5520 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_70
timestamp 1623890261
transform 1 0 7544 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0
timestamp 1623890261
transform -1 0 9936 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1623890261
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_82
timestamp 1623890261
transform 1 0 8648 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_87
timestamp 1623890261
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1623890261
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.delayen0
timestamp 1623890261
transform -1 0 12052 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__einvn_2  ringosc.iss.delayenb1
timestamp 1623890261
transform 1 0 10212 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_8_96
timestamp 1623890261
transform 1 0 9936 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_106
timestamp 1623890261
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_119
timestamp 1623890261
transform 1 0 12052 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_4  ringosc.iss.reseten0
timestamp 1623890261
transform 1 0 12236 0 -1 7072
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1623890261
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_132
timestamp 1623890261
transform 1 0 13248 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_140
timestamp 1623890261
transform 1 0 13984 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1623890261
transform -1 0 16100 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1623890261
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_156
timestamp 1623890261
transform 1 0 15456 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _186_
timestamp 1623890261
transform 1 0 2760 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _189_
timestamp 1623890261
transform 1 0 2024 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1623890261
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1623890261
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1623890261
transform 1 0 1932 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _139_
timestamp 1623890261
transform 1 0 3404 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _151_
timestamp 1623890261
transform 1 0 5060 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_28
timestamp 1623890261
transform 1 0 3680 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_40
timestamp 1623890261
transform 1 0 4784 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_46
timestamp 1623890261
transform 1 0 5336 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1623890261
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_54
timestamp 1623890261
transform 1 0 6072 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1623890261
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_70
timestamp 1623890261
transform 1 0 7544 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb0
timestamp 1623890261
transform 1 0 8188 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_9_76
timestamp 1623890261
transform 1 0 8096 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_84
timestamp 1623890261
transform 1 0 8832 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1623890261
transform 1 0 11040 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.delayen1
timestamp 1623890261
transform 1 0 10396 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1623890261
transform 1 0 11316 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1623890261
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_96
timestamp 1623890261
transform 1 0 9936 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_100
timestamp 1623890261
transform 1 0 10304 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1623890261
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_115
timestamp 1623890261
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb0
timestamp 1623890261
transform 1 0 13984 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_9_127
timestamp 1623890261
transform 1 0 12788 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_139
timestamp 1623890261
transform 1 0 13892 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen0
timestamp 1623890261
transform 1 0 14628 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1623890261
transform -1 0 16100 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_152
timestamp 1623890261
transform 1 0 15088 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _188_
timestamp 1623890261
transform -1 0 3404 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o221ai_2  _192_
timestamp 1623890261
transform 1 0 1840 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1623890261
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1623890261
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1623890261
transform 1 0 1748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o2111ai_4  _199_
timestamp 1623890261
transform 1 0 4232 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1623890261
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_25
timestamp 1623890261
transform 1 0 3404 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_30
timestamp 1623890261
transform 1 0 3864 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[0\].id.delayenb1
timestamp 1623890261
transform 1 0 7268 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_10_55
timestamp 1623890261
transform 1 0 6164 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1623890261
transform 1 0 8648 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen0
timestamp 1623890261
transform 1 0 8188 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1623890261
transform 1 0 9476 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1623890261
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_74
timestamp 1623890261
transform 1 0 7912 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1623890261
transform 1 0 8924 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1623890261
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_95
timestamp 1623890261
transform 1 0 9844 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  ringosc.dstage\[11\].id.delayen0
timestamp 1623890261
transform 1 0 11776 0 -1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_10_107
timestamp 1623890261
transform 1 0 10948 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_115
timestamp 1623890261
transform 1 0 11684 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1623890261
transform 1 0 13432 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1623890261
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_137
timestamp 1623890261
transform 1 0 13708 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1623890261
transform 1 0 14720 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1623890261
transform -1 0 14720 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1623890261
transform -1 0 16100 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_151
timestamp 1623890261
transform 1 0 14996 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_159
timestamp 1623890261
transform 1 0 15732 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_2  _190_
timestamp 1623890261
transform -1 0 2576 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1623890261
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1623890261
transform 1 0 1380 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_16
timestamp 1623890261
transform 1 0 2576 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _191_
timestamp 1623890261
transform -1 0 5520 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _208_
timestamp 1623890261
transform 1 0 3864 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_28
timestamp 1623890261
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__a22oi_2  _175_
timestamp 1623890261
transform 1 0 6440 0 1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _178_
timestamp 1623890261
transform 1 0 5612 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[0\].id.delayen1
timestamp 1623890261
transform 1 0 7360 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1623890261
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_48
timestamp 1623890261
transform 1 0 5520 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 1623890261
transform 1 0 8188 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_73
timestamp 1623890261
transform 1 0 7820 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_80
timestamp 1623890261
transform 1 0 8464 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_92
timestamp 1623890261
transform 1 0 9568 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp 1623890261
transform 1 0 11776 0 1 8160
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb0
timestamp 1623890261
transform 1 0 9936 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1623890261
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_103
timestamp 1623890261
transform 1 0 10580 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_111
timestamp 1623890261
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_115
timestamp 1623890261
transform 1 0 11684 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[10\].id.delayenb1
timestamp 1623890261
transform 1 0 14168 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen1
timestamp 1623890261
transform -1 0 14076 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_11_141
timestamp 1623890261
transform 1 0 14076 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1623890261
transform 1 0 15272 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[10\].id.delayen1
timestamp 1623890261
transform 1 0 14812 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1623890261
transform -1 0 16100 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_157
timestamp 1623890261
transform 1 0 15548 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _312_
timestamp 1623890261
transform 1 0 1380 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1623890261
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_23
timestamp 1623890261
transform 1 0 3220 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1623890261
transform 1 0 5152 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _193_
timestamp 1623890261
transform 1 0 4508 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _207_
timestamp 1623890261
transform 1 0 3864 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1623890261
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_36
timestamp 1623890261
transform 1 0 4416 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_47
timestamp 1623890261
transform 1 0 5428 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _176_
timestamp 1623890261
transform -1 0 6440 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1623890261
transform -1 0 5980 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_58
timestamp 1623890261
transform 1 0 6440 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_70
timestamp 1623890261
transform 1 0 7544 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen1
timestamp 1623890261
transform -1 0 10212 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[1\].id.delayenb1
timestamp 1623890261
transform 1 0 9108 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1623890261
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_82
timestamp 1623890261
transform 1 0 8648 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[1\].id.delayen0
timestamp 1623890261
transform 1 0 10212 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1623890261
transform 1 0 10672 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_107
timestamp 1623890261
transform 1 0 10948 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_119
timestamp 1623890261
transform 1 0 12052 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _300_
timestamp 1623890261
transform 1 0 13524 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[11\].id.delayenb1
timestamp 1623890261
transform 1 0 12512 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  ringosc.dstage\[11\].id.delayint0
timestamp 1623890261
transform -1 0 13524 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1623890261
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_123
timestamp 1623890261
transform 1 0 12420 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_138
timestamp 1623890261
transform 1 0 13800 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_142
timestamp 1623890261
transform 1 0 14168 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1623890261
transform -1 0 16100 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_144
timestamp 1623890261
transform 1 0 14352 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_156
timestamp 1623890261
transform 1 0 15456 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _291_
timestamp 1623890261
transform -1 0 2300 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1623890261
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1623890261
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1623890261
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_6
timestamp 1623890261
transform 1 0 1656 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _150_
timestamp 1623890261
transform -1 0 3404 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _240_
timestamp 1623890261
transform 1 0 2484 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_13_13
timestamp 1623890261
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_15
timestamp 1623890261
transform 1 0 2484 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_23
timestamp 1623890261
transform 1 0 3220 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1623890261
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _149_
timestamp 1623890261
transform -1 0 3772 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_4  _209_
timestamp 1623890261
transform -1 0 5520 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1623890261
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_25
timestamp 1623890261
transform 1 0 3404 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_37
timestamp 1623890261
transform 1 0 4508 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_30
timestamp 1623890261
transform 1 0 3864 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _235_
timestamp 1623890261
transform -1 0 6440 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _288_
timestamp 1623890261
transform -1 0 6808 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1623890261
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_49
timestamp 1623890261
transform 1 0 5612 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_48
timestamp 1623890261
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_58
timestamp 1623890261
transform 1 0 6440 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _265_
timestamp 1623890261
transform 1 0 7268 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_14_62
timestamp 1623890261
transform 1 0 6808 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_66
timestamp 1623890261
transform 1 0 7176 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _315_
timestamp 1623890261
transform 1 0 6440 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_2  _206_
timestamp 1623890261
transform -1 0 8832 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1623890261
transform -1 0 9844 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1623890261
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_84
timestamp 1623890261
transform 1 0 8832 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_95
timestamp 1623890261
transform 1 0 9844 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_74
timestamp 1623890261
transform 1 0 7912 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_87
timestamp 1623890261
transform 1 0 9108 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_95
timestamp 1623890261
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__o41a_2  _261_
timestamp 1623890261
transform 1 0 11684 0 -1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _263_
timestamp 1623890261
transform 1 0 10028 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1623890261
transform 1 0 10856 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1623890261
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_103
timestamp 1623890261
transform 1 0 10580 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_110
timestamp 1623890261
transform 1 0 11224 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_115
timestamp 1623890261
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_104
timestamp 1623890261
transform 1 0 10672 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_112
timestamp 1623890261
transform 1 0 11408 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _259_
timestamp 1623890261
transform -1 0 13432 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _262_
timestamp 1623890261
transform 1 0 13432 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1623890261
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_127
timestamp 1623890261
transform 1 0 12788 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_139
timestamp 1623890261
transform 1 0 13892 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_139
timestamp 1623890261
transform 1 0 13892 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1623890261
transform -1 0 15456 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen0
timestamp 1623890261
transform -1 0 15456 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb0
timestamp 1623890261
transform 1 0 14352 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1623890261
transform -1 0 16100 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1623890261
transform -1 0 16100 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1623890261
transform -1 0 15824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_151
timestamp 1623890261
transform 1 0 14996 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_156
timestamp 1623890261
transform 1 0 15456 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_156
timestamp 1623890261
transform 1 0 15456 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_1  _238_
timestamp 1623890261
transform 1 0 3036 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o22ai_1  _239_
timestamp 1623890261
transform 1 0 2576 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp 1623890261
transform -1 0 2208 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1623890261
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1623890261
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_12
timestamp 1623890261
transform 1 0 2208 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _211_
timestamp 1623890261
transform -1 0 4416 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _212_
timestamp 1623890261
transform -1 0 5060 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _234_
timestamp 1623890261
transform -1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1623890261
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_51
timestamp 1623890261
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_58
timestamp 1623890261
transform 1 0 6440 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_70
timestamp 1623890261
transform 1 0 7544 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_2  _270_
timestamp 1623890261
transform -1 0 8832 0 1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _271_
timestamp 1623890261
transform 1 0 8832 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_93
timestamp 1623890261
transform 1 0 9660 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _256_
timestamp 1623890261
transform 1 0 11684 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1623890261
transform 1 0 11040 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen1
timestamp 1623890261
transform 1 0 10580 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb1
timestamp 1623890261
transform 1 0 9936 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1623890261
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_111
timestamp 1623890261
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[9\].id.delayen1
timestamp 1623890261
transform 1 0 13892 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[9\].id.delayenb1
timestamp 1623890261
transform 1 0 13248 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_15_122
timestamp 1623890261
transform 1 0 12328 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_130
timestamp 1623890261
transform 1 0 13064 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1623890261
transform 1 0 14352 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1623890261
transform 1 0 14628 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1623890261
transform -1 0 16100 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_150
timestamp 1623890261
transform 1 0 14904 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_158
timestamp 1623890261
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _313_
timestamp 1623890261
transform 1 0 1380 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1623890261
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_23
timestamp 1623890261
transform 1 0 3220 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _198_
timestamp 1623890261
transform 1 0 4232 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _233_
timestamp 1623890261
transform 1 0 4968 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1623890261
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_30
timestamp 1623890261
transform 1 0 3864 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_39
timestamp 1623890261
transform 1 0 4692 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _147_
timestamp 1623890261
transform 1 0 7636 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _274_
timestamp 1623890261
transform -1 0 7636 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_51
timestamp 1623890261
transform 1 0 5796 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_59
timestamp 1623890261
transform 1 0 6532 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _272_
timestamp 1623890261
transform 1 0 9108 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1623890261
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_74
timestamp 1623890261
transform 1 0 7912 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_95
timestamp 1623890261
transform 1 0 9844 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1623890261
transform 1 0 10856 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_103
timestamp 1623890261
transform 1 0 10580 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1623890261
transform 1 0 11132 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1623890261
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1623890261
transform 1 0 12236 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_133
timestamp 1623890261
transform 1 0 13340 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1623890261
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1623890261
transform -1 0 15456 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1623890261
transform -1 0 16100 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_144
timestamp 1623890261
transform 1 0 14352 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_156
timestamp 1623890261
transform 1 0 15456 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1623890261
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1623890261
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1623890261
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1623890261
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1623890261
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _148_
timestamp 1623890261
transform 1 0 6072 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _195_
timestamp 1623890261
transform -1 0 6992 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1623890261
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_51
timestamp 1623890261
transform 1 0 5796 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_58
timestamp 1623890261
transform 1 0 6440 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_64
timestamp 1623890261
transform 1 0 6992 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_2  _268_
timestamp 1623890261
transform 1 0 9292 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _269_
timestamp 1623890261
transform 1 0 8556 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_76
timestamp 1623890261
transform 1 0 8096 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_80
timestamp 1623890261
transform 1 0 8464 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_95
timestamp 1623890261
transform 1 0 9844 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_2  _258_
timestamp 1623890261
transform 1 0 12052 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[2\].id.delayen0
timestamp 1623890261
transform 1 0 10672 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[2\].id.delayenb0
timestamp 1623890261
transform 1 0 9936 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1623890261
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_103
timestamp 1623890261
transform 1 0 10580 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_109
timestamp 1623890261
transform 1 0 11132 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1623890261
transform 1 0 11500 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_115
timestamp 1623890261
transform 1 0 11684 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_126
timestamp 1623890261
transform 1 0 12696 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_138
timestamp 1623890261
transform 1 0 13800 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1623890261
transform -1 0 16100 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_150
timestamp 1623890261
transform 1 0 14904 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_158
timestamp 1623890261
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _314_
timestamp 1623890261
transform -1 0 3312 0 -1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1623890261
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _194_
timestamp 1623890261
transform 1 0 4600 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _215_
timestamp 1623890261
transform -1 0 5704 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _236_
timestamp 1623890261
transform 1 0 3496 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _237_
timestamp 1623890261
transform 1 0 3864 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1623890261
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_24
timestamp 1623890261
transform 1 0 3312 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_41
timestamp 1623890261
transform 1 0 4876 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1623890261
transform 1 0 7268 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _197_
timestamp 1623890261
transform 1 0 6440 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _214_
timestamp 1623890261
transform -1 0 6348 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _278_
timestamp 1623890261
transform 1 0 7544 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_57
timestamp 1623890261
transform 1 0 6348 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp 1623890261
transform -1 0 8556 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _257_
timestamp 1623890261
transform 1 0 9844 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _267_
timestamp 1623890261
transform -1 0 9844 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1623890261
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_81
timestamp 1623890261
transform 1 0 8556 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1623890261
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1623890261
transform 1 0 11316 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_102
timestamp 1623890261
transform 1 0 10488 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_110
timestamp 1623890261
transform 1 0 11224 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_115
timestamp 1623890261
transform 1 0 11684 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_119
timestamp 1623890261
transform 1 0 12052 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o31a_1  _255_
timestamp 1623890261
transform -1 0 12788 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _276_
timestamp 1623890261
transform -1 0 13248 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb1
timestamp 1623890261
transform 1 0 13248 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1623890261
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_139
timestamp 1623890261
transform 1 0 13892 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen0
timestamp 1623890261
transform -1 0 15456 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[8\].id.delayenb0
timestamp 1623890261
transform 1 0 14352 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1623890261
transform -1 0 16100 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_156
timestamp 1623890261
transform 1 0 15456 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _289_
timestamp 1623890261
transform 1 0 2116 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1623890261
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1623890261
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1623890261
transform 1 0 1380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_14
timestamp 1623890261
transform 1 0 2392 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1623890261
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1623890261
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _232_
timestamp 1623890261
transform 1 0 3680 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1623890261
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_26
timestamp 1623890261
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1623890261
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_30
timestamp 1623890261
transform 1 0 3864 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _216_
timestamp 1623890261
transform -1 0 5428 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _230_
timestamp 1623890261
transform 1 0 5428 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_45
timestamp 1623890261
transform 1 0 5244 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_38
timestamp 1623890261
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_33
timestamp 1623890261
transform 1 0 4140 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _213_
timestamp 1623890261
transform 1 0 5612 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1623890261
transform 1 0 5888 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_50
timestamp 1623890261
transform 1 0 5704 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _146_
timestamp 1623890261
transform 1 0 6256 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _203_
timestamp 1623890261
transform 1 0 6900 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _254_
timestamp 1623890261
transform 1 0 6532 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1623890261
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_56
timestamp 1623890261
transform 1 0 6256 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_58
timestamp 1623890261
transform 1 0 6440 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_59
timestamp 1623890261
transform 1 0 6532 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _201_
timestamp 1623890261
transform 1 0 7176 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _264_
timestamp 1623890261
transform -1 0 8188 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _205_
timestamp 1623890261
transform 1 0 7912 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _266_
timestamp 1623890261
transform 1 0 8556 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _303_
timestamp 1623890261
transform -1 0 9936 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1623890261
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_73
timestamp 1623890261
transform 1 0 7820 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_79
timestamp 1623890261
transform 1 0 8372 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_91
timestamp 1623890261
transform 1 0 9476 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_77
timestamp 1623890261
transform 1 0 8188 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _273_
timestamp 1623890261
transform 1 0 9936 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb1
timestamp 1623890261
transform 1 0 10580 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_19_103
timestamp 1623890261
transform 1 0 10580 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_101
timestamp 1623890261
transform 1 0 10396 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1623890261
transform 1 0 11684 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen1
timestamp 1623890261
transform 1 0 11224 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1623890261
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_111
timestamp 1623890261
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_118
timestamp 1623890261
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_115
timestamp 1623890261
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _252_
timestamp 1623890261
transform 1 0 12144 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _277_
timestamp 1623890261
transform -1 0 13432 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1623890261
transform 1 0 14076 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[8\].id.delayen1
timestamp 1623890261
transform 1 0 13340 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1623890261
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_127
timestamp 1623890261
transform 1 0 12788 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_138
timestamp 1623890261
transform 1 0 13800 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_134
timestamp 1623890261
transform 1 0 13432 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_142
timestamp 1623890261
transform 1 0 14168 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1623890261
transform -1 0 15456 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1623890261
transform 1 0 14352 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1623890261
transform -1 0 16100 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1623890261
transform -1 0 16100 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1623890261
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_159
timestamp 1623890261
transform 1 0 15732 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_144
timestamp 1623890261
transform 1 0 14352 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_156
timestamp 1623890261
transform 1 0 15456 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _316_
timestamp 1623890261
transform -1 0 3312 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1623890261
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _217_
timestamp 1623890261
transform 1 0 5428 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _219_
timestamp 1623890261
transform 1 0 4692 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _221_
timestamp 1623890261
transform 1 0 4048 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _223_
timestamp 1623890261
transform -1 0 4048 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1623890261
transform -1 0 7268 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1623890261
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_54
timestamp 1623890261
transform 1 0 6072 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_58
timestamp 1623890261
transform 1 0 6440 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_67
timestamp 1623890261
transform 1 0 7268 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__o41a_1  _260_
timestamp 1623890261
transform 1 0 9200 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_79
timestamp 1623890261
transform 1 0 8372 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_87
timestamp 1623890261
transform 1 0 9108 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1623890261
transform 1 0 11684 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1623890261
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_97
timestamp 1623890261
transform 1 0 10028 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_109
timestamp 1623890261
transform 1 0 11132 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1623890261
transform 1 0 11500 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_118
timestamp 1623890261
transform 1 0 11960 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1623890261
transform 1 0 13892 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb0
timestamp 1623890261
transform 1 0 14168 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[7\].id.delayenb1
timestamp 1623890261
transform 1 0 13156 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_21_130
timestamp 1623890261
transform 1 0 13064 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_138
timestamp 1623890261
transform 1 0 13800 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen0
timestamp 1623890261
transform -1 0 15272 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1623890261
transform -1 0 16100 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_154
timestamp 1623890261
transform 1 0 15272 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1623890261
transform -1 0 3496 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _287_
timestamp 1623890261
transform -1 0 2208 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1623890261
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1623890261
transform 1 0 1380 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_12
timestamp 1623890261
transform 1 0 2208 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_20
timestamp 1623890261
transform 1 0 2944 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1623890261
transform 1 0 3496 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _225_
timestamp 1623890261
transform -1 0 5244 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _226_
timestamp 1623890261
transform -1 0 5612 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _231_
timestamp 1623890261
transform 1 0 3864 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1623890261
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_38
timestamp 1623890261
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen1
timestamp 1623890261
transform 1 0 7544 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb1
timestamp 1623890261
transform 1 0 6900 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_22_49
timestamp 1623890261
transform 1 0 5612 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_61
timestamp 1623890261
transform 1 0 6716 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1623890261
transform 1 0 8004 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1623890261
transform 1 0 8280 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1623890261
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_81
timestamp 1623890261
transform 1 0 8556 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1623890261
transform 1 0 8924 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_87
timestamp 1623890261
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[3\].id.delayen0
timestamp 1623890261
transform 1 0 11224 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[3\].id.delayenb0
timestamp 1623890261
transform 1 0 10488 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_22_99
timestamp 1623890261
transform 1 0 10212 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_109
timestamp 1623890261
transform 1 0 11132 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_115
timestamp 1623890261
transform 1 0 11684 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _253_
timestamp 1623890261
transform 1 0 12788 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[7\].id.delayen1
timestamp 1623890261
transform 1 0 13248 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1623890261
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_137
timestamp 1623890261
transform 1 0 13708 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1623890261
transform 1 0 14352 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1623890261
transform -1 0 16100 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_147
timestamp 1623890261
transform 1 0 14628 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_159
timestamp 1623890261
transform 1 0 15732 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1623890261
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1623890261
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1623890261
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1623890261
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1623890261
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_4  _144_
timestamp 1623890261
transform 1 0 6440 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1623890261
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_51
timestamp 1623890261
transform 1 0 5796 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_65
timestamp 1623890261
transform 1 0 7084 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[4\].id.delayen0
timestamp 1623890261
transform -1 0 9568 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[4\].id.delayenb0
timestamp 1623890261
transform -1 0 9108 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_23_77
timestamp 1623890261
transform 1 0 8188 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_92
timestamp 1623890261
transform 1 0 9568 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1623890261
transform -1 0 12052 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1623890261
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_104
timestamp 1623890261
transform 1 0 10672 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_112
timestamp 1623890261
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_119
timestamp 1623890261
transform 1 0 12052 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_131
timestamp 1623890261
transform 1 0 13156 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_143
timestamp 1623890261
transform 1 0 14260 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1623890261
transform -1 0 16100 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_155
timestamp 1623890261
transform 1 0 15364 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_159
timestamp 1623890261
transform 1 0 15732 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _210_
timestamp 1623890261
transform 1 0 3220 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _224_
timestamp 1623890261
transform -1 0 3220 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1623890261
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1623890261
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_15
timestamp 1623890261
transform 1 0 2484 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _228_
timestamp 1623890261
transform 1 0 4048 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _285_
timestamp 1623890261
transform 1 0 3496 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _317_
timestamp 1623890261
transform 1 0 4784 0 -1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1623890261
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_30
timestamp 1623890261
transform 1 0 3864 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_2  _275_
timestamp 1623890261
transform 1 0 6716 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_24_66
timestamp 1623890261
transform 1 0 7176 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1623890261
transform -1 0 9752 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1623890261
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_78
timestamp 1623890261
transform 1 0 8280 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_87
timestamp 1623890261
transform 1 0 9108 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_94
timestamp 1623890261
transform 1 0 9752 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_106
timestamp 1623890261
transform 1 0 10856 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_118
timestamp 1623890261
transform 1 0 11960 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen0
timestamp 1623890261
transform -1 0 14260 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[6\].id.delayen1
timestamp 1623890261
transform 1 0 13156 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb1
timestamp 1623890261
transform 1 0 12512 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1623890261
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_136
timestamp 1623890261
transform 1 0 13616 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[6\].id.delayenb0
timestamp 1623890261
transform 1 0 14352 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1623890261
transform -1 0 15364 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1623890261
transform -1 0 16100 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_155
timestamp 1623890261
transform 1 0 15364 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_159
timestamp 1623890261
transform 1 0 15732 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _318_
timestamp 1623890261
transform 1 0 2116 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1623890261
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1623890261
transform 1 0 1380 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1623890261
transform -1 0 5336 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1623890261
transform 1 0 5336 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _229_
timestamp 1623890261
transform -1 0 5060 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_32
timestamp 1623890261
transform 1 0 4048 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_38
timestamp 1623890261
transform 1 0 4600 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _145_
timestamp 1623890261
transform -1 0 6716 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp 1623890261
transform -1 0 5980 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_2  ringosc.dstage\[5\].id.delayenb1
timestamp 1623890261
transform 1 0 7268 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1623890261
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_49
timestamp 1623890261
transform 1 0 5612 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_53
timestamp 1623890261
transform 1 0 5980 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_61
timestamp 1623890261
transform 1 0 6716 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1623890261
transform 1 0 8372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.dstage\[5\].id.delayen1
timestamp 1623890261
transform 1 0 7912 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb0
timestamp 1623890261
transform -1 0 10212 0 1 15776
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1623890261
transform 1 0 8648 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_85
timestamp 1623890261
transform 1 0 8924 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1623890261
transform 1 0 10212 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__inv_1  ringosc.ibufp10
timestamp 1623890261
transform -1 0 11592 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ringosc.ibufp11
timestamp 1623890261
transform -1 0 11132 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1623890261
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_109
timestamp 1623890261
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_115
timestamp 1623890261
transform 1 0 11684 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1623890261
transform 1 0 12604 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1623890261
transform -1 0 13524 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1623890261
transform 1 0 13708 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1623890261
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_129
timestamp 1623890261
transform 1 0 12972 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_135
timestamp 1623890261
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_140
timestamp 1623890261
transform 1 0 13984 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1623890261
transform -1 0 16100 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_152
timestamp 1623890261
transform 1 0 15088 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1623890261
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1623890261
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_6
timestamp 1623890261
transform 1 0 1656 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_18
timestamp 1623890261
transform 1 0 2760 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1623890261
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1623890261
transform -1 0 5336 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_26
timestamp 1623890261
transform 1 0 3496 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1623890261
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_42
timestamp 1623890261
transform 1 0 4968 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_46
timestamp 1623890261
transform 1 0 5336 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1623890261
transform 1 0 6440 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_59
timestamp 1623890261
transform 1 0 6532 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_71
timestamp 1623890261
transform 1 0 7636 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1623890261
transform 1 0 9108 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_83
timestamp 1623890261
transform 1 0 8740 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_88
timestamp 1623890261
transform 1 0 9200 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1623890261
transform 1 0 11776 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output10
timestamp 1623890261
transform -1 0 11408 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_100
timestamp 1623890261
transform 1 0 10304 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_112
timestamp 1623890261
transform 1 0 11408 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1623890261
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1623890261
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1623890261
transform 1 0 14076 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1623890261
transform -1 0 16100 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1623890261
transform 1 0 14444 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1623890261
transform -1 0 15824 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_146
timestamp 1623890261
transform 1 0 14536 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_154
timestamp 1623890261
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
<< labels >>
rlabel metal2 s 5998 0 6054 800 4 clockp[0]
port 1 nsew
rlabel metal2 s 11058 18590 11114 19390 4 clockp[1]
port 2 nsew
rlabel metal2 s 5078 18590 5134 19390 4 div[0]
port 3 nsew
rlabel metal2 s 478 0 534 800 4 div[1]
port 4 nsew
rlabel metal2 s 16578 18590 16634 19390 4 div[2]
port 5 nsew
rlabel metal3 s 0 8848 800 8968 4 div[3]
port 6 nsew
rlabel metal3 s 0 17688 800 17808 4 div[4]
port 7 nsew
rlabel metal2 s 11978 0 12034 800 4 enable
port 8 nsew
rlabel metal3 s 16446 1368 17246 1488 4 osc
port 9 nsew
rlabel metal3 s 16446 10208 17246 10328 4 resetb
port 10 nsew
rlabel metal4 s 13441 2128 13761 16912 4 VPWR
port 11 nsew
rlabel metal4 s 8442 2128 8762 16912 4 VPWR
port 11 nsew
rlabel metal4 s 3443 2128 3763 16912 4 VPWR
port 11 nsew
rlabel metal5 s 1104 14208 16100 14528 4 VPWR
port 11 nsew
rlabel metal5 s 1104 9312 16100 9632 4 VPWR
port 11 nsew
rlabel metal5 s 1104 4416 16100 4736 4 VPWR
port 11 nsew
rlabel metal4 s 10941 2128 11261 16912 4 VGND
port 12 nsew
rlabel metal4 s 5943 2128 6263 16912 4 VGND
port 12 nsew
rlabel metal5 s 1104 11760 16100 12080 4 VGND
port 12 nsew
rlabel metal5 s 1104 6864 16100 7184 4 VGND
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 17246 19390
<< end >>
