magic
tech sky130A
magscale 1 2
timestamp 1619632579
<< obsli1 >>
rect 1104 2159 21959 22865
<< obsm1 >>
rect 474 2128 22158 22896
<< metal2 >>
rect 938 24323 994 25123
rect 2778 24323 2834 25123
rect 4618 24323 4674 25123
rect 5998 24323 6054 25123
rect 7838 24323 7894 25123
rect 9678 24323 9734 25123
rect 11518 24323 11574 25123
rect 12898 24323 12954 25123
rect 14738 24323 14794 25123
rect 16578 24323 16634 25123
rect 17958 24323 18014 25123
rect 19798 24323 19854 25123
rect 21638 24323 21694 25123
rect 478 0 534 800
rect 1858 0 1914 800
rect 3698 0 3754 800
rect 5538 0 5594 800
rect 6918 0 6974 800
rect 8758 0 8814 800
rect 10598 0 10654 800
rect 11978 0 12034 800
rect 13818 0 13874 800
rect 15658 0 15714 800
rect 17038 0 17094 800
rect 18878 0 18934 800
rect 20718 0 20774 800
rect 22098 0 22154 800
<< obsm2 >>
rect 480 24267 882 24323
rect 1050 24267 2722 24323
rect 2890 24267 4562 24323
rect 4730 24267 5942 24323
rect 6110 24267 7782 24323
rect 7950 24267 9622 24323
rect 9790 24267 11462 24323
rect 11630 24267 12842 24323
rect 13010 24267 14682 24323
rect 14850 24267 16522 24323
rect 16690 24267 17902 24323
rect 18070 24267 19742 24323
rect 19910 24267 21582 24323
rect 21750 24267 22152 24323
rect 480 856 22152 24267
rect 590 800 1802 856
rect 1970 800 3642 856
rect 3810 800 5482 856
rect 5650 800 6862 856
rect 7030 800 8702 856
rect 8870 800 10542 856
rect 10710 800 11922 856
rect 12090 800 13762 856
rect 13930 800 15602 856
rect 15770 800 16982 856
rect 17150 800 18822 856
rect 18990 800 20662 856
rect 20830 800 22042 856
<< metal3 >>
rect 0 23128 800 23248
rect 22179 23128 22979 23248
rect 0 20408 800 20528
rect 22179 20408 22979 20528
rect 0 17688 800 17808
rect 22179 17688 22979 17808
rect 0 15648 800 15768
rect 22179 15648 22979 15768
rect 0 12928 800 13048
rect 22179 12928 22979 13048
rect 0 10208 800 10328
rect 22179 10208 22979 10328
rect 0 8168 800 8288
rect 22179 8168 22979 8288
rect 0 5448 800 5568
rect 22179 5448 22979 5568
rect 0 2728 800 2848
rect 22179 2728 22979 2848
<< obsm3 >>
rect 880 23048 22099 23221
rect 800 20608 22179 23048
rect 880 20328 22099 20608
rect 800 17888 22179 20328
rect 880 17608 22099 17888
rect 800 15848 22179 17608
rect 880 15568 22099 15848
rect 800 13128 22179 15568
rect 880 12848 22099 13128
rect 800 10408 22179 12848
rect 880 10128 22099 10408
rect 800 8368 22179 10128
rect 880 8088 22099 8368
rect 800 5648 22179 8088
rect 880 5368 22099 5648
rect 800 2928 22179 5368
rect 880 2648 22099 2928
rect 800 2143 22179 2648
<< metal4 >>
rect 4394 2128 4714 22896
rect 7844 2128 8164 22896
rect 11294 2128 11614 22896
rect 14744 2128 15064 22896
rect 18194 2128 18514 22896
<< metal5 >>
rect 1104 19195 21804 19515
rect 1104 15749 21804 16069
rect 1104 12304 21804 12624
rect 1104 8859 21804 9179
rect 1104 5413 21804 5733
<< obsm5 >>
rect 1104 16389 21804 18875
rect 1104 12944 21804 15429
rect 1104 9499 21804 11984
<< labels >>
rlabel metal3 s 0 10208 800 10328 6 clockc
port 1 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 clockd[0]
port 2 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 clockd[1]
port 3 nsew signal output
rlabel metal3 s 22179 20408 22979 20528 6 clockd[2]
port 4 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 clockd[3]
port 5 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 clockp[0]
port 6 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 clockp[1]
port 7 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 dco
port 8 nsew signal input
rlabel metal3 s 22179 15648 22979 15768 6 div[0]
port 9 nsew signal input
rlabel metal2 s 19798 24323 19854 25123 6 div[1]
port 10 nsew signal input
rlabel metal2 s 7838 24323 7894 25123 6 div[2]
port 11 nsew signal input
rlabel metal2 s 478 0 534 800 6 div[3]
port 12 nsew signal input
rlabel metal2 s 14738 24323 14794 25123 6 div[4]
port 13 nsew signal input
rlabel metal2 s 16578 24323 16634 25123 6 ext_trim[0]
port 14 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 ext_trim[10]
port 15 nsew signal input
rlabel metal2 s 2778 24323 2834 25123 6 ext_trim[11]
port 16 nsew signal input
rlabel metal3 s 22179 5448 22979 5568 6 ext_trim[12]
port 17 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 ext_trim[13]
port 18 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 ext_trim[14]
port 19 nsew signal input
rlabel metal3 s 22179 17688 22979 17808 6 ext_trim[15]
port 20 nsew signal input
rlabel metal2 s 4618 24323 4674 25123 6 ext_trim[16]
port 21 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 ext_trim[17]
port 22 nsew signal input
rlabel metal2 s 5998 24323 6054 25123 6 ext_trim[18]
port 23 nsew signal input
rlabel metal3 s 22179 10208 22979 10328 6 ext_trim[19]
port 24 nsew signal input
rlabel metal2 s 12898 24323 12954 25123 6 ext_trim[1]
port 25 nsew signal input
rlabel metal2 s 11518 24323 11574 25123 6 ext_trim[20]
port 26 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 ext_trim[21]
port 27 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 ext_trim[22]
port 28 nsew signal input
rlabel metal3 s 22179 23128 22979 23248 6 ext_trim[23]
port 29 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 ext_trim[24]
port 30 nsew signal input
rlabel metal2 s 9678 24323 9734 25123 6 ext_trim[25]
port 31 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 ext_trim[2]
port 32 nsew signal input
rlabel metal3 s 22179 8168 22979 8288 6 ext_trim[3]
port 33 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 ext_trim[4]
port 34 nsew signal input
rlabel metal3 s 22179 12928 22979 13048 6 ext_trim[5]
port 35 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 ext_trim[6]
port 36 nsew signal input
rlabel metal2 s 938 24323 994 25123 6 ext_trim[7]
port 37 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 ext_trim[8]
port 38 nsew signal input
rlabel metal3 s 22179 2728 22979 2848 6 ext_trim[9]
port 39 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 extclk_sel
port 40 nsew signal input
rlabel metal2 s 17958 24323 18014 25123 6 osc
port 41 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 reset
port 42 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 sel[0]
port 43 nsew signal input
rlabel metal2 s 21638 24323 21694 25123 6 sel[1]
port 44 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 sel[2]
port 45 nsew signal input
rlabel metal4 s 18194 2128 18514 22896 6 VPWR
port 46 nsew power bidirectional
rlabel metal4 s 11294 2128 11614 22896 6 VPWR
port 47 nsew power bidirectional
rlabel metal4 s 4394 2128 4714 22896 6 VPWR
port 48 nsew power bidirectional
rlabel metal5 s 1104 19195 21804 19515 6 VPWR
port 49 nsew power bidirectional
rlabel metal5 s 1104 12304 21804 12624 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1104 5413 21804 5733 6 VPWR
port 51 nsew power bidirectional
rlabel metal4 s 14744 2128 15064 22896 6 VGND
port 52 nsew ground bidirectional
rlabel metal4 s 7844 2128 8164 22896 6 VGND
port 53 nsew ground bidirectional
rlabel metal5 s 1104 15749 21804 16069 6 VGND
port 54 nsew ground bidirectional
rlabel metal5 s 1104 8859 21804 9179 6 VGND
port 55 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 22979 25123
string LEFview TRUE
string GDS_FILE /openLANE_flow/designs/digital_pll/runs/sixth_run/results/magic/digital_pll.gds
string GDS_END 1462108
string GDS_START 590732
<< end >>

